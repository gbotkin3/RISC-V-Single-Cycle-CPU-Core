magic
tech sky130B
magscale 1 2
timestamp 1663363331
<< viali >>
rect 6469 54825 6503 54859
rect 14381 54825 14415 54859
rect 24777 54825 24811 54859
rect 29929 54825 29963 54859
rect 36369 54825 36403 54859
rect 38301 54825 38335 54859
rect 40877 54825 40911 54859
rect 47777 54825 47811 54859
rect 48605 54825 48639 54859
rect 51825 54825 51859 54859
rect 25237 54757 25271 54791
rect 3985 54689 4019 54723
rect 10977 54689 11011 54723
rect 12633 54689 12667 54723
rect 27353 54689 27387 54723
rect 27813 54689 27847 54723
rect 45201 54689 45235 54723
rect 1409 54621 1443 54655
rect 1685 54621 1719 54655
rect 4261 54621 4295 54655
rect 6653 54621 6687 54655
rect 7389 54621 7423 54655
rect 7849 54621 7883 54655
rect 10701 54621 10735 54655
rect 11897 54621 11931 54655
rect 12449 54621 12483 54655
rect 14565 54621 14599 54655
rect 17141 54621 17175 54655
rect 18705 54621 18739 54655
rect 19257 54621 19291 54655
rect 19533 54621 19567 54655
rect 23305 54621 23339 54655
rect 25421 54621 25455 54655
rect 28089 54621 28123 54655
rect 29745 54621 29779 54655
rect 32505 54621 32539 54655
rect 32689 54621 32723 54655
rect 36185 54621 36219 54655
rect 38945 54621 38979 54655
rect 40693 54621 40727 54655
rect 42809 54621 42843 54655
rect 43269 54621 43303 54655
rect 45477 54621 45511 54655
rect 47041 54621 47075 54655
rect 47593 54621 47627 54655
rect 49249 54621 49283 54655
rect 51181 54621 51215 54655
rect 51641 54621 51675 54655
rect 52929 54621 52963 54655
rect 53389 54621 53423 54655
rect 2789 54553 2823 54587
rect 22293 54553 22327 54587
rect 22477 54553 22511 54587
rect 23581 54553 23615 54587
rect 33149 54553 33183 54587
rect 33701 54553 33735 54587
rect 35265 54553 35299 54587
rect 2881 54485 2915 54519
rect 8033 54485 8067 54519
rect 15117 54485 15151 54519
rect 16957 54485 16991 54519
rect 17693 54485 17727 54519
rect 30481 54485 30515 54519
rect 31033 54485 31067 54519
rect 32597 54485 32631 54519
rect 35173 54485 35207 54519
rect 38853 54485 38887 54519
rect 40141 54485 40175 54519
rect 42625 54485 42659 54519
rect 49157 54485 49191 54519
rect 53573 54485 53607 54519
rect 2605 54281 2639 54315
rect 3893 54281 3927 54315
rect 6745 54281 6779 54315
rect 11529 54281 11563 54315
rect 22109 54281 22143 54315
rect 23213 54281 23247 54315
rect 34897 54281 34931 54315
rect 45109 54281 45143 54315
rect 1869 54213 1903 54247
rect 30389 54213 30423 54247
rect 52929 54213 52963 54247
rect 53573 54213 53607 54247
rect 28109 54145 28143 54179
rect 29377 54145 29411 54179
rect 29561 54145 29595 54179
rect 31401 54145 31435 54179
rect 32597 54145 32631 54179
rect 33241 54145 33275 54179
rect 33425 54145 33459 54179
rect 28365 54077 28399 54111
rect 32413 54077 32447 54111
rect 2053 54009 2087 54043
rect 53389 54009 53423 54043
rect 26985 53941 27019 53975
rect 28917 53941 28951 53975
rect 29469 53941 29503 53975
rect 30849 53941 30883 53975
rect 32781 53941 32815 53975
rect 33425 53941 33459 53975
rect 36093 53941 36127 53975
rect 1593 53737 1627 53771
rect 31401 53669 31435 53703
rect 33241 53669 33275 53703
rect 29561 53601 29595 53635
rect 30021 53601 30055 53635
rect 26893 53533 26927 53567
rect 28825 53533 28859 53567
rect 29009 53533 29043 53567
rect 29929 53533 29963 53567
rect 30573 53533 30607 53567
rect 30757 53533 30791 53567
rect 32781 53533 32815 53567
rect 27160 53465 27194 53499
rect 30665 53465 30699 53499
rect 32536 53465 32570 53499
rect 33609 53465 33643 53499
rect 52929 53465 52963 53499
rect 53573 53465 53607 53499
rect 24501 53397 24535 53431
rect 28273 53397 28307 53431
rect 28825 53397 28859 53431
rect 33425 53397 33459 53431
rect 33517 53397 33551 53431
rect 33793 53397 33827 53431
rect 53481 53397 53515 53431
rect 1409 53193 1443 53227
rect 24961 53193 24995 53227
rect 33701 53193 33735 53227
rect 34437 53193 34471 53227
rect 23857 53057 23891 53091
rect 24041 53057 24075 53091
rect 27905 53057 27939 53091
rect 31217 53057 31251 53091
rect 32137 53057 32171 53091
rect 33425 53057 33459 53091
rect 34345 53057 34379 53091
rect 34621 53057 34655 53091
rect 52929 53057 52963 53091
rect 53665 53057 53699 53091
rect 27997 52989 28031 53023
rect 28733 52989 28767 53023
rect 29009 52989 29043 53023
rect 31309 52989 31343 53023
rect 33517 52989 33551 53023
rect 33793 52989 33827 53023
rect 33885 52989 33919 53023
rect 30849 52921 30883 52955
rect 32597 52921 32631 52955
rect 23857 52853 23891 52887
rect 26249 52853 26283 52887
rect 26985 52853 27019 52887
rect 28273 52853 28307 52887
rect 30113 52853 30147 52887
rect 32229 52853 32263 52887
rect 33241 52853 33275 52887
rect 34805 52853 34839 52887
rect 35357 52853 35391 52887
rect 53481 52853 53515 52887
rect 29009 52649 29043 52683
rect 31493 52649 31527 52683
rect 1593 52581 1627 52615
rect 27997 52581 28031 52615
rect 32505 52581 32539 52615
rect 24409 52513 24443 52547
rect 24777 52513 24811 52547
rect 25605 52513 25639 52547
rect 26065 52513 26099 52547
rect 26617 52513 26651 52547
rect 29561 52513 29595 52547
rect 30021 52513 30055 52547
rect 31861 52513 31895 52547
rect 33333 52513 33367 52547
rect 34989 52513 35023 52547
rect 1409 52445 1443 52479
rect 23673 52445 23707 52479
rect 23857 52445 23891 52479
rect 24593 52445 24627 52479
rect 25697 52445 25731 52479
rect 26709 52445 26743 52479
rect 27537 52445 27571 52479
rect 27629 52445 27663 52479
rect 27813 52445 27847 52479
rect 28733 52445 28767 52479
rect 28825 52445 28859 52479
rect 29929 52445 29963 52479
rect 30205 52445 30239 52479
rect 30665 52445 30699 52479
rect 31033 52445 31067 52479
rect 31677 52445 31711 52479
rect 32413 52445 32447 52479
rect 32597 52445 32631 52479
rect 34161 52445 34195 52479
rect 35081 52445 35115 52479
rect 29009 52377 29043 52411
rect 30849 52377 30883 52411
rect 35725 52377 35759 52411
rect 23765 52309 23799 52343
rect 27077 52309 27111 52343
rect 34713 52309 34747 52343
rect 36277 52309 36311 52343
rect 1409 52105 1443 52139
rect 25145 52105 25179 52139
rect 26433 52105 26467 52139
rect 29837 52105 29871 52139
rect 31309 52105 31343 52139
rect 35357 52105 35391 52139
rect 36277 52105 36311 52139
rect 23765 52037 23799 52071
rect 29469 52037 29503 52071
rect 29653 52037 29687 52071
rect 30389 52037 30423 52071
rect 31493 52037 31527 52071
rect 33517 52037 33551 52071
rect 33609 52037 33643 52071
rect 23397 51969 23431 52003
rect 23581 51969 23615 52003
rect 23673 51969 23707 52003
rect 23857 51969 23891 52003
rect 24777 51969 24811 52003
rect 26249 51969 26283 52003
rect 27353 51969 27387 52003
rect 31217 51969 31251 52003
rect 32137 51969 32171 52003
rect 33379 51969 33413 52003
rect 33701 51969 33735 52003
rect 34529 51969 34563 52003
rect 35541 51969 35575 52003
rect 24685 51901 24719 51935
rect 26065 51901 26099 51935
rect 27629 51901 27663 51935
rect 33241 51901 33275 51935
rect 33885 51901 33919 51935
rect 34437 51901 34471 51935
rect 35725 51901 35759 51935
rect 35817 51901 35851 51935
rect 31493 51833 31527 51867
rect 22845 51765 22879 51799
rect 24041 51765 24075 51799
rect 28733 51765 28767 51799
rect 32781 51765 32815 51799
rect 34897 51765 34931 51799
rect 37289 51765 37323 51799
rect 22201 51561 22235 51595
rect 23213 51561 23247 51595
rect 26249 51561 26283 51595
rect 27629 51561 27663 51595
rect 35265 51561 35299 51595
rect 24869 51493 24903 51527
rect 36277 51493 36311 51527
rect 22753 51425 22787 51459
rect 26893 51425 26927 51459
rect 33333 51425 33367 51459
rect 23489 51357 23523 51391
rect 25513 51357 25547 51391
rect 25697 51357 25731 51391
rect 27353 51357 27387 51391
rect 27445 51357 27479 51391
rect 29009 51357 29043 51391
rect 30665 51357 30699 51391
rect 30849 51357 30883 51391
rect 31309 51357 31343 51391
rect 31493 51357 31527 51391
rect 33517 51357 33551 51391
rect 33793 51357 33827 51391
rect 34713 51357 34747 51391
rect 35081 51357 35115 51391
rect 23213 51289 23247 51323
rect 23397 51289 23431 51323
rect 27629 51289 27663 51323
rect 29561 51289 29595 51323
rect 30757 51289 30791 51323
rect 33701 51289 33735 51323
rect 34897 51289 34931 51323
rect 34989 51289 35023 51323
rect 25697 51221 25731 51255
rect 28089 51221 28123 51255
rect 30113 51221 30147 51255
rect 31401 51221 31435 51255
rect 31953 51221 31987 51255
rect 32597 51221 32631 51255
rect 35725 51221 35759 51255
rect 36921 51221 36955 51255
rect 23857 51017 23891 51051
rect 26157 51017 26191 51051
rect 31125 51017 31159 51051
rect 32873 51017 32907 51051
rect 35633 51017 35667 51051
rect 30021 50949 30055 50983
rect 30205 50949 30239 50983
rect 1409 50881 1443 50915
rect 22569 50881 22603 50915
rect 22753 50881 22787 50915
rect 23213 50881 23247 50915
rect 23397 50881 23431 50915
rect 23489 50881 23523 50915
rect 23581 50881 23615 50915
rect 25053 50881 25087 50915
rect 25881 50881 25915 50915
rect 30297 50881 30331 50915
rect 30941 50881 30975 50915
rect 32413 50881 32447 50915
rect 34897 50881 34931 50915
rect 52929 50881 52963 50915
rect 53573 50881 53607 50915
rect 24961 50813 24995 50847
rect 26157 50813 26191 50847
rect 30757 50813 30791 50847
rect 32137 50813 32171 50847
rect 34529 50813 34563 50847
rect 34989 50813 35023 50847
rect 25421 50745 25455 50779
rect 25973 50745 26007 50779
rect 28457 50745 28491 50779
rect 36185 50745 36219 50779
rect 1593 50677 1627 50711
rect 22017 50677 22051 50711
rect 22753 50677 22787 50711
rect 24317 50677 24351 50711
rect 27077 50677 27111 50711
rect 27997 50677 28031 50711
rect 29469 50677 29503 50711
rect 30021 50677 30055 50711
rect 32229 50677 32263 50711
rect 32321 50677 32355 50711
rect 33701 50677 33735 50711
rect 36737 50677 36771 50711
rect 53481 50677 53515 50711
rect 22845 50473 22879 50507
rect 23857 50473 23891 50507
rect 27169 50473 27203 50507
rect 30297 50473 30331 50507
rect 32689 50473 32723 50507
rect 34069 50473 34103 50507
rect 1409 50405 1443 50439
rect 31677 50405 31711 50439
rect 23397 50337 23431 50371
rect 25789 50337 25823 50371
rect 26249 50337 26283 50371
rect 28181 50337 28215 50371
rect 30389 50337 30423 50371
rect 20913 50269 20947 50303
rect 22477 50269 22511 50303
rect 22661 50269 22695 50303
rect 23489 50269 23523 50303
rect 25881 50269 25915 50303
rect 26709 50269 26743 50303
rect 26801 50269 26835 50303
rect 26985 50269 27019 50303
rect 30113 50269 30147 50303
rect 31125 50269 31159 50303
rect 31217 50269 31251 50303
rect 31401 50269 31435 50303
rect 31493 50269 31527 50303
rect 32505 50269 32539 50303
rect 32689 50269 32723 50303
rect 33149 50269 33183 50303
rect 33333 50269 33367 50303
rect 33517 50269 33551 50303
rect 34161 50269 34195 50303
rect 24869 50201 24903 50235
rect 25053 50201 25087 50235
rect 21465 50133 21499 50167
rect 22017 50133 22051 50167
rect 25237 50133 25271 50167
rect 28917 50133 28951 50167
rect 29929 50133 29963 50167
rect 32321 50133 32355 50167
rect 34713 50133 34747 50167
rect 35265 50133 35299 50167
rect 35909 50133 35943 50167
rect 22753 49929 22787 49963
rect 26433 49929 26467 49963
rect 31401 49929 31435 49963
rect 34253 49929 34287 49963
rect 35173 49929 35207 49963
rect 21281 49861 21315 49895
rect 22201 49861 22235 49895
rect 31033 49861 31067 49895
rect 34437 49861 34471 49895
rect 34621 49861 34655 49895
rect 22661 49793 22695 49827
rect 22845 49793 22879 49827
rect 23673 49793 23707 49827
rect 23857 49793 23891 49827
rect 24317 49793 24351 49827
rect 24501 49793 24535 49827
rect 25329 49793 25363 49827
rect 25513 49793 25547 49827
rect 26249 49793 26283 49827
rect 29754 49793 29788 49827
rect 30941 49793 30975 49827
rect 31217 49793 31251 49827
rect 32137 49793 32171 49827
rect 25421 49725 25455 49759
rect 26065 49725 26099 49759
rect 27077 49725 27111 49759
rect 28089 49725 28123 49759
rect 30021 49725 30055 49759
rect 32413 49725 32447 49759
rect 23765 49589 23799 49623
rect 24409 49589 24443 49623
rect 28641 49589 28675 49623
rect 33701 49589 33735 49623
rect 35633 49589 35667 49623
rect 36185 49589 36219 49623
rect 22293 49385 22327 49419
rect 29561 49385 29595 49419
rect 32689 49385 32723 49419
rect 36829 49385 36863 49419
rect 37289 49385 37323 49419
rect 23857 49317 23891 49351
rect 23581 49249 23615 49283
rect 30021 49249 30055 49283
rect 32505 49249 32539 49283
rect 33425 49249 33459 49283
rect 35633 49249 35667 49283
rect 23489 49181 23523 49215
rect 24409 49181 24443 49215
rect 24501 49181 24535 49215
rect 24685 49181 24719 49215
rect 25513 49181 25547 49215
rect 25973 49181 26007 49215
rect 26157 49181 26191 49215
rect 26801 49181 26835 49215
rect 27997 49181 28031 49215
rect 28181 49181 28215 49215
rect 28825 49181 28859 49215
rect 29009 49181 29043 49215
rect 29745 49181 29779 49215
rect 29929 49181 29963 49215
rect 30665 49181 30699 49215
rect 31309 49181 31343 49215
rect 31493 49181 31527 49215
rect 32321 49181 32355 49215
rect 32413 49181 32447 49215
rect 32689 49181 32723 49215
rect 33333 49181 33367 49215
rect 33517 49181 33551 49215
rect 33609 49181 33643 49215
rect 33793 49181 33827 49215
rect 34897 49181 34931 49215
rect 35541 49181 35575 49215
rect 35725 49181 35759 49215
rect 26617 49113 26651 49147
rect 26985 49113 27019 49147
rect 30481 49113 30515 49147
rect 30849 49113 30883 49147
rect 35081 49113 35115 49147
rect 21741 49045 21775 49079
rect 22845 49045 22879 49079
rect 24869 49045 24903 49079
rect 25421 49045 25455 49079
rect 26157 49045 26191 49079
rect 27537 49045 27571 49079
rect 28181 49045 28215 49079
rect 28825 49045 28859 49079
rect 31309 49045 31343 49079
rect 33149 49045 33183 49079
rect 34713 49045 34747 49079
rect 36185 49045 36219 49079
rect 23489 48841 23523 48875
rect 25329 48841 25363 48875
rect 34345 48841 34379 48875
rect 33517 48773 33551 48807
rect 34437 48773 34471 48807
rect 34621 48773 34655 48807
rect 21281 48705 21315 48739
rect 22477 48705 22511 48739
rect 23857 48705 23891 48739
rect 24685 48705 24719 48739
rect 24869 48705 24903 48739
rect 24961 48705 24995 48739
rect 25053 48705 25087 48739
rect 26249 48705 26283 48739
rect 26433 48705 26467 48739
rect 27169 48705 27203 48739
rect 28549 48705 28583 48739
rect 30113 48705 30147 48739
rect 30205 48705 30239 48739
rect 30389 48705 30423 48739
rect 30849 48705 30883 48739
rect 31033 48705 31067 48739
rect 33701 48705 33735 48739
rect 34345 48705 34379 48739
rect 35081 48705 35115 48739
rect 35265 48705 35299 48739
rect 52929 48705 52963 48739
rect 53573 48705 53607 48739
rect 23673 48637 23707 48671
rect 23765 48637 23799 48671
rect 23949 48637 23983 48671
rect 27261 48637 27295 48671
rect 28457 48637 28491 48671
rect 21925 48569 21959 48603
rect 22937 48569 22971 48603
rect 27537 48569 27571 48603
rect 28917 48569 28951 48603
rect 32689 48569 32723 48603
rect 35173 48569 35207 48603
rect 53389 48569 53423 48603
rect 26341 48501 26375 48535
rect 29377 48501 29411 48535
rect 30113 48501 30147 48535
rect 30941 48501 30975 48535
rect 31493 48501 31527 48535
rect 32229 48501 32263 48535
rect 33885 48501 33919 48535
rect 35725 48501 35759 48535
rect 36369 48501 36403 48535
rect 24961 48297 24995 48331
rect 29745 48297 29779 48331
rect 21833 48229 21867 48263
rect 23857 48229 23891 48263
rect 26709 48229 26743 48263
rect 27169 48229 27203 48263
rect 29009 48229 29043 48263
rect 36093 48229 36127 48263
rect 26433 48161 26467 48195
rect 29929 48161 29963 48195
rect 30021 48161 30055 48195
rect 30757 48161 30791 48195
rect 32689 48161 32723 48195
rect 33609 48161 33643 48195
rect 34805 48161 34839 48195
rect 34989 48161 35023 48195
rect 35541 48161 35575 48195
rect 37289 48161 37323 48195
rect 1685 48093 1719 48127
rect 21189 48093 21223 48127
rect 24501 48093 24535 48127
rect 24777 48093 24811 48127
rect 25421 48093 25455 48127
rect 25605 48093 25639 48127
rect 26341 48093 26375 48127
rect 27307 48093 27341 48127
rect 27537 48093 27571 48127
rect 27720 48093 27754 48127
rect 27813 48093 27847 48127
rect 28365 48093 28399 48127
rect 28549 48093 28583 48127
rect 28641 48093 28675 48127
rect 30113 48093 30147 48127
rect 30205 48093 30239 48127
rect 30941 48093 30975 48127
rect 31125 48093 31159 48127
rect 31217 48093 31251 48127
rect 32229 48093 32263 48127
rect 32321 48093 32355 48127
rect 32505 48093 32539 48127
rect 33517 48093 33551 48127
rect 34713 48093 34747 48127
rect 35449 48093 35483 48127
rect 35633 48093 35667 48127
rect 2237 48025 2271 48059
rect 24593 48025 24627 48059
rect 27445 48025 27479 48059
rect 1501 47957 1535 47991
rect 20729 47957 20763 47991
rect 22293 47957 22327 47991
rect 22937 47957 22971 47991
rect 25605 47957 25639 47991
rect 31677 47957 31711 47991
rect 33149 47957 33183 47991
rect 34989 47957 35023 47991
rect 36645 47957 36679 47991
rect 23489 47753 23523 47787
rect 24041 47753 24075 47787
rect 24593 47753 24627 47787
rect 26433 47753 26467 47787
rect 29009 47753 29043 47787
rect 30573 47753 30607 47787
rect 31217 47753 31251 47787
rect 35265 47753 35299 47787
rect 25329 47685 25363 47719
rect 25513 47685 25547 47719
rect 27721 47685 27755 47719
rect 29285 47685 29319 47719
rect 22293 47617 22327 47651
rect 23305 47617 23339 47651
rect 24501 47617 24535 47651
rect 24685 47617 24719 47651
rect 25145 47617 25179 47651
rect 26065 47617 26099 47651
rect 26249 47617 26283 47651
rect 26985 47617 27019 47651
rect 27261 47617 27295 47651
rect 27537 47617 27571 47651
rect 29188 47617 29222 47651
rect 29377 47617 29411 47651
rect 29560 47617 29594 47651
rect 29653 47617 29687 47651
rect 31033 47617 31067 47651
rect 32137 47617 32171 47651
rect 32321 47617 32355 47651
rect 32965 47617 32999 47651
rect 33149 47617 33183 47651
rect 33241 47617 33275 47651
rect 33425 47617 33459 47651
rect 34529 47617 34563 47651
rect 35173 47617 35207 47651
rect 35357 47617 35391 47651
rect 22385 47549 22419 47583
rect 23121 47549 23155 47583
rect 25973 47549 26007 47583
rect 30941 47549 30975 47583
rect 32229 47549 32263 47583
rect 33333 47549 33367 47583
rect 34621 47549 34655 47583
rect 22661 47481 22695 47515
rect 27813 47481 27847 47515
rect 34161 47481 34195 47515
rect 36369 47481 36403 47515
rect 20177 47413 20211 47447
rect 20729 47413 20763 47447
rect 21281 47413 21315 47447
rect 28549 47413 28583 47447
rect 33701 47413 33735 47447
rect 35817 47413 35851 47447
rect 37381 47413 37415 47447
rect 26709 47209 26743 47243
rect 28641 47209 28675 47243
rect 30297 47209 30331 47243
rect 30757 47209 30791 47243
rect 32965 47209 32999 47243
rect 34161 47209 34195 47243
rect 23581 47141 23615 47175
rect 27169 47141 27203 47175
rect 35357 47141 35391 47175
rect 23305 47073 23339 47107
rect 24501 47073 24535 47107
rect 28181 47073 28215 47107
rect 29837 47073 29871 47107
rect 32505 47073 32539 47107
rect 37473 47073 37507 47107
rect 20269 47005 20303 47039
rect 23213 47005 23247 47039
rect 24961 47005 24995 47039
rect 25145 47005 25179 47039
rect 25237 47005 25271 47039
rect 25329 47005 25363 47039
rect 26065 47005 26099 47039
rect 26249 47005 26283 47039
rect 26341 47005 26375 47039
rect 26433 47005 26467 47039
rect 27169 47005 27203 47039
rect 27445 47005 27479 47039
rect 28825 47005 28859 47039
rect 29929 47005 29963 47039
rect 30113 47005 30147 47039
rect 31125 47005 31159 47039
rect 32229 47005 32263 47039
rect 32321 47005 32355 47039
rect 33144 47005 33178 47039
rect 33461 47005 33495 47039
rect 33584 47005 33618 47039
rect 36921 47005 36955 47039
rect 20729 46937 20763 46971
rect 21373 46937 21407 46971
rect 25605 46937 25639 46971
rect 27353 46937 27387 46971
rect 29009 46937 29043 46971
rect 30941 46937 30975 46971
rect 31677 46937 31711 46971
rect 33241 46937 33275 46971
rect 33333 46937 33367 46971
rect 34713 46937 34747 46971
rect 35909 46937 35943 46971
rect 19625 46869 19659 46903
rect 21833 46869 21867 46903
rect 22385 46869 22419 46903
rect 32505 46869 32539 46903
rect 36461 46869 36495 46903
rect 21281 46665 21315 46699
rect 23581 46665 23615 46699
rect 24593 46665 24627 46699
rect 25513 46665 25547 46699
rect 29193 46665 29227 46699
rect 30021 46665 30055 46699
rect 30757 46665 30791 46699
rect 31309 46665 31343 46699
rect 32689 46665 32723 46699
rect 34069 46665 34103 46699
rect 28825 46597 28859 46631
rect 29041 46597 29075 46631
rect 29929 46597 29963 46631
rect 33149 46597 33183 46631
rect 34621 46597 34655 46631
rect 23397 46529 23431 46563
rect 23581 46529 23615 46563
rect 24225 46529 24259 46563
rect 25697 46529 25731 46563
rect 25881 46529 25915 46563
rect 26985 46529 27019 46563
rect 27261 46529 27295 46563
rect 29653 46529 29687 46563
rect 29837 46529 29871 46563
rect 30665 46529 30699 46563
rect 30849 46529 30883 46563
rect 32321 46529 32355 46563
rect 33333 46529 33367 46563
rect 33609 46529 33643 46563
rect 34805 46529 34839 46563
rect 36001 46529 36035 46563
rect 53389 46529 53423 46563
rect 20729 46461 20763 46495
rect 24317 46461 24351 46495
rect 25789 46461 25823 46495
rect 25973 46461 26007 46495
rect 30205 46461 30239 46495
rect 32229 46461 32263 46495
rect 33517 46461 33551 46495
rect 35541 46461 35575 46495
rect 52837 46461 52871 46495
rect 22845 46393 22879 46427
rect 18889 46325 18923 46359
rect 19349 46325 19383 46359
rect 19993 46325 20027 46359
rect 22385 46325 22419 46359
rect 27077 46325 27111 46359
rect 27445 46325 27479 46359
rect 28273 46325 28307 46359
rect 29009 46325 29043 46359
rect 34989 46325 35023 46359
rect 36645 46325 36679 46359
rect 37289 46325 37323 46359
rect 37841 46325 37875 46359
rect 53573 46325 53607 46359
rect 18705 46121 18739 46155
rect 21005 46121 21039 46155
rect 23213 46121 23247 46155
rect 25605 46121 25639 46155
rect 29561 46121 29595 46155
rect 32321 46121 32355 46155
rect 32965 46121 32999 46155
rect 33149 46121 33183 46155
rect 35173 46053 35207 46087
rect 22201 45985 22235 46019
rect 27997 45985 28031 46019
rect 33241 45985 33275 46019
rect 20177 45917 20211 45951
rect 20361 45917 20395 45951
rect 21649 45917 21683 45951
rect 25513 45917 25547 45951
rect 25697 45917 25731 45951
rect 27730 45917 27764 45951
rect 29745 45917 29779 45951
rect 29837 45917 29871 45951
rect 30389 45917 30423 45951
rect 33333 45917 33367 45951
rect 34069 45917 34103 45951
rect 34161 45917 34195 45951
rect 34713 45917 34747 45951
rect 34989 45917 35023 45951
rect 35633 45917 35667 45951
rect 35817 45917 35851 45951
rect 36277 45917 36311 45951
rect 37381 45917 37415 45951
rect 1869 45849 1903 45883
rect 2053 45849 2087 45883
rect 19717 45849 19751 45883
rect 23857 45849 23891 45883
rect 29561 45849 29595 45883
rect 32137 45849 32171 45883
rect 32337 45849 32371 45883
rect 33885 45849 33919 45883
rect 17509 45781 17543 45815
rect 20269 45781 20303 45815
rect 22753 45781 22787 45815
rect 24501 45781 24535 45815
rect 25053 45781 25087 45815
rect 26617 45781 26651 45815
rect 28457 45781 28491 45815
rect 30849 45781 30883 45815
rect 31493 45781 31527 45815
rect 32505 45781 32539 45815
rect 33977 45781 34011 45815
rect 34805 45781 34839 45815
rect 35817 45781 35851 45815
rect 36921 45781 36955 45815
rect 1593 45577 1627 45611
rect 20085 45577 20119 45611
rect 22477 45577 22511 45611
rect 27445 45577 27479 45611
rect 30297 45577 30331 45611
rect 31217 45577 31251 45611
rect 32321 45577 32355 45611
rect 33625 45577 33659 45611
rect 34437 45577 34471 45611
rect 34621 45577 34655 45611
rect 35449 45577 35483 45611
rect 19441 45509 19475 45543
rect 25789 45509 25823 45543
rect 26341 45509 26375 45543
rect 29101 45509 29135 45543
rect 32505 45509 32539 45543
rect 33425 45509 33459 45543
rect 36277 45509 36311 45543
rect 19349 45441 19383 45475
rect 19533 45441 19567 45475
rect 19993 45441 20027 45475
rect 20269 45441 20303 45475
rect 20729 45441 20763 45475
rect 20913 45441 20947 45475
rect 22937 45441 22971 45475
rect 23121 45441 23155 45475
rect 23581 45441 23615 45475
rect 27261 45441 27295 45475
rect 32229 45441 32263 45475
rect 34713 45441 34747 45475
rect 35633 45441 35667 45475
rect 17785 45373 17819 45407
rect 23029 45373 23063 45407
rect 23857 45373 23891 45407
rect 25329 45373 25363 45407
rect 34345 45373 34379 45407
rect 34805 45373 34839 45407
rect 35817 45373 35851 45407
rect 18337 45305 18371 45339
rect 20269 45305 20303 45339
rect 32505 45305 32539 45339
rect 33793 45305 33827 45339
rect 37841 45305 37875 45339
rect 17233 45237 17267 45271
rect 18889 45237 18923 45271
rect 20821 45237 20855 45271
rect 21925 45237 21959 45271
rect 23673 45237 23707 45271
rect 23765 45237 23799 45271
rect 24777 45237 24811 45271
rect 27997 45237 28031 45271
rect 28549 45237 28583 45271
rect 29653 45237 29687 45271
rect 33609 45237 33643 45271
rect 34989 45237 35023 45271
rect 37381 45237 37415 45271
rect 16497 45033 16531 45067
rect 19257 45033 19291 45067
rect 22753 45033 22787 45067
rect 30941 45033 30975 45067
rect 31953 45033 31987 45067
rect 36001 45033 36035 45067
rect 37841 45033 37875 45067
rect 17233 44965 17267 44999
rect 18705 44965 18739 44999
rect 21189 44965 21223 44999
rect 23857 44965 23891 44999
rect 24501 44965 24535 44999
rect 25421 44965 25455 44999
rect 26985 44965 27019 44999
rect 29009 44965 29043 44999
rect 19809 44897 19843 44931
rect 20913 44897 20947 44931
rect 23397 44897 23431 44931
rect 24961 44897 24995 44931
rect 29561 44897 29595 44931
rect 33609 44897 33643 44931
rect 34713 44897 34747 44931
rect 34989 44897 35023 44931
rect 35173 44897 35207 44931
rect 36737 44897 36771 44931
rect 16957 44829 16991 44863
rect 17693 44829 17727 44863
rect 17877 44829 17911 44863
rect 19993 44829 20027 44863
rect 20821 44829 20855 44863
rect 21649 44829 21683 44863
rect 21833 44829 21867 44863
rect 22385 44829 22419 44863
rect 22569 44829 22603 44863
rect 23567 44829 23601 44863
rect 24409 44829 24443 44863
rect 24685 44829 24719 44863
rect 24777 44829 24811 44863
rect 25697 44829 25731 44863
rect 27261 44829 27295 44863
rect 28733 44829 28767 44863
rect 29837 44829 29871 44863
rect 31953 44829 31987 44863
rect 32597 44829 32631 44863
rect 32781 44829 32815 44863
rect 33425 44829 33459 44863
rect 33701 44829 33735 44863
rect 34897 44829 34931 44863
rect 35081 44829 35115 44863
rect 35725 44829 35759 44863
rect 36185 44829 36219 44863
rect 36645 44829 36679 44863
rect 36829 44829 36863 44863
rect 17233 44761 17267 44795
rect 25421 44761 25455 44795
rect 26433 44761 26467 44795
rect 26985 44761 27019 44795
rect 29009 44761 29043 44795
rect 35817 44761 35851 44795
rect 37289 44761 37323 44795
rect 38393 44761 38427 44795
rect 15301 44693 15335 44727
rect 15853 44693 15887 44727
rect 17049 44693 17083 44727
rect 17877 44693 17911 44727
rect 20177 44693 20211 44727
rect 21741 44693 21775 44727
rect 25605 44693 25639 44727
rect 27169 44693 27203 44727
rect 28181 44693 28215 44727
rect 28825 44693 28859 44727
rect 32689 44693 32723 44727
rect 33241 44693 33275 44727
rect 38945 44693 38979 44727
rect 19365 44489 19399 44523
rect 22033 44489 22067 44523
rect 25145 44489 25179 44523
rect 26433 44489 26467 44523
rect 30849 44489 30883 44523
rect 33517 44489 33551 44523
rect 34345 44489 34379 44523
rect 35357 44489 35391 44523
rect 36185 44489 36219 44523
rect 37289 44489 37323 44523
rect 18705 44421 18739 44455
rect 19165 44421 19199 44455
rect 20085 44421 20119 44455
rect 20269 44421 20303 44455
rect 20913 44421 20947 44455
rect 21833 44421 21867 44455
rect 22753 44421 22787 44455
rect 23305 44421 23339 44455
rect 28641 44421 28675 44455
rect 31217 44421 31251 44455
rect 34161 44421 34195 44455
rect 15577 44353 15611 44387
rect 15761 44353 15795 44387
rect 16681 44353 16715 44387
rect 16865 44353 16899 44387
rect 17325 44353 17359 44387
rect 17509 44353 17543 44387
rect 18429 44353 18463 44387
rect 18521 44353 18555 44387
rect 21097 44353 21131 44387
rect 22661 44353 22695 44387
rect 22845 44353 22879 44387
rect 23489 44353 23523 44387
rect 24317 44353 24351 44387
rect 25329 44353 25363 44387
rect 25513 44353 25547 44387
rect 25605 44353 25639 44387
rect 26065 44353 26099 44387
rect 26249 44353 26283 44387
rect 27721 44353 27755 44387
rect 30389 44353 30423 44387
rect 31033 44353 31067 44387
rect 31309 44353 31343 44387
rect 32137 44353 32171 44387
rect 32321 44353 32355 44387
rect 32781 44353 32815 44387
rect 32965 44353 32999 44387
rect 33057 44353 33091 44387
rect 33333 44353 33367 44387
rect 34437 44353 34471 44387
rect 35541 44353 35575 44387
rect 36369 44353 36403 44387
rect 36553 44353 36587 44387
rect 24225 44285 24259 44319
rect 24685 44285 24719 44319
rect 27997 44285 28031 44319
rect 32229 44285 32263 44319
rect 33149 44285 33183 44319
rect 35725 44285 35759 44319
rect 15669 44217 15703 44251
rect 18705 44217 18739 44251
rect 19533 44217 19567 44251
rect 22201 44217 22235 44251
rect 27905 44217 27939 44251
rect 34161 44217 34195 44251
rect 38393 44217 38427 44251
rect 13737 44149 13771 44183
rect 14473 44149 14507 44183
rect 15025 44149 15059 44183
rect 16865 44149 16899 44183
rect 17693 44149 17727 44183
rect 19349 44149 19383 44183
rect 20453 44149 20487 44183
rect 21281 44149 21315 44183
rect 22017 44149 22051 44183
rect 23673 44149 23707 44183
rect 27169 44149 27203 44183
rect 27813 44149 27847 44183
rect 37841 44149 37875 44183
rect 39037 44149 39071 44183
rect 13461 43945 13495 43979
rect 17417 43945 17451 43979
rect 18429 43945 18463 43979
rect 21189 43945 21223 43979
rect 23857 43945 23891 43979
rect 25145 43945 25179 43979
rect 28365 43945 28399 43979
rect 32873 43945 32907 43979
rect 33425 43945 33459 43979
rect 35265 43945 35299 43979
rect 36369 43945 36403 43979
rect 15669 43877 15703 43911
rect 20453 43877 20487 43911
rect 22017 43877 22051 43911
rect 26249 43877 26283 43911
rect 37933 43877 37967 43911
rect 17233 43809 17267 43843
rect 22569 43809 22603 43843
rect 23765 43809 23799 43843
rect 25053 43809 25087 43843
rect 25513 43809 25547 43843
rect 26985 43809 27019 43843
rect 29561 43809 29595 43843
rect 33793 43809 33827 43843
rect 35909 43809 35943 43843
rect 2053 43741 2087 43775
rect 14749 43741 14783 43775
rect 14933 43741 14967 43775
rect 15393 43741 15427 43775
rect 15485 43741 15519 43775
rect 15669 43741 15703 43775
rect 17141 43741 17175 43775
rect 17969 43741 18003 43775
rect 18245 43741 18279 43775
rect 19533 43741 19567 43775
rect 20453 43741 20487 43775
rect 20729 43741 20763 43775
rect 21189 43741 21223 43775
rect 21465 43741 21499 43775
rect 21925 43741 21959 43775
rect 22109 43741 22143 43775
rect 22753 43741 22787 43775
rect 23581 43741 23615 43775
rect 25329 43741 25363 43775
rect 26065 43741 26099 43775
rect 26157 43741 26191 43775
rect 26341 43741 26375 43775
rect 26525 43741 26559 43775
rect 27261 43741 27295 43775
rect 29817 43741 29851 43775
rect 31493 43741 31527 43775
rect 31760 43741 31794 43775
rect 33609 43741 33643 43775
rect 36001 43741 36035 43775
rect 53389 43741 53423 43775
rect 1869 43673 1903 43707
rect 16129 43673 16163 43707
rect 16313 43673 16347 43707
rect 18061 43673 18095 43707
rect 19625 43673 19659 43707
rect 19809 43673 19843 43707
rect 20637 43673 20671 43707
rect 22937 43673 22971 43707
rect 23857 43673 23891 43707
rect 34713 43673 34747 43707
rect 37473 43673 37507 43707
rect 14197 43605 14231 43639
rect 14933 43605 14967 43639
rect 16497 43605 16531 43639
rect 19717 43605 19751 43639
rect 21373 43605 21407 43639
rect 23397 43605 23431 43639
rect 24409 43605 24443 43639
rect 30941 43605 30975 43639
rect 36829 43605 36863 43639
rect 38577 43605 38611 43639
rect 39129 43605 39163 43639
rect 52837 43605 52871 43639
rect 53573 43605 53607 43639
rect 1593 43401 1627 43435
rect 14473 43401 14507 43435
rect 14933 43401 14967 43435
rect 18521 43401 18555 43435
rect 19533 43401 19567 43435
rect 25789 43401 25823 43435
rect 27721 43401 27755 43435
rect 30113 43401 30147 43435
rect 31033 43401 31067 43435
rect 14105 43333 14139 43367
rect 18797 43333 18831 43367
rect 20821 43333 20855 43367
rect 22753 43333 22787 43367
rect 24501 43333 24535 43367
rect 30849 43333 30883 43367
rect 31401 43333 31435 43367
rect 34897 43333 34931 43367
rect 36461 43333 36495 43367
rect 37289 43333 37323 43367
rect 37841 43333 37875 43367
rect 38393 43333 38427 43367
rect 13093 43265 13127 43299
rect 13645 43265 13679 43299
rect 14289 43265 14323 43299
rect 15393 43265 15427 43299
rect 16865 43265 16899 43299
rect 16957 43265 16991 43299
rect 17141 43265 17175 43299
rect 17233 43265 17267 43299
rect 17877 43265 17911 43299
rect 18521 43265 18555 43299
rect 18613 43265 18647 43299
rect 19441 43265 19475 43299
rect 19717 43265 19751 43299
rect 21925 43265 21959 43299
rect 22109 43265 22143 43299
rect 22569 43265 22603 43299
rect 23397 43265 23431 43299
rect 23581 43265 23615 43299
rect 23673 43265 23707 43299
rect 23765 43265 23799 43299
rect 24777 43265 24811 43299
rect 25605 43265 25639 43299
rect 27077 43265 27111 43299
rect 27537 43265 27571 43299
rect 28641 43265 28675 43299
rect 31125 43265 31159 43299
rect 31217 43265 31251 43299
rect 32689 43265 32723 43299
rect 33793 43265 33827 43299
rect 34253 43265 34287 43299
rect 34437 43265 34471 43299
rect 35541 43265 35575 43299
rect 35725 43265 35759 43299
rect 36185 43265 36219 43299
rect 36277 43265 36311 43299
rect 15301 43197 15335 43231
rect 16129 43197 16163 43231
rect 17693 43197 17727 43231
rect 18061 43197 18095 43231
rect 22017 43197 22051 43231
rect 24593 43197 24627 43231
rect 25421 43197 25455 43231
rect 27261 43197 27295 43231
rect 27353 43197 27387 43231
rect 32781 43197 32815 43231
rect 33057 43197 33091 43231
rect 33517 43197 33551 43231
rect 35633 43197 35667 43231
rect 15577 43129 15611 43163
rect 21189 43129 21223 43163
rect 27445 43129 27479 43163
rect 33701 43129 33735 43163
rect 16681 43061 16715 43095
rect 19901 43061 19935 43095
rect 21281 43061 21315 43095
rect 22937 43061 22971 43095
rect 24041 43061 24075 43095
rect 24777 43061 24811 43095
rect 24961 43061 24995 43095
rect 26433 43061 26467 43095
rect 33609 43061 33643 43095
rect 34345 43061 34379 43095
rect 36461 43061 36495 43095
rect 38945 43061 38979 43095
rect 39497 43061 39531 43095
rect 40049 43061 40083 43095
rect 13001 42857 13035 42891
rect 14197 42857 14231 42891
rect 17693 42857 17727 42891
rect 18613 42857 18647 42891
rect 21281 42857 21315 42891
rect 28457 42857 28491 42891
rect 28649 42857 28683 42891
rect 32137 42857 32171 42891
rect 35541 42857 35575 42891
rect 36001 42857 36035 42891
rect 16957 42789 16991 42823
rect 23581 42789 23615 42823
rect 27261 42789 27295 42823
rect 34069 42789 34103 42823
rect 38301 42789 38335 42823
rect 15117 42721 15151 42755
rect 16865 42721 16899 42755
rect 19349 42721 19383 42755
rect 20913 42721 20947 42755
rect 21833 42721 21867 42755
rect 23029 42721 23063 42755
rect 25329 42721 25363 42755
rect 29745 42721 29779 42755
rect 29929 42721 29963 42755
rect 36369 42721 36403 42755
rect 38853 42721 38887 42755
rect 14105 42653 14139 42687
rect 14289 42653 14323 42687
rect 15761 42653 15795 42687
rect 16037 42653 16071 42687
rect 16773 42653 16807 42687
rect 17049 42653 17083 42687
rect 17693 42653 17727 42687
rect 17785 42653 17819 42687
rect 19901 42653 19935 42687
rect 20361 42653 20395 42687
rect 21005 42653 21039 42687
rect 22937 42653 22971 42687
rect 23121 42653 23155 42687
rect 23581 42653 23615 42687
rect 23857 42653 23891 42687
rect 24593 42653 24627 42687
rect 24777 42653 24811 42687
rect 25237 42653 25271 42687
rect 25421 42653 25455 42687
rect 26801 42653 26835 42687
rect 27813 42653 27847 42687
rect 29009 42653 29043 42687
rect 29837 42653 29871 42687
rect 30021 42653 30055 42687
rect 32045 42653 32079 42687
rect 32229 42653 32263 42687
rect 32873 42653 32907 42687
rect 33057 42653 33091 42687
rect 33793 42653 33827 42687
rect 34713 42653 34747 42687
rect 34897 42653 34931 42687
rect 35357 42653 35391 42687
rect 35541 42653 35575 42687
rect 36185 42653 36219 42687
rect 36921 42653 36955 42687
rect 37013 42655 37047 42689
rect 37197 42653 37231 42687
rect 37657 42653 37691 42687
rect 37841 42653 37875 42687
rect 14749 42585 14783 42619
rect 14933 42585 14967 42619
rect 16221 42585 16255 42619
rect 20269 42585 20303 42619
rect 23765 42585 23799 42619
rect 24409 42585 24443 42619
rect 27629 42585 27663 42619
rect 31125 42585 31159 42619
rect 32689 42585 32723 42619
rect 34069 42585 34103 42619
rect 40417 42585 40451 42619
rect 13553 42517 13587 42551
rect 15853 42517 15887 42551
rect 17233 42517 17267 42551
rect 18061 42517 18095 42551
rect 20177 42517 20211 42551
rect 22385 42517 22419 42551
rect 26249 42517 26283 42551
rect 27445 42517 27479 42551
rect 27537 42517 27571 42551
rect 28641 42517 28675 42551
rect 29561 42517 29595 42551
rect 30573 42517 30607 42551
rect 33885 42517 33919 42551
rect 34713 42517 34747 42551
rect 37749 42517 37783 42551
rect 39957 42517 39991 42551
rect 40969 42517 41003 42551
rect 14933 42313 14967 42347
rect 17049 42313 17083 42347
rect 17601 42313 17635 42347
rect 19809 42313 19843 42347
rect 22109 42313 22143 42347
rect 22385 42313 22419 42347
rect 23397 42313 23431 42347
rect 24593 42313 24627 42347
rect 26341 42313 26375 42347
rect 27813 42313 27847 42347
rect 27981 42313 28015 42347
rect 29561 42313 29595 42347
rect 31401 42313 31435 42347
rect 34989 42313 35023 42347
rect 35157 42313 35191 42347
rect 36461 42313 36495 42347
rect 39405 42313 39439 42347
rect 40509 42313 40543 42347
rect 15853 42245 15887 42279
rect 16037 42245 16071 42279
rect 18981 42245 19015 42279
rect 22201 42245 22235 42279
rect 23949 42245 23983 42279
rect 28181 42245 28215 42279
rect 28825 42245 28859 42279
rect 35357 42245 35391 42279
rect 37381 42245 37415 42279
rect 41061 42245 41095 42279
rect 14749 42177 14783 42211
rect 14933 42177 14967 42211
rect 16129 42177 16163 42211
rect 16681 42177 16715 42211
rect 16865 42177 16899 42211
rect 17509 42177 17543 42211
rect 17693 42177 17727 42211
rect 19625 42177 19659 42211
rect 20453 42177 20487 42211
rect 20729 42177 20763 42211
rect 20913 42177 20947 42211
rect 22017 42177 22051 42211
rect 23213 42177 23247 42211
rect 23397 42177 23431 42211
rect 24409 42177 24443 42211
rect 24593 42177 24627 42211
rect 27169 42177 27203 42211
rect 27353 42177 27387 42211
rect 28641 42177 28675 42211
rect 28917 42177 28951 42211
rect 30674 42177 30708 42211
rect 30941 42177 30975 42211
rect 32137 42177 32171 42211
rect 33149 42177 33183 42211
rect 34069 42177 34103 42211
rect 34345 42177 34379 42211
rect 35909 42177 35943 42211
rect 36093 42177 36127 42211
rect 36185 42177 36219 42211
rect 36277 42177 36311 42211
rect 37289 42177 37323 42211
rect 37565 42177 37599 42211
rect 38393 42177 38427 42211
rect 14289 42109 14323 42143
rect 19441 42109 19475 42143
rect 25237 42109 25271 42143
rect 33241 42109 33275 42143
rect 34161 42109 34195 42143
rect 38853 42109 38887 42143
rect 16129 42041 16163 42075
rect 21833 42041 21867 42075
rect 25881 42041 25915 42075
rect 28641 42041 28675 42075
rect 33517 42041 33551 42075
rect 34253 42041 34287 42075
rect 38301 42041 38335 42075
rect 41613 42041 41647 42075
rect 13645 41973 13679 42007
rect 18429 41973 18463 42007
rect 20269 41973 20303 42007
rect 27353 41973 27387 42007
rect 27997 41973 28031 42007
rect 32321 41973 32355 42007
rect 34529 41973 34563 42007
rect 35173 41973 35207 42007
rect 37749 41973 37783 42007
rect 40049 41973 40083 42007
rect 14381 41769 14415 41803
rect 17601 41769 17635 41803
rect 19717 41769 19751 41803
rect 30389 41769 30423 41803
rect 33517 41769 33551 41803
rect 35633 41769 35667 41803
rect 38945 41769 38979 41803
rect 39957 41769 39991 41803
rect 41521 41769 41555 41803
rect 22201 41701 22235 41735
rect 27261 41701 27295 41735
rect 37657 41701 37691 41735
rect 15485 41633 15519 41667
rect 16589 41633 16623 41667
rect 21741 41633 21775 41667
rect 25053 41633 25087 41667
rect 32137 41633 32171 41667
rect 36369 41633 36403 41667
rect 17785 41565 17819 41599
rect 17969 41565 18003 41599
rect 18061 41565 18095 41599
rect 20269 41565 20303 41599
rect 20453 41565 20487 41599
rect 20637 41565 20671 41599
rect 21005 41565 21039 41599
rect 21189 41565 21223 41599
rect 21833 41565 21867 41599
rect 23489 41565 23523 41599
rect 24869 41565 24903 41599
rect 25513 41565 25547 41599
rect 25697 41565 25731 41599
rect 26985 41565 27019 41599
rect 27077 41565 27111 41599
rect 27353 41565 27387 41599
rect 27813 41565 27847 41599
rect 27997 41565 28031 41599
rect 31677 41565 31711 41599
rect 32404 41565 32438 41599
rect 34713 41565 34747 41599
rect 34897 41565 34931 41599
rect 36461 41565 36495 41599
rect 37289 41565 37323 41599
rect 38485 41565 38519 41599
rect 38945 41565 38979 41599
rect 39129 41565 39163 41599
rect 17141 41497 17175 41531
rect 22937 41497 22971 41531
rect 24685 41497 24719 41531
rect 25881 41497 25915 41531
rect 27905 41497 27939 41531
rect 29009 41497 29043 41531
rect 34069 41497 34103 41531
rect 37473 41497 37507 41531
rect 38301 41497 38335 41531
rect 53389 41497 53423 41531
rect 53573 41497 53607 41531
rect 16037 41429 16071 41463
rect 18705 41429 18739 41463
rect 20177 41429 20211 41463
rect 26801 41429 26835 41463
rect 35081 41429 35115 41463
rect 36093 41429 36127 41463
rect 37105 41429 37139 41463
rect 37381 41429 37415 41463
rect 38117 41429 38151 41463
rect 40509 41429 40543 41463
rect 41061 41429 41095 41463
rect 42073 41429 42107 41463
rect 42625 41429 42659 41463
rect 52929 41429 52963 41463
rect 16037 41225 16071 41259
rect 17877 41225 17911 41259
rect 25237 41225 25271 41259
rect 28365 41225 28399 41259
rect 30297 41225 30331 41259
rect 32229 41225 32263 41259
rect 36645 41225 36679 41259
rect 38025 41225 38059 41259
rect 38393 41225 38427 41259
rect 40969 41225 41003 41259
rect 30757 41157 30791 41191
rect 33517 41157 33551 41191
rect 33635 41157 33669 41191
rect 41521 41157 41555 41191
rect 1685 41089 1719 41123
rect 17693 41089 17727 41123
rect 17969 41089 18003 41123
rect 18613 41089 18647 41123
rect 19717 41089 19751 41123
rect 21281 41089 21315 41123
rect 22661 41089 22695 41123
rect 23673 41089 23707 41123
rect 23857 41089 23891 41123
rect 24593 41089 24627 41123
rect 25053 41089 25087 41123
rect 25237 41089 25271 41123
rect 29561 41089 29595 41123
rect 29745 41095 29779 41129
rect 30124 41089 30158 41123
rect 30941 41089 30975 41123
rect 31033 41089 31067 41123
rect 31309 41089 31343 41123
rect 32413 41089 32447 41123
rect 32597 41089 32631 41123
rect 33333 41089 33367 41123
rect 33425 41089 33459 41123
rect 34437 41089 34471 41123
rect 34621 41089 34655 41123
rect 35633 41089 35667 41123
rect 36461 41089 36495 41123
rect 36737 41089 36771 41123
rect 37749 41089 37783 41123
rect 38117 41089 38151 41123
rect 39037 41089 39071 41123
rect 39129 41089 39163 41123
rect 39313 41089 39347 41123
rect 39405 41089 39439 41123
rect 18429 41021 18463 41055
rect 20637 41021 20671 41055
rect 24317 41021 24351 41055
rect 26985 41021 27019 41055
rect 27261 41021 27295 41055
rect 29837 41021 29871 41055
rect 29929 41021 29963 41055
rect 33793 41021 33827 41055
rect 35449 41021 35483 41055
rect 38234 41021 38268 41055
rect 39865 41021 39899 41055
rect 2237 40953 2271 40987
rect 17049 40953 17083 40987
rect 18797 40953 18831 40987
rect 22017 40953 22051 40987
rect 25881 40953 25915 40987
rect 38853 40953 38887 40987
rect 1501 40885 1535 40919
rect 17509 40885 17543 40919
rect 23121 40885 23155 40919
rect 23765 40885 23799 40919
rect 24409 40885 24443 40919
rect 24501 40885 24535 40919
rect 26341 40885 26375 40919
rect 31217 40885 31251 40919
rect 33149 40885 33183 40919
rect 34253 40885 34287 40919
rect 35817 40885 35851 40919
rect 36277 40885 36311 40919
rect 40417 40885 40451 40919
rect 42441 40885 42475 40919
rect 16037 40681 16071 40715
rect 17141 40681 17175 40715
rect 17969 40681 18003 40715
rect 20545 40681 20579 40715
rect 26985 40681 27019 40715
rect 30113 40681 30147 40715
rect 33701 40681 33735 40715
rect 35449 40681 35483 40715
rect 41061 40681 41095 40715
rect 16681 40613 16715 40647
rect 31401 40613 31435 40647
rect 34805 40613 34839 40647
rect 15577 40545 15611 40579
rect 20085 40545 20119 40579
rect 24501 40545 24535 40579
rect 26617 40545 26651 40579
rect 28917 40545 28951 40579
rect 29837 40545 29871 40579
rect 33241 40545 33275 40579
rect 33333 40545 33367 40579
rect 36277 40545 36311 40579
rect 17969 40477 18003 40511
rect 18429 40477 18463 40511
rect 18613 40477 18647 40511
rect 20729 40477 20763 40511
rect 20913 40477 20947 40511
rect 22845 40477 22879 40511
rect 23029 40477 23063 40511
rect 23489 40477 23523 40511
rect 23673 40477 23707 40511
rect 24593 40477 24627 40511
rect 26249 40477 26283 40511
rect 26433 40477 26467 40511
rect 26525 40477 26559 40511
rect 26801 40477 26835 40511
rect 27721 40477 27755 40511
rect 28457 40477 28491 40511
rect 29745 40477 29779 40511
rect 30757 40477 30791 40511
rect 30849 40477 30883 40511
rect 31585 40477 31619 40511
rect 31677 40477 31711 40511
rect 32229 40477 32263 40511
rect 32413 40477 32447 40511
rect 33425 40477 33459 40511
rect 33517 40477 33551 40511
rect 34713 40477 34747 40511
rect 34897 40477 34931 40511
rect 35357 40477 35391 40511
rect 35541 40477 35575 40511
rect 36645 40477 36679 40511
rect 36921 40477 36955 40511
rect 37289 40477 37323 40511
rect 39221 40477 39255 40511
rect 39865 40477 39899 40511
rect 40049 40477 40083 40511
rect 17693 40409 17727 40443
rect 17877 40409 17911 40443
rect 19533 40409 19567 40443
rect 36185 40409 36219 40443
rect 38485 40409 38519 40443
rect 41613 40409 41647 40443
rect 18521 40341 18555 40375
rect 21833 40341 21867 40375
rect 22385 40341 22419 40375
rect 22937 40341 22971 40375
rect 23857 40341 23891 40375
rect 24961 40341 24995 40375
rect 25789 40341 25823 40375
rect 30573 40341 30607 40375
rect 32321 40341 32355 40375
rect 39957 40341 39991 40375
rect 40509 40341 40543 40375
rect 17249 40137 17283 40171
rect 18337 40137 18371 40171
rect 23121 40137 23155 40171
rect 28089 40137 28123 40171
rect 30481 40137 30515 40171
rect 32229 40137 32263 40171
rect 34253 40137 34287 40171
rect 39405 40137 39439 40171
rect 40509 40137 40543 40171
rect 41061 40137 41095 40171
rect 17049 40069 17083 40103
rect 19165 40069 19199 40103
rect 34437 40069 34471 40103
rect 16129 40001 16163 40035
rect 18981 40001 19015 40035
rect 19625 40001 19659 40035
rect 19809 40001 19843 40035
rect 20729 40001 20763 40035
rect 22201 40001 22235 40035
rect 22385 40001 22419 40035
rect 23213 40001 23247 40035
rect 23305 40001 23339 40035
rect 23949 40001 23983 40035
rect 24225 40001 24259 40035
rect 24869 40001 24903 40035
rect 25053 40001 25087 40035
rect 25513 40001 25547 40035
rect 26433 40001 26467 40035
rect 27353 40001 27387 40035
rect 27905 40001 27939 40035
rect 29009 40001 29043 40035
rect 30113 40001 30147 40035
rect 30941 40001 30975 40035
rect 31125 40001 31159 40035
rect 33057 40001 33091 40035
rect 33149 40001 33183 40035
rect 33333 40001 33367 40035
rect 34621 40001 34655 40035
rect 35541 40001 35575 40035
rect 35725 40001 35759 40035
rect 36185 40001 36219 40035
rect 36369 40001 36403 40035
rect 37473 40001 37507 40035
rect 37657 40001 37691 40035
rect 38117 40001 38151 40035
rect 38301 40001 38335 40035
rect 38577 40001 38611 40035
rect 38945 40001 38979 40035
rect 39681 40001 39715 40035
rect 39773 40001 39807 40035
rect 39865 40001 39899 40035
rect 40049 40001 40083 40035
rect 52929 40001 52963 40035
rect 53573 40001 53607 40035
rect 17877 39933 17911 39967
rect 19717 39933 19751 39967
rect 22845 39933 22879 39967
rect 24133 39933 24167 39967
rect 25789 39933 25823 39967
rect 27077 39933 27111 39967
rect 27261 39933 27295 39967
rect 30021 39933 30055 39967
rect 31033 39933 31067 39967
rect 36277 39933 36311 39967
rect 53389 39933 53423 39967
rect 17417 39865 17451 39899
rect 18153 39865 18187 39899
rect 22293 39865 22327 39899
rect 25605 39865 25639 39899
rect 38301 39865 38335 39899
rect 41613 39865 41647 39899
rect 17233 39797 17267 39831
rect 18797 39797 18831 39831
rect 21189 39797 21223 39831
rect 23765 39797 23799 39831
rect 24685 39797 24719 39831
rect 24869 39797 24903 39831
rect 25513 39797 25547 39831
rect 27169 39797 27203 39831
rect 33333 39797 33367 39831
rect 35725 39797 35759 39831
rect 37565 39797 37599 39831
rect 21373 39593 21407 39627
rect 22385 39593 22419 39627
rect 31585 39593 31619 39627
rect 32689 39593 32723 39627
rect 33333 39593 33367 39627
rect 41521 39593 41555 39627
rect 18613 39525 18647 39559
rect 19993 39525 20027 39559
rect 23581 39525 23615 39559
rect 26525 39525 26559 39559
rect 34989 39525 35023 39559
rect 39865 39525 39899 39559
rect 17693 39457 17727 39491
rect 18153 39457 18187 39491
rect 23489 39457 23523 39491
rect 23857 39457 23891 39491
rect 26985 39457 27019 39491
rect 29745 39457 29779 39491
rect 30297 39457 30331 39491
rect 35541 39457 35575 39491
rect 36553 39457 36587 39491
rect 38393 39457 38427 39491
rect 15945 39389 15979 39423
rect 16129 39389 16163 39423
rect 16773 39389 16807 39423
rect 16957 39389 16991 39423
rect 17049 39389 17083 39423
rect 17785 39389 17819 39423
rect 19717 39389 19751 39423
rect 20453 39389 20487 39423
rect 20637 39389 20671 39423
rect 23213 39389 23247 39423
rect 23397 39389 23431 39423
rect 23673 39389 23707 39423
rect 24409 39389 24443 39423
rect 24593 39389 24627 39423
rect 24685 39389 24719 39423
rect 24777 39389 24811 39423
rect 24961 39389 24995 39423
rect 26249 39389 26283 39423
rect 27261 39389 27295 39423
rect 29837 39389 29871 39423
rect 30757 39389 30791 39423
rect 34713 39389 34747 39423
rect 35449 39389 35483 39423
rect 35633 39389 35667 39423
rect 36369 39389 36403 39423
rect 37473 39389 37507 39423
rect 37749 39389 37783 39423
rect 38485 39389 38519 39423
rect 14933 39321 14967 39355
rect 16589 39321 16623 39355
rect 19993 39321 20027 39355
rect 22569 39321 22603 39355
rect 22753 39321 22787 39355
rect 25789 39321 25823 39355
rect 26525 39321 26559 39355
rect 30435 39321 30469 39355
rect 30573 39321 30607 39355
rect 30665 39321 30699 39355
rect 31553 39321 31587 39355
rect 31769 39321 31803 39355
rect 33301 39321 33335 39355
rect 33517 39321 33551 39355
rect 34989 39321 35023 39355
rect 37657 39321 37691 39355
rect 40969 39321 41003 39355
rect 15485 39253 15519 39287
rect 16037 39253 16071 39287
rect 17509 39253 17543 39287
rect 19809 39253 19843 39287
rect 20545 39253 20579 39287
rect 21925 39253 21959 39287
rect 25145 39253 25179 39287
rect 26341 39253 26375 39287
rect 28365 39253 28399 39287
rect 30941 39253 30975 39287
rect 31401 39253 31435 39287
rect 33149 39253 33183 39287
rect 33977 39253 34011 39287
rect 34805 39253 34839 39287
rect 36185 39253 36219 39287
rect 37289 39253 37323 39287
rect 39313 39253 39347 39287
rect 40417 39253 40451 39287
rect 17601 39049 17635 39083
rect 17969 39049 18003 39083
rect 20177 39049 20211 39083
rect 20637 39049 20671 39083
rect 22385 39049 22419 39083
rect 23213 39049 23247 39083
rect 23857 39049 23891 39083
rect 24777 39049 24811 39083
rect 25329 39049 25363 39083
rect 26985 39049 27019 39083
rect 29009 39049 29043 39083
rect 29561 39049 29595 39083
rect 29929 39049 29963 39083
rect 35081 39049 35115 39083
rect 37447 39049 37481 39083
rect 38485 39049 38519 39083
rect 39497 39049 39531 39083
rect 40049 39049 40083 39083
rect 16037 38981 16071 39015
rect 16865 38981 16899 39015
rect 17049 38981 17083 39015
rect 18705 38981 18739 39015
rect 19809 38981 19843 39015
rect 20009 38981 20043 39015
rect 31585 38981 31619 39015
rect 35173 38981 35207 39015
rect 36461 38981 36495 39015
rect 37657 38981 37691 39015
rect 1869 38913 1903 38947
rect 15945 38913 15979 38947
rect 16129 38913 16163 38947
rect 17509 38913 17543 38947
rect 17785 38913 17819 38947
rect 18429 38913 18463 38947
rect 18521 38913 18555 38947
rect 21097 38913 21131 38947
rect 22017 38913 22051 38947
rect 23121 38913 23155 38947
rect 23305 38913 23339 38947
rect 23765 38913 23799 38947
rect 24041 38913 24075 38947
rect 27169 38913 27203 38947
rect 27353 38913 27387 38947
rect 27445 38913 27479 38947
rect 29469 38913 29503 38947
rect 29745 38913 29779 38947
rect 30665 38913 30699 38947
rect 30757 38913 30791 38947
rect 30941 38913 30975 38947
rect 31033 38913 31067 38947
rect 32404 38913 32438 38947
rect 34253 38913 34287 38947
rect 34437 38913 34471 38947
rect 35265 38913 35299 38947
rect 35449 38913 35483 38947
rect 36645 38913 36679 38947
rect 36737 38913 36771 38947
rect 38853 38913 38887 38947
rect 19349 38845 19383 38879
rect 21005 38845 21039 38879
rect 21281 38845 21315 38879
rect 21925 38845 21959 38879
rect 32137 38845 32171 38879
rect 34897 38845 34931 38879
rect 38945 38845 38979 38879
rect 18613 38777 18647 38811
rect 27905 38777 27939 38811
rect 1961 38709 1995 38743
rect 16681 38709 16715 38743
rect 19993 38709 20027 38743
rect 24225 38709 24259 38743
rect 25789 38709 25823 38743
rect 26341 38709 26375 38743
rect 30481 38709 30515 38743
rect 33517 38709 33551 38743
rect 34069 38709 34103 38743
rect 34437 38709 34471 38743
rect 36001 38709 36035 38743
rect 36461 38709 36495 38743
rect 37289 38709 37323 38743
rect 37473 38709 37507 38743
rect 40601 38709 40635 38743
rect 1593 38505 1627 38539
rect 16681 38505 16715 38539
rect 29009 38505 29043 38539
rect 30665 38505 30699 38539
rect 32965 38505 32999 38539
rect 34805 38505 34839 38539
rect 34989 38505 35023 38539
rect 36231 38505 36265 38539
rect 37013 38505 37047 38539
rect 23857 38437 23891 38471
rect 26709 38437 26743 38471
rect 27445 38437 27479 38471
rect 23029 38369 23063 38403
rect 27997 38369 28031 38403
rect 29929 38369 29963 38403
rect 31033 38369 31067 38403
rect 36369 38369 36403 38403
rect 15301 38301 15335 38335
rect 17233 38301 17267 38335
rect 17509 38301 17543 38335
rect 18153 38301 18187 38335
rect 18337 38301 18371 38335
rect 19257 38301 19291 38335
rect 19441 38301 19475 38335
rect 20177 38301 20211 38335
rect 20453 38301 20487 38335
rect 20913 38301 20947 38335
rect 21189 38301 21223 38335
rect 21833 38301 21867 38335
rect 22201 38301 22235 38335
rect 22845 38301 22879 38335
rect 24409 38301 24443 38335
rect 25237 38301 25271 38335
rect 25421 38301 25455 38335
rect 26065 38301 26099 38335
rect 26249 38301 26283 38335
rect 26709 38301 26743 38335
rect 26985 38301 27019 38335
rect 28733 38301 28767 38335
rect 28825 38301 28859 38335
rect 29837 38301 29871 38335
rect 31309 38301 31343 38335
rect 31953 38301 31987 38335
rect 32045 38301 32079 38335
rect 33241 38301 33275 38335
rect 33609 38301 33643 38335
rect 33701 38301 33735 38335
rect 36093 38301 36127 38335
rect 36553 38301 36587 38335
rect 37289 38301 37323 38335
rect 37473 38301 37507 38335
rect 38485 38301 38519 38335
rect 16313 38233 16347 38267
rect 16497 38233 16531 38267
rect 17325 38233 17359 38267
rect 19349 38233 19383 38267
rect 19993 38233 20027 38267
rect 21925 38233 21959 38267
rect 22661 38233 22695 38267
rect 24593 38233 24627 38267
rect 29009 38233 29043 38267
rect 30824 38233 30858 38267
rect 33333 38233 33367 38267
rect 35173 38233 35207 38267
rect 37933 38233 37967 38267
rect 39037 38233 39071 38267
rect 15853 38165 15887 38199
rect 17693 38165 17727 38199
rect 18153 38165 18187 38199
rect 20361 38165 20395 38199
rect 21005 38165 21039 38199
rect 21373 38165 21407 38199
rect 22017 38165 22051 38199
rect 22109 38165 22143 38199
rect 24777 38165 24811 38199
rect 25237 38165 25271 38199
rect 26157 38165 26191 38199
rect 26893 38165 26927 38199
rect 30205 38165 30239 38199
rect 30941 38165 30975 38199
rect 31769 38165 31803 38199
rect 33425 38165 33459 38199
rect 34973 38165 35007 38199
rect 36553 38165 36587 38199
rect 37197 38165 37231 38199
rect 39865 38165 39899 38199
rect 15577 37961 15611 37995
rect 17509 37961 17543 37995
rect 21833 37961 21867 37995
rect 25237 37961 25271 37995
rect 25421 37961 25455 37995
rect 33333 37961 33367 37995
rect 34069 37961 34103 37995
rect 35449 37961 35483 37995
rect 36185 37961 36219 37995
rect 16957 37893 16991 37927
rect 18429 37893 18463 37927
rect 18629 37893 18663 37927
rect 30113 37893 30147 37927
rect 17417 37825 17451 37859
rect 17693 37825 17727 37859
rect 19993 37825 20027 37859
rect 20177 37825 20211 37859
rect 21097 37825 21131 37859
rect 22017 37825 22051 37859
rect 22109 37825 22143 37859
rect 23397 37825 23431 37859
rect 23581 37825 23615 37859
rect 24501 37825 24535 37859
rect 25145 37825 25179 37859
rect 25513 37825 25547 37859
rect 25973 37825 26007 37859
rect 26433 37825 26467 37859
rect 26985 37825 27019 37859
rect 27241 37825 27275 37859
rect 30849 37825 30883 37859
rect 31401 37825 31435 37859
rect 32597 37825 32631 37859
rect 33057 37825 33091 37859
rect 33149 37825 33183 37859
rect 33977 37825 34011 37859
rect 34161 37825 34195 37859
rect 35541 37825 35575 37859
rect 36093 37825 36127 37859
rect 36277 37825 36311 37859
rect 37779 37825 37813 37859
rect 37933 37825 37967 37859
rect 20637 37757 20671 37791
rect 21005 37757 21039 37791
rect 21833 37757 21867 37791
rect 25329 37757 25363 37791
rect 26065 37757 26099 37791
rect 26295 37757 26329 37791
rect 29009 37757 29043 37791
rect 33333 37757 33367 37791
rect 18797 37689 18831 37723
rect 19993 37689 20027 37723
rect 23581 37689 23615 37723
rect 37565 37689 37599 37723
rect 16037 37621 16071 37655
rect 17877 37621 17911 37655
rect 18613 37621 18647 37655
rect 19717 37621 19751 37655
rect 21281 37621 21315 37655
rect 22937 37621 22971 37655
rect 24041 37621 24075 37655
rect 24225 37621 24259 37655
rect 26157 37621 26191 37655
rect 28365 37621 28399 37655
rect 32137 37621 32171 37655
rect 32505 37621 32539 37655
rect 34621 37621 34655 37655
rect 38393 37621 38427 37655
rect 38945 37621 38979 37655
rect 16589 37417 16623 37451
rect 17509 37417 17543 37451
rect 17601 37417 17635 37451
rect 18705 37417 18739 37451
rect 23857 37417 23891 37451
rect 26893 37417 26927 37451
rect 30849 37417 30883 37451
rect 33517 37417 33551 37451
rect 36369 37417 36403 37451
rect 38209 37417 38243 37451
rect 39037 37417 39071 37451
rect 52837 37417 52871 37451
rect 17417 37349 17451 37383
rect 19257 37349 19291 37383
rect 20269 37349 20303 37383
rect 22385 37349 22419 37383
rect 27077 37349 27111 37383
rect 29837 37349 29871 37383
rect 34161 37349 34195 37383
rect 35357 37349 35391 37383
rect 37289 37349 37323 37383
rect 37381 37349 37415 37383
rect 16037 37281 16071 37315
rect 17877 37281 17911 37315
rect 21833 37281 21867 37315
rect 23765 37281 23799 37315
rect 37013 37281 37047 37315
rect 17141 37213 17175 37247
rect 18429 37213 18463 37247
rect 18705 37213 18739 37247
rect 19625 37213 19659 37247
rect 20085 37213 20119 37247
rect 20269 37213 20303 37247
rect 20821 37213 20855 37247
rect 21005 37213 21039 37247
rect 22845 37213 22879 37247
rect 23029 37213 23063 37247
rect 23857 37213 23891 37247
rect 24685 37213 24719 37247
rect 24777 37213 24811 37247
rect 24869 37213 24903 37247
rect 25053 37213 25087 37247
rect 25789 37213 25823 37247
rect 28365 37213 28399 37247
rect 28549 37213 28583 37247
rect 29745 37213 29779 37247
rect 29929 37213 29963 37247
rect 30021 37213 30055 37247
rect 30205 37213 30239 37247
rect 31033 37213 31067 37247
rect 31309 37213 31343 37247
rect 31769 37213 31803 37247
rect 32873 37213 32907 37247
rect 33977 37213 34011 37247
rect 34161 37213 34195 37247
rect 34713 37213 34747 37247
rect 34897 37213 34931 37247
rect 36369 37213 36403 37247
rect 36553 37213 36587 37247
rect 37197 37213 37231 37247
rect 37473 37213 37507 37247
rect 37657 37213 37691 37247
rect 38117 37213 38151 37247
rect 53389 37213 53423 37247
rect 19441 37145 19475 37179
rect 22937 37145 22971 37179
rect 25513 37145 25547 37179
rect 25697 37145 25731 37179
rect 26709 37145 26743 37179
rect 26909 37145 26943 37179
rect 31217 37145 31251 37179
rect 17233 37077 17267 37111
rect 18521 37077 18555 37111
rect 21005 37077 21039 37111
rect 23489 37077 23523 37111
rect 24409 37077 24443 37111
rect 25611 37077 25645 37111
rect 27629 37077 27663 37111
rect 28457 37077 28491 37111
rect 29561 37077 29595 37111
rect 32413 37077 32447 37111
rect 34805 37077 34839 37111
rect 38577 37077 38611 37111
rect 53573 37077 53607 37111
rect 18245 36873 18279 36907
rect 19717 36873 19751 36907
rect 21005 36873 21039 36907
rect 22017 36873 22051 36907
rect 23765 36873 23799 36907
rect 28089 36873 28123 36907
rect 30941 36873 30975 36907
rect 33701 36873 33735 36907
rect 37657 36873 37691 36907
rect 17509 36805 17543 36839
rect 20269 36805 20303 36839
rect 30389 36805 30423 36839
rect 34989 36805 35023 36839
rect 17417 36737 17451 36771
rect 17693 36737 17727 36771
rect 18153 36737 18187 36771
rect 18429 36737 18463 36771
rect 21005 36737 21039 36771
rect 23029 36737 23063 36771
rect 23213 36737 23247 36771
rect 23673 36737 23707 36771
rect 23857 36737 23891 36771
rect 24501 36737 24535 36771
rect 24593 36737 24627 36771
rect 25697 36737 25731 36771
rect 26985 36737 27019 36771
rect 27077 36737 27111 36771
rect 30849 36737 30883 36771
rect 31033 36737 31067 36771
rect 32137 36737 32171 36771
rect 33425 36737 33459 36771
rect 33517 36737 33551 36771
rect 34345 36737 34379 36771
rect 35173 36737 35207 36771
rect 36553 36737 36587 36771
rect 38301 36737 38335 36771
rect 38669 36737 38703 36771
rect 39313 36737 39347 36771
rect 39405 36737 39439 36771
rect 39497 36737 39531 36771
rect 20729 36669 20763 36703
rect 22569 36669 22603 36703
rect 24409 36669 24443 36703
rect 24685 36669 24719 36703
rect 25421 36669 25455 36703
rect 27261 36669 27295 36703
rect 32781 36669 32815 36703
rect 34161 36669 34195 36703
rect 36645 36669 36679 36703
rect 17601 36601 17635 36635
rect 20913 36601 20947 36635
rect 23121 36601 23155 36635
rect 25513 36601 25547 36635
rect 29101 36601 29135 36635
rect 36185 36601 36219 36635
rect 39681 36601 39715 36635
rect 18613 36533 18647 36567
rect 19165 36533 19199 36567
rect 24869 36533 24903 36567
rect 25881 36533 25915 36567
rect 26341 36533 26375 36567
rect 27169 36533 27203 36567
rect 31493 36533 31527 36567
rect 34529 36533 34563 36567
rect 35357 36533 35391 36567
rect 20637 36329 20671 36363
rect 23489 36329 23523 36363
rect 24777 36329 24811 36363
rect 30573 36329 30607 36363
rect 35541 36329 35575 36363
rect 38761 36329 38795 36363
rect 17877 36261 17911 36295
rect 17969 36261 18003 36295
rect 29653 36261 29687 36295
rect 34989 36261 35023 36295
rect 20545 36193 20579 36227
rect 21649 36193 21683 36227
rect 22201 36193 22235 36227
rect 26617 36193 26651 36227
rect 26893 36193 26927 36227
rect 28733 36193 28767 36227
rect 31033 36193 31067 36227
rect 32689 36193 32723 36227
rect 32965 36193 32999 36227
rect 33885 36193 33919 36227
rect 35725 36193 35759 36227
rect 36645 36193 36679 36227
rect 37105 36193 37139 36227
rect 37657 36193 37691 36227
rect 37841 36193 37875 36227
rect 38301 36193 38335 36227
rect 17785 36125 17819 36159
rect 18061 36125 18095 36159
rect 18245 36125 18279 36159
rect 19441 36125 19475 36159
rect 19533 36125 19567 36159
rect 20453 36125 20487 36159
rect 21465 36125 21499 36159
rect 22109 36125 22143 36159
rect 22293 36125 22327 36159
rect 24593 36125 24627 36159
rect 24777 36125 24811 36159
rect 29009 36125 29043 36159
rect 29653 36125 29687 36159
rect 30757 36125 30791 36159
rect 30849 36125 30883 36159
rect 31125 36125 31159 36159
rect 32597 36125 32631 36159
rect 33609 36125 33643 36159
rect 33793 36125 33827 36159
rect 33977 36123 34011 36157
rect 34161 36127 34195 36161
rect 34713 36125 34747 36159
rect 35449 36125 35483 36159
rect 37013 36125 37047 36159
rect 37933 36125 37967 36159
rect 38761 36125 38795 36159
rect 38945 36125 38979 36159
rect 1869 36057 1903 36091
rect 17141 36057 17175 36091
rect 19257 36057 19291 36091
rect 23673 36057 23707 36091
rect 23857 36057 23891 36091
rect 25237 36057 25271 36091
rect 34989 36057 35023 36091
rect 1961 35989 1995 36023
rect 16589 35989 16623 36023
rect 17601 35989 17635 36023
rect 19533 35989 19567 36023
rect 20821 35989 20855 36023
rect 21281 35989 21315 36023
rect 23029 35989 23063 36023
rect 27445 35989 27479 36023
rect 31585 35989 31619 36023
rect 33425 35989 33459 36023
rect 34805 35989 34839 36023
rect 35725 35989 35759 36023
rect 39865 35989 39899 36023
rect 40509 35989 40543 36023
rect 1685 35785 1719 35819
rect 18061 35785 18095 35819
rect 19257 35785 19291 35819
rect 20009 35785 20043 35819
rect 20177 35785 20211 35819
rect 25237 35785 25271 35819
rect 26341 35785 26375 35819
rect 34345 35785 34379 35819
rect 34805 35785 34839 35819
rect 36553 35785 36587 35819
rect 37289 35785 37323 35819
rect 38853 35785 38887 35819
rect 39497 35785 39531 35819
rect 17509 35717 17543 35751
rect 19809 35717 19843 35751
rect 25789 35717 25823 35751
rect 30389 35717 30423 35751
rect 36737 35717 36771 35751
rect 37457 35717 37491 35751
rect 37657 35717 37691 35751
rect 40509 35717 40543 35751
rect 17417 35649 17451 35683
rect 17601 35649 17635 35683
rect 18521 35649 18555 35683
rect 19073 35649 19107 35683
rect 19349 35649 19383 35683
rect 20637 35649 20671 35683
rect 20821 35649 20855 35683
rect 21097 35649 21131 35683
rect 22017 35649 22051 35683
rect 24133 35649 24167 35683
rect 24317 35649 24351 35683
rect 24409 35649 24443 35683
rect 26065 35649 26099 35683
rect 27169 35649 27203 35683
rect 32137 35649 32171 35683
rect 32316 35649 32350 35683
rect 32413 35649 32447 35683
rect 32505 35649 32539 35683
rect 33885 35649 33919 35683
rect 34161 35649 34195 35683
rect 34979 35649 35013 35683
rect 35081 35649 35115 35683
rect 35265 35649 35299 35683
rect 36461 35649 36495 35683
rect 38117 35649 38151 35683
rect 38301 35649 38335 35683
rect 38761 35649 38795 35683
rect 38945 35649 38979 35683
rect 20913 35581 20947 35615
rect 21925 35581 21959 35615
rect 22385 35581 22419 35615
rect 25697 35581 25731 35615
rect 26188 35581 26222 35615
rect 26985 35581 27019 35615
rect 31401 35581 31435 35615
rect 34069 35581 34103 35615
rect 35173 35581 35207 35615
rect 38209 35581 38243 35615
rect 19073 35513 19107 35547
rect 21005 35513 21039 35547
rect 22937 35513 22971 35547
rect 24225 35513 24259 35547
rect 27353 35513 27387 35547
rect 29101 35513 29135 35547
rect 33977 35513 34011 35547
rect 36737 35513 36771 35547
rect 16037 35445 16071 35479
rect 16865 35445 16899 35479
rect 18245 35445 18279 35479
rect 19993 35445 20027 35479
rect 21281 35445 21315 35479
rect 23397 35445 23431 35479
rect 23949 35445 23983 35479
rect 28089 35445 28123 35479
rect 30941 35445 30975 35479
rect 32781 35445 32815 35479
rect 33241 35445 33275 35479
rect 35817 35445 35851 35479
rect 37473 35445 37507 35479
rect 40049 35445 40083 35479
rect 16957 35241 16991 35275
rect 20821 35241 20855 35275
rect 21005 35241 21039 35275
rect 21741 35241 21775 35275
rect 23765 35241 23799 35275
rect 24501 35241 24535 35275
rect 24777 35241 24811 35275
rect 26157 35241 26191 35275
rect 28825 35241 28859 35275
rect 37473 35241 37507 35275
rect 38393 35241 38427 35275
rect 39865 35241 39899 35275
rect 22937 35173 22971 35207
rect 29653 35173 29687 35207
rect 33793 35173 33827 35207
rect 36185 35173 36219 35207
rect 36737 35173 36771 35207
rect 17509 35105 17543 35139
rect 17969 35105 18003 35139
rect 21097 35105 21131 35139
rect 21833 35105 21867 35139
rect 22753 35105 22787 35139
rect 26617 35105 26651 35139
rect 15853 35037 15887 35071
rect 16865 35037 16899 35071
rect 17049 35037 17083 35071
rect 17693 35037 17727 35071
rect 18061 35037 18095 35071
rect 18521 35037 18555 35071
rect 18705 35037 18739 35071
rect 19441 35037 19475 35071
rect 19809 35037 19843 35071
rect 19901 35037 19935 35071
rect 21005 35037 21039 35071
rect 21741 35037 21775 35071
rect 22569 35037 22603 35071
rect 22937 35037 22971 35071
rect 24777 35037 24811 35071
rect 24961 35037 24995 35071
rect 26893 35037 26927 35071
rect 28273 35037 28307 35071
rect 29929 35037 29963 35071
rect 31697 35037 31731 35071
rect 31953 35037 31987 35071
rect 32413 35037 32447 35071
rect 32680 35037 32714 35071
rect 34713 35037 34747 35071
rect 35449 35037 35483 35071
rect 35633 35037 35667 35071
rect 37841 35037 37875 35071
rect 18613 34969 18647 35003
rect 19579 34969 19613 35003
rect 19717 34969 19751 35003
rect 21281 34969 21315 35003
rect 29653 34969 29687 35003
rect 37657 34969 37691 35003
rect 52929 34969 52963 35003
rect 53573 34969 53607 35003
rect 16313 34901 16347 34935
rect 20085 34901 20119 34935
rect 22109 34901 22143 34935
rect 22661 34901 22695 34935
rect 25605 34901 25639 34935
rect 29837 34901 29871 34935
rect 30573 34901 30607 34935
rect 34897 34901 34931 34935
rect 35449 34901 35483 34935
rect 38853 34901 38887 34935
rect 53481 34901 53515 34935
rect 15485 34697 15519 34731
rect 16129 34697 16163 34731
rect 17601 34697 17635 34731
rect 18889 34697 18923 34731
rect 21281 34697 21315 34731
rect 25145 34697 25179 34731
rect 26433 34697 26467 34731
rect 30757 34697 30791 34731
rect 31486 34697 31520 34731
rect 34161 34697 34195 34731
rect 36553 34697 36587 34731
rect 37565 34697 37599 34731
rect 38669 34697 38703 34731
rect 39221 34697 39255 34731
rect 16773 34629 16807 34663
rect 17233 34629 17267 34663
rect 17449 34629 17483 34663
rect 19073 34629 19107 34663
rect 22385 34629 22419 34663
rect 23581 34629 23615 34663
rect 25424 34629 25458 34663
rect 28641 34629 28675 34663
rect 31401 34629 31435 34663
rect 31585 34629 31619 34663
rect 32137 34629 32171 34663
rect 33393 34629 33427 34663
rect 33609 34629 33643 34663
rect 35265 34629 35299 34663
rect 1869 34561 1903 34595
rect 18245 34561 18279 34595
rect 19257 34561 19291 34595
rect 19901 34561 19935 34595
rect 21005 34561 21039 34595
rect 21097 34561 21131 34595
rect 22201 34561 22235 34595
rect 25283 34561 25317 34595
rect 25513 34561 25547 34595
rect 25641 34561 25675 34595
rect 25789 34561 25823 34595
rect 26985 34561 27019 34595
rect 27169 34561 27203 34595
rect 28825 34561 28859 34595
rect 29101 34561 29135 34595
rect 29837 34561 29871 34595
rect 30665 34561 30699 34595
rect 30849 34561 30883 34595
rect 31309 34561 31343 34595
rect 32413 34561 32447 34595
rect 32505 34561 32539 34595
rect 32597 34561 32631 34595
rect 32781 34561 32815 34595
rect 34529 34561 34563 34595
rect 35173 34561 35207 34595
rect 35357 34561 35391 34595
rect 35817 34561 35851 34595
rect 36001 34561 36035 34595
rect 37381 34561 37415 34595
rect 37565 34561 37599 34595
rect 2053 34493 2087 34527
rect 18429 34493 18463 34527
rect 19809 34493 19843 34527
rect 21281 34493 21315 34527
rect 29009 34493 29043 34527
rect 29929 34493 29963 34527
rect 30205 34493 30239 34527
rect 34621 34493 34655 34527
rect 20269 34425 20303 34459
rect 24133 34425 24167 34459
rect 28917 34425 28951 34459
rect 17417 34357 17451 34391
rect 18061 34357 18095 34391
rect 22569 34357 22603 34391
rect 24685 34357 24719 34391
rect 27169 34357 27203 34391
rect 28181 34357 28215 34391
rect 33241 34357 33275 34391
rect 33425 34357 33459 34391
rect 35909 34357 35943 34391
rect 38025 34357 38059 34391
rect 17417 34153 17451 34187
rect 17969 34153 18003 34187
rect 19901 34153 19935 34187
rect 19993 34153 20027 34187
rect 25513 34153 25547 34187
rect 26065 34153 26099 34187
rect 26249 34153 26283 34187
rect 26893 34153 26927 34187
rect 27813 34153 27847 34187
rect 32505 34153 32539 34187
rect 32689 34153 32723 34187
rect 35909 34153 35943 34187
rect 36553 34153 36587 34187
rect 1593 34085 1627 34119
rect 19349 34085 19383 34119
rect 23857 34085 23891 34119
rect 28917 34085 28951 34119
rect 34069 34085 34103 34119
rect 34989 34085 35023 34119
rect 16405 34017 16439 34051
rect 20085 34017 20119 34051
rect 22109 34017 22143 34051
rect 23581 34017 23615 34051
rect 25329 34017 25363 34051
rect 27905 34017 27939 34051
rect 28457 34017 28491 34051
rect 29837 34017 29871 34051
rect 31217 34017 31251 34051
rect 35081 34017 35115 34051
rect 18153 33949 18187 33983
rect 19809 33949 19843 33983
rect 20913 33949 20947 33983
rect 22017 33949 22051 33983
rect 22201 33949 22235 33983
rect 22661 33949 22695 33983
rect 22845 33949 22879 33983
rect 23489 33949 23523 33983
rect 25237 33949 25271 33983
rect 26893 33949 26927 33983
rect 27169 33949 27203 33983
rect 27629 33949 27663 33983
rect 27721 33949 27755 33983
rect 28549 33949 28583 33983
rect 29745 33949 29779 33983
rect 30849 33949 30883 33983
rect 31309 33949 31343 33983
rect 32781 33949 32815 33983
rect 32873 33949 32907 33983
rect 33885 33949 33919 33983
rect 34161 33949 34195 33983
rect 34897 33949 34931 33983
rect 35173 33949 35207 33983
rect 38853 33949 38887 33983
rect 18337 33881 18371 33915
rect 22753 33881 22787 33915
rect 26433 33881 26467 33915
rect 34713 33881 34747 33915
rect 35893 33881 35927 33915
rect 36093 33881 36127 33915
rect 37105 33881 37139 33915
rect 16865 33813 16899 33847
rect 21465 33813 21499 33847
rect 24501 33813 24535 33847
rect 26228 33813 26262 33847
rect 27077 33813 27111 33847
rect 30113 33813 30147 33847
rect 33701 33813 33735 33847
rect 35725 33813 35759 33847
rect 37657 33813 37691 33847
rect 38209 33813 38243 33847
rect 39957 33813 39991 33847
rect 18061 33609 18095 33643
rect 18981 33609 19015 33643
rect 24685 33609 24719 33643
rect 26433 33609 26467 33643
rect 29377 33609 29411 33643
rect 31309 33609 31343 33643
rect 32866 33609 32900 33643
rect 33517 33609 33551 33643
rect 35081 33609 35115 33643
rect 35909 33609 35943 33643
rect 17509 33541 17543 33575
rect 24041 33541 24075 33575
rect 25237 33541 25271 33575
rect 30481 33541 30515 33575
rect 30697 33541 30731 33575
rect 16957 33473 16991 33507
rect 17969 33473 18003 33507
rect 18153 33473 18187 33507
rect 22477 33473 22511 33507
rect 22661 33473 22695 33507
rect 23305 33473 23339 33507
rect 27169 33473 27203 33507
rect 27261 33473 27295 33507
rect 27537 33473 27571 33507
rect 28089 33473 28123 33507
rect 28549 33473 28583 33507
rect 28733 33473 28767 33507
rect 29607 33473 29641 33507
rect 29742 33473 29776 33507
rect 29837 33473 29871 33507
rect 30021 33473 30055 33507
rect 31309 33473 31343 33507
rect 31493 33473 31527 33507
rect 32689 33473 32723 33507
rect 32781 33473 32815 33507
rect 32965 33473 32999 33507
rect 34437 33473 34471 33507
rect 35265 33473 35299 33507
rect 35449 33473 35483 33507
rect 36093 33473 36127 33507
rect 36277 33473 36311 33507
rect 37473 33473 37507 33507
rect 38945 33473 38979 33507
rect 39129 33473 39163 33507
rect 39773 33473 39807 33507
rect 40417 33473 40451 33507
rect 40969 33473 41003 33507
rect 20085 33405 20119 33439
rect 21833 33405 21867 33439
rect 23581 33405 23615 33439
rect 27445 33405 27479 33439
rect 28917 33405 28951 33439
rect 32229 33405 32263 33439
rect 34345 33405 34379 33439
rect 37381 33405 37415 33439
rect 37841 33405 37875 33439
rect 39957 33405 39991 33439
rect 20729 33337 20763 33371
rect 22569 33337 22603 33371
rect 34069 33337 34103 33371
rect 39589 33337 39623 33371
rect 19441 33269 19475 33303
rect 21189 33269 21223 33303
rect 23121 33269 23155 33303
rect 23489 33269 23523 33303
rect 25789 33269 25823 33303
rect 26985 33269 27019 33303
rect 30665 33269 30699 33303
rect 30849 33269 30883 33303
rect 39037 33269 39071 33303
rect 19257 33065 19291 33099
rect 33609 33065 33643 33099
rect 35357 33065 35391 33099
rect 37933 33065 37967 33099
rect 38945 33065 38979 33099
rect 26617 32997 26651 33031
rect 28917 32997 28951 33031
rect 38393 32997 38427 33031
rect 18337 32929 18371 32963
rect 20821 32929 20855 32963
rect 22937 32929 22971 32963
rect 24501 32929 24535 32963
rect 29653 32929 29687 32963
rect 39865 32929 39899 32963
rect 18061 32861 18095 32895
rect 18153 32861 18187 32895
rect 19257 32861 19291 32895
rect 19349 32861 19383 32895
rect 20085 32861 20119 32895
rect 20269 32861 20303 32895
rect 22109 32861 22143 32895
rect 23121 32861 23155 32895
rect 24593 32861 24627 32895
rect 25421 32861 25455 32895
rect 25605 32861 25639 32895
rect 25697 32861 25731 32895
rect 25789 32861 25823 32895
rect 27997 32861 28031 32895
rect 28825 32861 28859 32895
rect 29009 32861 29043 32895
rect 30297 32861 30331 32895
rect 31125 32861 31159 32895
rect 31309 32861 31343 32895
rect 32321 32861 32355 32895
rect 32413 32861 32447 32895
rect 33057 32861 33091 32895
rect 34161 32861 34195 32895
rect 35081 32861 35115 32895
rect 35357 32861 35391 32895
rect 35817 32861 35851 32895
rect 36645 32861 36679 32895
rect 36829 32861 36863 32895
rect 21925 32793 21959 32827
rect 26065 32793 26099 32827
rect 27730 32793 27764 32827
rect 30113 32793 30147 32827
rect 32137 32793 32171 32827
rect 36001 32793 36035 32827
rect 16865 32725 16899 32759
rect 18337 32725 18371 32759
rect 19625 32725 19659 32759
rect 20177 32725 20211 32759
rect 21373 32725 21407 32759
rect 22293 32725 22327 32759
rect 23305 32725 23339 32759
rect 23857 32725 23891 32759
rect 24961 32725 24995 32759
rect 30481 32725 30515 32759
rect 30941 32725 30975 32759
rect 35173 32725 35207 32759
rect 36185 32725 36219 32759
rect 36737 32725 36771 32759
rect 37381 32725 37415 32759
rect 40417 32725 40451 32759
rect 18153 32521 18187 32555
rect 19349 32521 19383 32555
rect 25605 32521 25639 32555
rect 28457 32521 28491 32555
rect 29009 32521 29043 32555
rect 29653 32521 29687 32555
rect 32873 32521 32907 32555
rect 33701 32521 33735 32555
rect 35817 32521 35851 32555
rect 37289 32521 37323 32555
rect 38209 32521 38243 32555
rect 38669 32521 38703 32555
rect 18981 32453 19015 32487
rect 19197 32453 19231 32487
rect 20085 32453 20119 32487
rect 26985 32453 27019 32487
rect 30593 32453 30627 32487
rect 1685 32385 1719 32419
rect 2237 32385 2271 32419
rect 17417 32385 17451 32419
rect 18337 32385 18371 32419
rect 18429 32385 18463 32419
rect 19809 32385 19843 32419
rect 19901 32385 19935 32419
rect 20821 32385 20855 32419
rect 21925 32385 21959 32419
rect 22109 32385 22143 32419
rect 22569 32385 22603 32419
rect 22753 32385 22787 32419
rect 23213 32385 23247 32419
rect 23581 32385 23615 32419
rect 24225 32385 24259 32419
rect 24409 32385 24443 32419
rect 24501 32385 24535 32419
rect 25513 32385 25547 32419
rect 25697 32385 25731 32419
rect 29561 32385 29595 32419
rect 29745 32385 29779 32419
rect 30205 32385 30239 32419
rect 30298 32385 30332 32419
rect 30481 32385 30515 32419
rect 30711 32385 30745 32419
rect 31309 32385 31343 32419
rect 32321 32385 32355 32419
rect 32413 32385 32447 32419
rect 32873 32385 32907 32419
rect 33149 32385 33183 32419
rect 35633 32385 35667 32419
rect 35817 32385 35851 32419
rect 36277 32385 36311 32419
rect 37473 32385 37507 32419
rect 52929 32385 52963 32419
rect 53573 32385 53607 32419
rect 16957 32317 16991 32351
rect 17693 32317 17727 32351
rect 20729 32317 20763 32351
rect 22017 32317 22051 32351
rect 31585 32317 31619 32351
rect 32137 32317 32171 32351
rect 37657 32317 37691 32351
rect 17601 32249 17635 32283
rect 20085 32249 20119 32283
rect 21189 32249 21223 32283
rect 30849 32249 30883 32283
rect 32965 32249 32999 32283
rect 53389 32249 53423 32283
rect 1501 32181 1535 32215
rect 17509 32181 17543 32215
rect 19165 32181 19199 32215
rect 22661 32181 22695 32215
rect 23305 32181 23339 32215
rect 23765 32181 23799 32215
rect 24225 32181 24259 32215
rect 24685 32181 24719 32215
rect 26157 32181 26191 32215
rect 31401 32181 31435 32215
rect 31493 32181 31527 32215
rect 32229 32181 32263 32215
rect 34253 32181 34287 32215
rect 34713 32181 34747 32215
rect 36369 32181 36403 32215
rect 15485 31977 15519 32011
rect 16037 31977 16071 32011
rect 18153 31977 18187 32011
rect 18521 31977 18555 32011
rect 23489 31977 23523 32011
rect 24501 31977 24535 32011
rect 26433 31977 26467 32011
rect 31677 31977 31711 32011
rect 19257 31909 19291 31943
rect 25605 31909 25639 31943
rect 29009 31909 29043 31943
rect 29745 31909 29779 31943
rect 33057 31909 33091 31943
rect 33701 31909 33735 31943
rect 34713 31909 34747 31943
rect 36093 31909 36127 31943
rect 36829 31909 36863 31943
rect 17601 31841 17635 31875
rect 21649 31841 21683 31875
rect 24685 31841 24719 31875
rect 30665 31841 30699 31875
rect 31217 31841 31251 31875
rect 32597 31841 32631 31875
rect 36645 31841 36679 31875
rect 37565 31841 37599 31875
rect 37933 31841 37967 31875
rect 16589 31773 16623 31807
rect 16773 31773 16807 31807
rect 17417 31773 17451 31807
rect 18061 31773 18095 31807
rect 19625 31773 19659 31807
rect 20453 31773 20487 31807
rect 20729 31773 20763 31807
rect 21465 31773 21499 31807
rect 22201 31773 22235 31807
rect 22293 31773 22327 31807
rect 23213 31773 23247 31807
rect 23489 31773 23523 31807
rect 24409 31773 24443 31807
rect 25789 31773 25823 31807
rect 25881 31773 25915 31807
rect 26985 31773 27019 31807
rect 30389 31773 30423 31807
rect 30481 31773 30515 31807
rect 30757 31773 30791 31807
rect 31401 31773 31435 31807
rect 31493 31773 31527 31807
rect 31769 31773 31803 31807
rect 32229 31773 32263 31807
rect 32413 31773 32447 31807
rect 33057 31773 33091 31807
rect 33241 31773 33275 31807
rect 33885 31773 33919 31807
rect 34161 31773 34195 31807
rect 35357 31773 35391 31807
rect 36553 31773 36587 31807
rect 37473 31773 37507 31807
rect 38485 31773 38519 31807
rect 19441 31705 19475 31739
rect 20637 31705 20671 31739
rect 21281 31705 21315 31739
rect 22477 31705 22511 31739
rect 25605 31705 25639 31739
rect 34069 31705 34103 31739
rect 36093 31705 36127 31739
rect 16681 31637 16715 31671
rect 17233 31637 17267 31671
rect 20269 31637 20303 31671
rect 23305 31637 23339 31671
rect 24961 31637 24995 31671
rect 30205 31637 30239 31671
rect 37289 31637 37323 31671
rect 16037 31433 16071 31467
rect 17693 31433 17727 31467
rect 22753 31433 22787 31467
rect 23673 31433 23707 31467
rect 25973 31433 26007 31467
rect 33793 31433 33827 31467
rect 35909 31433 35943 31467
rect 37657 31433 37691 31467
rect 22661 31365 22695 31399
rect 23581 31365 23615 31399
rect 31585 31365 31619 31399
rect 35265 31365 35299 31399
rect 16957 31297 16991 31331
rect 17141 31297 17175 31331
rect 17601 31297 17635 31331
rect 17785 31297 17819 31331
rect 18245 31297 18279 31331
rect 18408 31297 18442 31331
rect 18521 31297 18555 31331
rect 18659 31297 18693 31331
rect 19533 31297 19567 31331
rect 20545 31297 20579 31331
rect 21925 31297 21959 31331
rect 22109 31297 22143 31331
rect 22569 31297 22603 31331
rect 22845 31297 22879 31331
rect 23765 31297 23799 31331
rect 24501 31297 24535 31331
rect 25421 31297 25455 31331
rect 25697 31297 25731 31331
rect 25789 31297 25823 31331
rect 26985 31297 27019 31331
rect 27261 31297 27295 31331
rect 29377 31297 29411 31331
rect 29561 31297 29595 31331
rect 31309 31297 31343 31331
rect 32137 31297 32171 31331
rect 32229 31297 32263 31331
rect 32505 31297 32539 31331
rect 33149 31297 33183 31331
rect 34069 31297 34103 31331
rect 34161 31297 34195 31331
rect 34253 31297 34287 31331
rect 34437 31297 34471 31331
rect 35081 31297 35115 31331
rect 36277 31297 36311 31331
rect 37749 31297 37783 31331
rect 19625 31229 19659 31263
rect 19901 31229 19935 31263
rect 20453 31229 20487 31263
rect 23305 31229 23339 31263
rect 23397 31229 23431 31263
rect 30021 31229 30055 31263
rect 31585 31229 31619 31263
rect 32321 31229 32355 31263
rect 33333 31229 33367 31263
rect 36369 31229 36403 31263
rect 37289 31229 37323 31263
rect 20913 31161 20947 31195
rect 25513 31161 25547 31195
rect 30757 31161 30791 31195
rect 31401 31161 31435 31195
rect 35449 31161 35483 31195
rect 16957 31093 16991 31127
rect 18889 31093 18923 31127
rect 22017 31093 22051 31127
rect 24041 31093 24075 31127
rect 24593 31093 24627 31127
rect 28365 31093 28399 31127
rect 29561 31093 29595 31127
rect 32505 31093 32539 31127
rect 32965 31093 32999 31127
rect 37473 31093 37507 31127
rect 38209 31093 38243 31127
rect 21649 30889 21683 30923
rect 23397 30889 23431 30923
rect 25973 30889 26007 30923
rect 26065 30889 26099 30923
rect 27261 30889 27295 30923
rect 28273 30889 28307 30923
rect 31125 30889 31159 30923
rect 31953 30889 31987 30923
rect 32321 30889 32355 30923
rect 32781 30889 32815 30923
rect 34713 30889 34747 30923
rect 35633 30889 35667 30923
rect 18613 30821 18647 30855
rect 21005 30821 21039 30855
rect 22753 30821 22787 30855
rect 18337 30753 18371 30787
rect 20361 30753 20395 30787
rect 20821 30753 20855 30787
rect 24685 30753 24719 30787
rect 25881 30753 25915 30787
rect 29561 30753 29595 30787
rect 33793 30753 33827 30787
rect 36369 30753 36403 30787
rect 36461 30753 36495 30787
rect 36645 30753 36679 30787
rect 18245 30685 18279 30719
rect 19901 30685 19935 30719
rect 20177 30685 20211 30719
rect 21097 30685 21131 30719
rect 21557 30685 21591 30719
rect 21741 30685 21775 30719
rect 23213 30685 23247 30719
rect 23489 30685 23523 30719
rect 24777 30685 24811 30719
rect 26157 30685 26191 30719
rect 26709 30685 26743 30719
rect 29837 30685 29871 30719
rect 31953 30685 31987 30719
rect 32045 30685 32079 30719
rect 33701 30685 33735 30719
rect 35541 30685 35575 30719
rect 35725 30685 35759 30719
rect 36553 30685 36587 30719
rect 19441 30617 19475 30651
rect 19993 30617 20027 30651
rect 23305 30617 23339 30651
rect 37289 30617 37323 30651
rect 37749 30617 37783 30651
rect 16957 30549 16991 30583
rect 17509 30549 17543 30583
rect 20821 30549 20855 30583
rect 24409 30549 24443 30583
rect 27721 30549 27755 30583
rect 33333 30549 33367 30583
rect 36185 30549 36219 30583
rect 23029 30345 23063 30379
rect 23765 30345 23799 30379
rect 25697 30345 25731 30379
rect 31033 30345 31067 30379
rect 33517 30345 33551 30379
rect 34069 30345 34103 30379
rect 36277 30345 36311 30379
rect 37381 30345 37415 30379
rect 18705 30277 18739 30311
rect 19257 30277 19291 30311
rect 21925 30277 21959 30311
rect 24961 30277 24995 30311
rect 32404 30277 32438 30311
rect 20821 30209 20855 30243
rect 21005 30209 21039 30243
rect 21833 30209 21867 30243
rect 22017 30209 22051 30243
rect 22937 30209 22971 30243
rect 23121 30209 23155 30243
rect 23581 30209 23615 30243
rect 23765 30209 23799 30243
rect 24225 30209 24259 30243
rect 24409 30209 24443 30243
rect 24869 30209 24903 30243
rect 25237 30209 25271 30243
rect 25881 30209 25915 30243
rect 26985 30209 27019 30243
rect 28641 30209 28675 30243
rect 34989 30209 35023 30243
rect 35173 30209 35207 30243
rect 35265 30209 35299 30243
rect 36185 30209 36219 30243
rect 36369 30209 36403 30243
rect 52929 30209 52963 30243
rect 53573 30209 53607 30243
rect 24317 30141 24351 30175
rect 25053 30141 25087 30175
rect 26065 30141 26099 30175
rect 27261 30141 27295 30175
rect 32137 30141 32171 30175
rect 25237 30073 25271 30107
rect 17969 30005 18003 30039
rect 19809 30005 19843 30039
rect 20361 30005 20395 30039
rect 20913 30005 20947 30039
rect 35265 30005 35299 30039
rect 53481 30005 53515 30039
rect 18705 29801 18739 29835
rect 23581 29801 23615 29835
rect 25145 29801 25179 29835
rect 26157 29801 26191 29835
rect 30205 29801 30239 29835
rect 33057 29801 33091 29835
rect 34069 29801 34103 29835
rect 36461 29801 36495 29835
rect 20729 29733 20763 29767
rect 23029 29733 23063 29767
rect 24501 29733 24535 29767
rect 21189 29665 21223 29699
rect 22201 29665 22235 29699
rect 24685 29665 24719 29699
rect 26617 29665 26651 29699
rect 31953 29665 31987 29699
rect 34713 29665 34747 29699
rect 1409 29597 1443 29631
rect 19625 29597 19659 29631
rect 19809 29597 19843 29631
rect 21557 29597 21591 29631
rect 21649 29597 21683 29631
rect 22109 29597 22143 29631
rect 22753 29597 22787 29631
rect 23489 29597 23523 29631
rect 23673 29597 23707 29631
rect 24409 29597 24443 29631
rect 25329 29597 25363 29631
rect 25605 29597 25639 29631
rect 26893 29597 26927 29631
rect 28825 29597 28859 29631
rect 29009 29597 29043 29631
rect 29561 29597 29595 29631
rect 31677 29599 31711 29633
rect 31861 29597 31895 29631
rect 32045 29597 32079 29631
rect 32229 29597 32263 29631
rect 32873 29597 32907 29631
rect 33057 29597 33091 29631
rect 35725 29597 35759 29631
rect 36737 29597 36771 29631
rect 23029 29529 23063 29563
rect 24685 29529 24719 29563
rect 1593 29461 1627 29495
rect 18153 29461 18187 29495
rect 19717 29461 19751 29495
rect 21465 29461 21499 29495
rect 22845 29461 22879 29495
rect 25513 29461 25547 29495
rect 27997 29461 28031 29495
rect 29009 29461 29043 29495
rect 30665 29461 30699 29495
rect 32413 29461 32447 29495
rect 33517 29461 33551 29495
rect 36277 29461 36311 29495
rect 1409 29257 1443 29291
rect 19257 29257 19291 29291
rect 20729 29257 20763 29291
rect 21925 29257 21959 29291
rect 23305 29257 23339 29291
rect 23857 29257 23891 29291
rect 33793 29257 33827 29291
rect 18153 29189 18187 29223
rect 20177 29189 20211 29223
rect 25129 29189 25163 29223
rect 25329 29189 25363 29223
rect 19165 29121 19199 29155
rect 19349 29121 19383 29155
rect 19993 29121 20027 29155
rect 20637 29121 20671 29155
rect 20913 29121 20947 29155
rect 21833 29121 21867 29155
rect 22109 29121 22143 29155
rect 23029 29121 23063 29155
rect 23121 29121 23155 29155
rect 25965 29121 25999 29155
rect 26065 29121 26099 29155
rect 26985 29121 27019 29155
rect 27169 29121 27203 29155
rect 28457 29121 28491 29155
rect 28713 29121 28747 29155
rect 30757 29121 30791 29155
rect 31217 29121 31251 29155
rect 31401 29121 31435 29155
rect 32137 29121 32171 29155
rect 32689 29121 32723 29155
rect 33599 29121 33633 29155
rect 33793 29121 33827 29155
rect 34897 29121 34931 29155
rect 35265 29121 35299 29155
rect 35817 29121 35851 29155
rect 36001 29121 36035 29155
rect 17601 29053 17635 29087
rect 23305 29053 23339 29087
rect 24501 29053 24535 29087
rect 26157 29053 26191 29087
rect 26249 29053 26283 29087
rect 34345 29053 34379 29087
rect 36093 29053 36127 29087
rect 36461 29053 36495 29087
rect 18705 28985 18739 29019
rect 22201 28985 22235 29019
rect 27629 28985 27663 29019
rect 29837 28985 29871 29019
rect 31493 28985 31527 29019
rect 19809 28917 19843 28951
rect 20913 28917 20947 28951
rect 22293 28917 22327 28951
rect 22569 28917 22603 28951
rect 24961 28917 24995 28951
rect 25145 28917 25179 28951
rect 25789 28917 25823 28951
rect 26985 28917 27019 28951
rect 32229 28917 32263 28951
rect 18521 28713 18555 28747
rect 21281 28713 21315 28747
rect 28273 28713 28307 28747
rect 30481 28713 30515 28747
rect 35817 28713 35851 28747
rect 19717 28645 19751 28679
rect 29561 28645 29595 28679
rect 36645 28645 36679 28679
rect 37197 28645 37231 28679
rect 18705 28577 18739 28611
rect 20453 28577 20487 28611
rect 21373 28577 21407 28611
rect 25053 28577 25087 28611
rect 25237 28577 25271 28611
rect 27813 28577 27847 28611
rect 28733 28577 28767 28611
rect 32505 28577 32539 28611
rect 33241 28577 33275 28611
rect 34069 28577 34103 28611
rect 18429 28509 18463 28543
rect 19533 28509 19567 28543
rect 19625 28509 19659 28543
rect 19809 28509 19843 28543
rect 20821 28509 20855 28543
rect 21281 28509 21315 28543
rect 22109 28509 22143 28543
rect 22293 28509 22327 28543
rect 22569 28509 22603 28543
rect 25145 28509 25179 28543
rect 25329 28509 25363 28543
rect 27546 28509 27580 28543
rect 28457 28509 28491 28543
rect 28641 28509 28675 28543
rect 29837 28509 29871 28543
rect 30297 28509 30331 28543
rect 32249 28509 32283 28543
rect 32965 28509 32999 28543
rect 33977 28509 34011 28543
rect 34161 28509 34195 28543
rect 34988 28509 35022 28543
rect 35081 28509 35115 28543
rect 35173 28509 35207 28543
rect 35357 28509 35391 28543
rect 36185 28509 36219 28543
rect 37749 28509 37783 28543
rect 18705 28441 18739 28475
rect 20637 28441 20671 28475
rect 22753 28441 22787 28475
rect 23213 28441 23247 28475
rect 23397 28441 23431 28475
rect 29561 28441 29595 28475
rect 34713 28441 34747 28475
rect 36001 28441 36035 28475
rect 19349 28373 19383 28407
rect 21649 28373 21683 28407
rect 23581 28373 23615 28407
rect 24869 28373 24903 28407
rect 26433 28373 26467 28407
rect 29745 28373 29779 28407
rect 31125 28373 31159 28407
rect 19717 28169 19751 28203
rect 20913 28169 20947 28203
rect 23213 28169 23247 28203
rect 23949 28169 23983 28203
rect 25329 28169 25363 28203
rect 26341 28169 26375 28203
rect 27813 28169 27847 28203
rect 30481 28169 30515 28203
rect 31585 28169 31619 28203
rect 35541 28169 35575 28203
rect 36277 28169 36311 28203
rect 37841 28169 37875 28203
rect 19257 28101 19291 28135
rect 20545 28101 20579 28135
rect 20745 28101 20779 28135
rect 22201 28101 22235 28135
rect 24133 28101 24167 28135
rect 25513 28101 25547 28135
rect 27077 28101 27111 28135
rect 28733 28101 28767 28135
rect 28917 28101 28951 28135
rect 31217 28101 31251 28135
rect 31309 28101 31343 28135
rect 35081 28101 35115 28135
rect 19901 28033 19935 28067
rect 22017 28033 22051 28067
rect 22293 28033 22327 28067
rect 23121 28033 23155 28067
rect 23397 28033 23431 28067
rect 23857 28033 23891 28067
rect 24593 28033 24627 28067
rect 24685 28033 24719 28067
rect 26985 28033 27019 28067
rect 27261 28033 27295 28067
rect 28089 28033 28123 28067
rect 30113 28033 30147 28067
rect 30941 28033 30975 28067
rect 31089 28033 31123 28067
rect 31447 28033 31481 28067
rect 32321 28033 32355 28067
rect 32781 28033 32815 28067
rect 32965 28033 32999 28067
rect 35541 28033 35575 28067
rect 35725 28033 35759 28067
rect 36185 28033 36219 28067
rect 36369 28033 36403 28067
rect 18705 27965 18739 27999
rect 20085 27965 20119 27999
rect 24869 27965 24903 27999
rect 27813 27965 27847 27999
rect 27997 27965 28031 27999
rect 30021 27965 30055 27999
rect 34253 27965 34287 27999
rect 53389 27965 53423 27999
rect 53665 27965 53699 27999
rect 23397 27897 23431 27931
rect 24133 27897 24167 27931
rect 25881 27897 25915 27931
rect 27261 27897 27295 27931
rect 37289 27897 37323 27931
rect 20729 27829 20763 27863
rect 21833 27829 21867 27863
rect 24777 27829 24811 27863
rect 25513 27829 25547 27863
rect 28549 27829 28583 27863
rect 29469 27829 29503 27863
rect 19533 27625 19567 27659
rect 21649 27625 21683 27659
rect 27905 27625 27939 27659
rect 31309 27625 31343 27659
rect 36461 27625 36495 27659
rect 37013 27625 37047 27659
rect 37565 27625 37599 27659
rect 53665 27625 53699 27659
rect 19901 27557 19935 27591
rect 22937 27557 22971 27591
rect 25605 27557 25639 27591
rect 25881 27557 25915 27591
rect 26341 27557 26375 27591
rect 29009 27557 29043 27591
rect 29653 27557 29687 27591
rect 31493 27557 31527 27591
rect 21465 27489 21499 27523
rect 23765 27489 23799 27523
rect 24685 27489 24719 27523
rect 25513 27489 25547 27523
rect 30205 27489 30239 27523
rect 30665 27489 30699 27523
rect 31953 27489 31987 27523
rect 34805 27489 34839 27523
rect 1685 27421 1719 27455
rect 19533 27421 19567 27455
rect 19717 27421 19751 27455
rect 20729 27421 20763 27455
rect 21373 27421 21407 27455
rect 22753 27421 22787 27455
rect 24593 27421 24627 27455
rect 25237 27421 25271 27455
rect 25421 27421 25455 27455
rect 25697 27421 25731 27455
rect 26525 27421 26559 27455
rect 26617 27421 26651 27455
rect 28365 27421 28399 27455
rect 28733 27421 28767 27455
rect 28825 27421 28859 27455
rect 30297 27421 30331 27455
rect 32137 27421 32171 27455
rect 32689 27421 32723 27455
rect 33793 27421 33827 27455
rect 35357 27421 35391 27455
rect 2237 27353 2271 27387
rect 22385 27353 22419 27387
rect 22661 27353 22695 27387
rect 28503 27353 28537 27387
rect 28641 27353 28675 27387
rect 31125 27353 31159 27387
rect 1501 27285 1535 27319
rect 22569 27285 22603 27319
rect 27169 27285 27203 27319
rect 31325 27285 31359 27319
rect 35909 27285 35943 27319
rect 20361 27081 20395 27115
rect 22661 27081 22695 27115
rect 24317 27081 24351 27115
rect 25513 27081 25547 27115
rect 26157 27081 26191 27115
rect 28641 27081 28675 27115
rect 29561 27081 29595 27115
rect 30389 27081 30423 27115
rect 31493 27081 31527 27115
rect 32597 27081 32631 27115
rect 19901 27013 19935 27047
rect 21281 27013 21315 27047
rect 23213 27013 23247 27047
rect 25329 27013 25363 27047
rect 32229 27013 32263 27047
rect 32413 27013 32447 27047
rect 34897 27013 34931 27047
rect 21005 26945 21039 26979
rect 21097 26945 21131 26979
rect 22201 26945 22235 26979
rect 22293 26945 22327 26979
rect 22477 26945 22511 26979
rect 24225 26945 24259 26979
rect 24409 26945 24443 26979
rect 25145 26945 25179 26979
rect 26249 26945 26283 26979
rect 26433 26945 26467 26979
rect 27445 26945 27479 26979
rect 27905 26945 27939 26979
rect 27997 26945 28031 26979
rect 28181 26945 28215 26979
rect 29377 26945 29411 26979
rect 30113 26945 30147 26979
rect 30849 26945 30883 26979
rect 31033 26945 31067 26979
rect 33149 26945 33183 26979
rect 33977 26945 34011 26979
rect 35725 26945 35759 26979
rect 21281 26877 21315 26911
rect 22385 26877 22419 26911
rect 23765 26877 23799 26911
rect 26985 26877 27019 26911
rect 29193 26877 29227 26911
rect 30389 26877 30423 26911
rect 34069 26877 34103 26911
rect 28181 26809 28215 26843
rect 30849 26809 30883 26843
rect 25973 26741 26007 26775
rect 27169 26741 27203 26775
rect 30205 26741 30239 26775
rect 36185 26741 36219 26775
rect 22109 26537 22143 26571
rect 24501 26537 24535 26571
rect 25973 26537 26007 26571
rect 27629 26537 27663 26571
rect 28181 26537 28215 26571
rect 29009 26537 29043 26571
rect 30389 26537 30423 26571
rect 30757 26537 30791 26571
rect 32505 26537 32539 26571
rect 34069 26537 34103 26571
rect 20453 26469 20487 26503
rect 22753 26469 22787 26503
rect 19993 26401 20027 26435
rect 21925 26401 21959 26435
rect 25513 26401 25547 26435
rect 26157 26401 26191 26435
rect 26433 26401 26467 26435
rect 30481 26401 30515 26435
rect 34805 26401 34839 26435
rect 20085 26333 20119 26367
rect 21833 26333 21867 26367
rect 22661 26333 22695 26367
rect 22845 26333 22879 26367
rect 24409 26333 24443 26367
rect 24593 26333 24627 26367
rect 26249 26333 26283 26367
rect 26341 26333 26375 26367
rect 26985 26333 27019 26367
rect 27077 26333 27111 26367
rect 27460 26333 27494 26367
rect 28089 26333 28123 26367
rect 28273 26333 28307 26367
rect 28733 26333 28767 26367
rect 29009 26333 29043 26367
rect 29929 26333 29963 26367
rect 30389 26333 30423 26367
rect 31217 26333 31251 26367
rect 31401 26333 31435 26367
rect 31953 26333 31987 26367
rect 32965 26333 32999 26367
rect 35633 26333 35667 26367
rect 23765 26265 23799 26299
rect 27261 26265 27295 26299
rect 27353 26265 27387 26299
rect 28825 26265 28859 26299
rect 29745 26265 29779 26299
rect 33609 26265 33643 26299
rect 36093 26265 36127 26299
rect 21097 26197 21131 26231
rect 29561 26197 29595 26231
rect 31309 26197 31343 26231
rect 20085 25993 20119 26027
rect 24409 25993 24443 26027
rect 24869 25993 24903 26027
rect 26341 25993 26375 26027
rect 27537 25993 27571 26027
rect 28733 25993 28767 26027
rect 30205 25993 30239 26027
rect 32781 25993 32815 26027
rect 33333 25993 33367 26027
rect 33793 25993 33827 26027
rect 34345 25993 34379 26027
rect 24225 25925 24259 25959
rect 31033 25925 31067 25959
rect 19993 25857 20027 25891
rect 20177 25857 20211 25891
rect 20637 25857 20671 25891
rect 20821 25857 20855 25891
rect 22937 25857 22971 25891
rect 24041 25857 24075 25891
rect 24869 25857 24903 25891
rect 25053 25857 25087 25891
rect 25973 25857 26007 25891
rect 26157 25857 26191 25891
rect 27077 25857 27111 25891
rect 27997 25857 28031 25891
rect 28733 25857 28767 25891
rect 28917 25857 28951 25891
rect 29837 25857 29871 25891
rect 30021 25857 30055 25891
rect 31217 25857 31251 25891
rect 27169 25789 27203 25823
rect 27261 25789 27295 25823
rect 27353 25789 27387 25823
rect 23581 25721 23615 25755
rect 19441 25653 19475 25687
rect 20729 25653 20763 25687
rect 21833 25653 21867 25687
rect 22477 25653 22511 25687
rect 30849 25653 30883 25687
rect 32229 25653 32263 25687
rect 19993 25449 20027 25483
rect 21189 25449 21223 25483
rect 24685 25449 24719 25483
rect 25789 25449 25823 25483
rect 27169 25449 27203 25483
rect 29009 25449 29043 25483
rect 29653 25449 29687 25483
rect 32045 25449 32079 25483
rect 52837 25449 52871 25483
rect 26433 25381 26467 25415
rect 32597 25381 32631 25415
rect 20177 25313 20211 25347
rect 20729 25313 20763 25347
rect 27629 25313 27663 25347
rect 30481 25313 30515 25347
rect 19717 25245 19751 25279
rect 19809 25245 19843 25279
rect 20821 25245 20855 25279
rect 26341 25245 26375 25279
rect 26525 25245 26559 25279
rect 26985 25245 27019 25279
rect 27169 25245 27203 25279
rect 28825 25245 28859 25279
rect 29009 25245 29043 25279
rect 29561 25245 29595 25279
rect 29745 25245 29779 25279
rect 30389 25245 30423 25279
rect 30849 25245 30883 25279
rect 31309 25245 31343 25279
rect 31493 25245 31527 25279
rect 53389 25245 53423 25279
rect 1869 25177 1903 25211
rect 1961 25109 1995 25143
rect 21741 25109 21775 25143
rect 22937 25109 22971 25143
rect 25145 25109 25179 25143
rect 28273 25109 28307 25143
rect 30205 25109 30239 25143
rect 31309 25109 31343 25143
rect 53573 25109 53607 25143
rect 1685 24905 1719 24939
rect 19901 24905 19935 24939
rect 21833 24905 21867 24939
rect 24593 24905 24627 24939
rect 25145 24905 25179 24939
rect 25973 24905 26007 24939
rect 29193 24905 29227 24939
rect 29653 24905 29687 24939
rect 32229 24905 32263 24939
rect 20085 24769 20119 24803
rect 20269 24769 20303 24803
rect 20913 24769 20947 24803
rect 21281 24769 21315 24803
rect 21833 24769 21867 24803
rect 22017 24769 22051 24803
rect 27077 24769 27111 24803
rect 30021 24769 30055 24803
rect 31033 24769 31067 24803
rect 21097 24701 21131 24735
rect 29929 24701 29963 24735
rect 30941 24701 30975 24735
rect 21189 24633 21223 24667
rect 30665 24633 30699 24667
rect 19349 24565 19383 24599
rect 27629 24565 27663 24599
rect 28089 24565 28123 24599
rect 20085 24361 20119 24395
rect 21373 24361 21407 24395
rect 26801 24361 26835 24395
rect 27353 24361 27387 24395
rect 30481 24361 30515 24395
rect 20913 24293 20947 24327
rect 22109 24225 22143 24259
rect 22661 24225 22695 24259
rect 30113 24225 30147 24259
rect 21373 24157 21407 24191
rect 21557 24157 21591 24191
rect 30205 24157 30239 24191
rect 19533 24089 19567 24123
rect 20545 24089 20579 24123
rect 20729 24089 20763 24123
rect 31033 24021 31067 24055
rect 20821 23817 20855 23851
rect 30021 23817 30055 23851
rect 52837 23817 52871 23851
rect 20637 23681 20671 23715
rect 20821 23681 20855 23715
rect 53389 23681 53423 23715
rect 21833 23613 21867 23647
rect 20085 23477 20119 23511
rect 53573 23477 53607 23511
rect 20913 23273 20947 23307
rect 1409 22593 1443 22627
rect 1685 22525 1719 22559
rect 1409 22185 1443 22219
rect 53389 21505 53423 21539
rect 52837 21369 52871 21403
rect 53573 21301 53607 21335
rect 1409 20893 1443 20927
rect 1593 20757 1627 20791
rect 1409 20485 1443 20519
rect 53389 18649 53423 18683
rect 53573 18649 53607 18683
rect 52929 18581 52963 18615
rect 1869 18241 1903 18275
rect 2145 18037 2179 18071
rect 1593 17765 1627 17799
rect 52837 16609 52871 16643
rect 53389 16541 53423 16575
rect 53573 16405 53607 16439
rect 1409 16065 1443 16099
rect 1593 15861 1627 15895
rect 1409 15657 1443 15691
rect 1685 13889 1719 13923
rect 2237 13889 2271 13923
rect 52929 13889 52963 13923
rect 53665 13889 53699 13923
rect 53481 13753 53515 13787
rect 1501 13685 1535 13719
rect 53389 11713 53423 11747
rect 52837 11577 52871 11611
rect 53573 11577 53607 11611
rect 1869 11033 1903 11067
rect 2237 11033 2271 11067
rect 1593 10761 1627 10795
rect 53389 9945 53423 9979
rect 53573 9945 53607 9979
rect 52929 9877 52963 9911
rect 1685 8925 1719 8959
rect 2237 8857 2271 8891
rect 1501 8789 1535 8823
rect 1869 7361 1903 7395
rect 52929 7361 52963 7395
rect 53665 7361 53699 7395
rect 53481 7225 53515 7259
rect 1961 7157 1995 7191
rect 1685 6953 1719 6987
rect 53389 5185 53423 5219
rect 52837 5049 52871 5083
rect 53573 4981 53607 5015
rect 1685 4573 1719 4607
rect 2237 4573 2271 4607
rect 1501 4437 1535 4471
rect 53389 3485 53423 3519
rect 52837 3417 52871 3451
rect 1593 3349 1627 3383
rect 2145 3349 2179 3383
rect 53573 3349 53607 3383
rect 51457 3145 51491 3179
rect 1869 3009 1903 3043
rect 53389 3009 53423 3043
rect 2145 2941 2179 2975
rect 13461 2873 13495 2907
rect 52837 2873 52871 2907
rect 2789 2805 2823 2839
rect 6469 2805 6503 2839
rect 19349 2805 19383 2839
rect 22109 2805 22143 2839
rect 32229 2805 32263 2839
rect 34897 2805 34931 2839
rect 45109 2805 45143 2839
rect 47777 2805 47811 2839
rect 50353 2805 50387 2839
rect 52193 2805 52227 2839
rect 53573 2805 53607 2839
rect 2145 2601 2179 2635
rect 22385 2601 22419 2635
rect 25973 2601 26007 2635
rect 50721 2601 50755 2635
rect 6745 2533 6779 2567
rect 15117 2533 15151 2567
rect 24593 2533 24627 2567
rect 32505 2533 32539 2567
rect 35357 2533 35391 2567
rect 38945 2533 38979 2567
rect 41613 2533 41647 2567
rect 53297 2533 53331 2567
rect 2973 2465 3007 2499
rect 10977 2465 11011 2499
rect 11529 2465 11563 2499
rect 19717 2465 19751 2499
rect 30665 2465 30699 2499
rect 2789 2397 2823 2431
rect 4261 2397 4295 2431
rect 6561 2397 6595 2431
rect 8953 2397 8987 2431
rect 10701 2397 10735 2431
rect 13277 2397 13311 2431
rect 14473 2397 14507 2431
rect 14933 2397 14967 2431
rect 17141 2397 17175 2431
rect 19441 2397 19475 2431
rect 22293 2397 22327 2431
rect 24409 2397 24443 2431
rect 29929 2397 29963 2431
rect 30389 2397 30423 2431
rect 32321 2397 32355 2431
rect 36737 2397 36771 2431
rect 37565 2397 37599 2431
rect 38301 2397 38335 2431
rect 38761 2397 38795 2431
rect 43269 2397 43303 2431
rect 45201 2397 45235 2431
rect 50629 2397 50663 2431
rect 51641 2397 51675 2431
rect 1869 2329 1903 2363
rect 25421 2329 25455 2363
rect 26065 2329 26099 2363
rect 27353 2329 27387 2363
rect 27905 2329 27939 2363
rect 28089 2329 28123 2363
rect 35173 2329 35207 2363
rect 40877 2329 40911 2363
rect 41429 2329 41463 2363
rect 48053 2329 48087 2363
rect 53573 2329 53607 2363
rect 4077 2261 4111 2295
rect 4813 2261 4847 2295
rect 8401 2261 8435 2295
rect 9137 2261 9171 2295
rect 13093 2261 13127 2295
rect 16957 2261 16991 2295
rect 17693 2261 17727 2295
rect 23857 2261 23891 2295
rect 37381 2261 37415 2295
rect 42809 2261 42843 2295
rect 43453 2261 43487 2295
rect 45385 2261 45419 2295
rect 48145 2261 48179 2295
rect 51825 2261 51859 2295
<< metal1 >>
rect 1104 54970 54372 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 54372 54970
rect 1104 54896 54372 54918
rect 5810 54816 5816 54868
rect 5868 54856 5874 54868
rect 6457 54859 6515 54865
rect 6457 54856 6469 54859
rect 5868 54828 6469 54856
rect 5868 54816 5874 54828
rect 6457 54825 6469 54828
rect 6503 54825 6515 54859
rect 6457 54819 6515 54825
rect 14182 54816 14188 54868
rect 14240 54856 14246 54868
rect 14369 54859 14427 54865
rect 14369 54856 14381 54859
rect 14240 54828 14381 54856
rect 14240 54816 14246 54828
rect 14369 54825 14381 54828
rect 14415 54825 14427 54859
rect 24670 54856 24676 54868
rect 14369 54819 14427 54825
rect 14476 54828 24676 54856
rect 14476 54788 14504 54828
rect 24670 54816 24676 54828
rect 24728 54816 24734 54868
rect 24765 54859 24823 54865
rect 24765 54825 24777 54859
rect 24811 54856 24823 54859
rect 25130 54856 25136 54868
rect 24811 54828 25136 54856
rect 24811 54825 24823 54828
rect 24765 54819 24823 54825
rect 25130 54816 25136 54828
rect 25188 54816 25194 54868
rect 29638 54816 29644 54868
rect 29696 54856 29702 54868
rect 29917 54859 29975 54865
rect 29917 54856 29929 54859
rect 29696 54828 29929 54856
rect 29696 54816 29702 54828
rect 29917 54825 29929 54828
rect 29963 54825 29975 54859
rect 29917 54819 29975 54825
rect 36078 54816 36084 54868
rect 36136 54856 36142 54868
rect 36357 54859 36415 54865
rect 36357 54856 36369 54859
rect 36136 54828 36369 54856
rect 36136 54816 36142 54828
rect 36357 54825 36369 54828
rect 36403 54825 36415 54859
rect 36357 54819 36415 54825
rect 38289 54859 38347 54865
rect 38289 54825 38301 54859
rect 38335 54856 38347 54859
rect 38654 54856 38660 54868
rect 38335 54828 38660 54856
rect 38335 54825 38347 54828
rect 38289 54819 38347 54825
rect 38654 54816 38660 54828
rect 38712 54816 38718 54868
rect 40586 54816 40592 54868
rect 40644 54856 40650 54868
rect 40865 54859 40923 54865
rect 40865 54856 40877 54859
rect 40644 54828 40877 54856
rect 40644 54816 40650 54828
rect 40865 54825 40877 54828
rect 40911 54825 40923 54859
rect 40865 54819 40923 54825
rect 47026 54816 47032 54868
rect 47084 54856 47090 54868
rect 47765 54859 47823 54865
rect 47765 54856 47777 54859
rect 47084 54828 47777 54856
rect 47084 54816 47090 54828
rect 47765 54825 47777 54828
rect 47811 54825 47823 54859
rect 47765 54819 47823 54825
rect 48593 54859 48651 54865
rect 48593 54825 48605 54859
rect 48639 54856 48651 54859
rect 48958 54856 48964 54868
rect 48639 54828 48964 54856
rect 48639 54825 48651 54828
rect 48593 54819 48651 54825
rect 48958 54816 48964 54828
rect 49016 54816 49022 54868
rect 51534 54816 51540 54868
rect 51592 54856 51598 54868
rect 51813 54859 51871 54865
rect 51813 54856 51825 54859
rect 51592 54828 51825 54856
rect 51592 54816 51598 54828
rect 51813 54825 51825 54828
rect 51859 54825 51871 54859
rect 51813 54819 51871 54825
rect 6886 54760 14504 54788
rect 3878 54680 3884 54732
rect 3936 54720 3942 54732
rect 3973 54723 4031 54729
rect 3973 54720 3985 54723
rect 3936 54692 3985 54720
rect 3936 54680 3942 54692
rect 3973 54689 3985 54692
rect 4019 54689 4031 54723
rect 3973 54683 4031 54689
rect 1394 54652 1400 54664
rect 1355 54624 1400 54652
rect 1394 54612 1400 54624
rect 1452 54612 1458 54664
rect 1670 54652 1676 54664
rect 1631 54624 1676 54652
rect 1670 54612 1676 54624
rect 1728 54612 1734 54664
rect 4249 54655 4307 54661
rect 4249 54621 4261 54655
rect 4295 54621 4307 54655
rect 6638 54652 6644 54664
rect 6599 54624 6644 54652
rect 4249 54615 4307 54621
rect 2774 54584 2780 54596
rect 2735 54556 2780 54584
rect 2774 54544 2780 54556
rect 2832 54544 2838 54596
rect 4264 54584 4292 54615
rect 6638 54612 6644 54624
rect 6696 54652 6702 54664
rect 6886 54652 6914 54760
rect 14642 54748 14648 54800
rect 14700 54788 14706 54800
rect 22186 54788 22192 54800
rect 14700 54760 22192 54788
rect 14700 54748 14706 54760
rect 22186 54748 22192 54760
rect 22244 54748 22250 54800
rect 22370 54748 22376 54800
rect 22428 54788 22434 54800
rect 25225 54791 25283 54797
rect 25225 54788 25237 54791
rect 22428 54760 25237 54788
rect 22428 54748 22434 54760
rect 25225 54757 25237 54760
rect 25271 54757 25283 54791
rect 25225 54751 25283 54757
rect 26896 54760 31754 54788
rect 10318 54680 10324 54732
rect 10376 54720 10382 54732
rect 10962 54720 10968 54732
rect 10376 54692 10968 54720
rect 10376 54680 10382 54692
rect 10962 54680 10968 54692
rect 11020 54680 11026 54732
rect 12621 54723 12679 54729
rect 12621 54689 12633 54723
rect 12667 54720 12679 54723
rect 26896 54720 26924 54760
rect 12667 54692 26924 54720
rect 27341 54723 27399 54729
rect 12667 54689 12679 54692
rect 12621 54683 12679 54689
rect 27341 54689 27353 54723
rect 27387 54720 27399 54723
rect 27706 54720 27712 54732
rect 27387 54692 27712 54720
rect 27387 54689 27399 54692
rect 27341 54683 27399 54689
rect 27706 54680 27712 54692
rect 27764 54720 27770 54732
rect 27801 54723 27859 54729
rect 27801 54720 27813 54723
rect 27764 54692 27813 54720
rect 27764 54680 27770 54692
rect 27801 54689 27813 54692
rect 27847 54689 27859 54723
rect 27801 54683 27859 54689
rect 6696 54624 6914 54652
rect 7377 54655 7435 54661
rect 6696 54612 6702 54624
rect 7377 54621 7389 54655
rect 7423 54652 7435 54655
rect 7742 54652 7748 54664
rect 7423 54624 7748 54652
rect 7423 54621 7435 54624
rect 7377 54615 7435 54621
rect 7742 54612 7748 54624
rect 7800 54652 7806 54664
rect 7837 54655 7895 54661
rect 7837 54652 7849 54655
rect 7800 54624 7849 54652
rect 7800 54612 7806 54624
rect 7837 54621 7849 54624
rect 7883 54621 7895 54655
rect 10686 54652 10692 54664
rect 10647 54624 10692 54652
rect 7837 54615 7895 54621
rect 10686 54612 10692 54624
rect 10744 54612 10750 54664
rect 11885 54655 11943 54661
rect 11885 54621 11897 54655
rect 11931 54652 11943 54655
rect 12250 54652 12256 54664
rect 11931 54624 12256 54652
rect 11931 54621 11943 54624
rect 11885 54615 11943 54621
rect 12250 54612 12256 54624
rect 12308 54652 12314 54664
rect 12437 54655 12495 54661
rect 12437 54652 12449 54655
rect 12308 54624 12449 54652
rect 12308 54612 12314 54624
rect 12437 54621 12449 54624
rect 12483 54621 12495 54655
rect 12437 54615 12495 54621
rect 14553 54655 14611 54661
rect 14553 54621 14565 54655
rect 14599 54652 14611 54655
rect 17129 54655 17187 54661
rect 14599 54624 15148 54652
rect 14599 54621 14611 54624
rect 14553 54615 14611 54621
rect 14642 54584 14648 54596
rect 4264 54556 14648 54584
rect 14642 54544 14648 54556
rect 14700 54544 14706 54596
rect 15120 54528 15148 54624
rect 17129 54621 17141 54655
rect 17175 54652 17187 54655
rect 18690 54652 18696 54664
rect 17175 54624 17724 54652
rect 18651 54624 18696 54652
rect 17175 54621 17187 54624
rect 17129 54615 17187 54621
rect 2866 54516 2872 54528
rect 2827 54488 2872 54516
rect 2866 54476 2872 54488
rect 2924 54476 2930 54528
rect 8018 54516 8024 54528
rect 7979 54488 8024 54516
rect 8018 54476 8024 54488
rect 8076 54476 8082 54528
rect 15102 54516 15108 54528
rect 15063 54488 15108 54516
rect 15102 54476 15108 54488
rect 15160 54476 15166 54528
rect 16758 54476 16764 54528
rect 16816 54516 16822 54528
rect 17696 54525 17724 54624
rect 18690 54612 18696 54624
rect 18748 54652 18754 54664
rect 19245 54655 19303 54661
rect 19245 54652 19257 54655
rect 18748 54624 19257 54652
rect 18748 54612 18754 54624
rect 19245 54621 19257 54624
rect 19291 54621 19303 54655
rect 19245 54615 19303 54621
rect 19521 54655 19579 54661
rect 19521 54621 19533 54655
rect 19567 54621 19579 54655
rect 19521 54615 19579 54621
rect 19536 54584 19564 54615
rect 21266 54612 21272 54664
rect 21324 54652 21330 54664
rect 21324 54624 22324 54652
rect 21324 54612 21330 54624
rect 22296 54596 22324 54624
rect 23198 54612 23204 54664
rect 23256 54652 23262 54664
rect 23293 54655 23351 54661
rect 23293 54652 23305 54655
rect 23256 54624 23305 54652
rect 23256 54612 23262 54624
rect 23293 54621 23305 54624
rect 23339 54621 23351 54655
rect 23293 54615 23351 54621
rect 23492 54624 24992 54652
rect 22278 54584 22284 54596
rect 19536 54556 22094 54584
rect 22239 54556 22284 54584
rect 16945 54519 17003 54525
rect 16945 54516 16957 54519
rect 16816 54488 16957 54516
rect 16816 54476 16822 54488
rect 16945 54485 16957 54488
rect 16991 54485 17003 54519
rect 16945 54479 17003 54485
rect 17681 54519 17739 54525
rect 17681 54485 17693 54519
rect 17727 54516 17739 54519
rect 18874 54516 18880 54528
rect 17727 54488 18880 54516
rect 17727 54485 17739 54488
rect 17681 54479 17739 54485
rect 18874 54476 18880 54488
rect 18932 54476 18938 54528
rect 22066 54516 22094 54556
rect 22278 54544 22284 54556
rect 22336 54544 22342 54596
rect 22465 54587 22523 54593
rect 22465 54553 22477 54587
rect 22511 54584 22523 54587
rect 23492 54584 23520 54624
rect 22511 54556 23520 54584
rect 23569 54587 23627 54593
rect 22511 54553 22523 54556
rect 22465 54547 22523 54553
rect 23569 54553 23581 54587
rect 23615 54584 23627 54587
rect 24854 54584 24860 54596
rect 23615 54556 24860 54584
rect 23615 54553 23627 54556
rect 23569 54547 23627 54553
rect 24854 54544 24860 54556
rect 24912 54544 24918 54596
rect 24964 54584 24992 54624
rect 25222 54612 25228 54664
rect 25280 54652 25286 54664
rect 25409 54655 25467 54661
rect 25409 54652 25421 54655
rect 25280 54624 25421 54652
rect 25280 54612 25286 54624
rect 25409 54621 25421 54624
rect 25455 54621 25467 54655
rect 25409 54615 25467 54621
rect 27890 54612 27896 54664
rect 27948 54652 27954 54664
rect 28077 54655 28135 54661
rect 28077 54652 28089 54655
rect 27948 54624 28089 54652
rect 27948 54612 27954 54624
rect 28077 54621 28089 54624
rect 28123 54621 28135 54655
rect 28077 54615 28135 54621
rect 28166 54612 28172 54664
rect 28224 54652 28230 54664
rect 29733 54655 29791 54661
rect 29733 54652 29745 54655
rect 28224 54624 29745 54652
rect 28224 54612 28230 54624
rect 29733 54621 29745 54624
rect 29779 54621 29791 54655
rect 30466 54652 30472 54664
rect 29733 54615 29791 54621
rect 29932 54624 30472 54652
rect 29932 54584 29960 54624
rect 30466 54612 30472 54624
rect 30524 54612 30530 54664
rect 24964 54556 29960 54584
rect 31726 54584 31754 54760
rect 33870 54720 33876 54732
rect 32324 54692 33876 54720
rect 32324 54584 32352 54692
rect 33870 54680 33876 54692
rect 33928 54680 33934 54732
rect 45094 54680 45100 54732
rect 45152 54720 45158 54732
rect 45189 54723 45247 54729
rect 45189 54720 45201 54723
rect 45152 54692 45201 54720
rect 45152 54680 45158 54692
rect 45189 54689 45201 54692
rect 45235 54689 45247 54723
rect 45189 54683 45247 54689
rect 32493 54655 32551 54661
rect 32493 54621 32505 54655
rect 32539 54652 32551 54655
rect 32674 54652 32680 54664
rect 32539 54624 32573 54652
rect 32635 54624 32680 54652
rect 32539 54621 32551 54624
rect 32493 54615 32551 54621
rect 31726 54556 32352 54584
rect 32398 54544 32404 54596
rect 32456 54584 32462 54596
rect 32508 54584 32536 54615
rect 32674 54612 32680 54624
rect 32732 54612 32738 54664
rect 36078 54612 36084 54664
rect 36136 54652 36142 54664
rect 36173 54655 36231 54661
rect 36173 54652 36185 54655
rect 36136 54624 36185 54652
rect 36136 54612 36142 54624
rect 36173 54621 36185 54624
rect 36219 54621 36231 54655
rect 36173 54615 36231 54621
rect 38654 54612 38660 54664
rect 38712 54652 38718 54664
rect 38933 54655 38991 54661
rect 38933 54652 38945 54655
rect 38712 54624 38945 54652
rect 38712 54612 38718 54624
rect 38933 54621 38945 54624
rect 38979 54621 38991 54655
rect 40681 54655 40739 54661
rect 40681 54652 40693 54655
rect 38933 54615 38991 54621
rect 40144 54624 40693 54652
rect 33137 54587 33195 54593
rect 33137 54584 33149 54587
rect 32456 54556 33149 54584
rect 32456 54544 32462 54556
rect 33137 54553 33149 54556
rect 33183 54584 33195 54587
rect 33689 54587 33747 54593
rect 33689 54584 33701 54587
rect 33183 54556 33701 54584
rect 33183 54553 33195 54556
rect 33137 54547 33195 54553
rect 33689 54553 33701 54556
rect 33735 54553 33747 54587
rect 33689 54547 33747 54553
rect 34514 54544 34520 54596
rect 34572 54584 34578 54596
rect 35253 54587 35311 54593
rect 35253 54584 35265 54587
rect 34572 54556 35265 54584
rect 34572 54544 34578 54556
rect 35253 54553 35265 54556
rect 35299 54553 35311 54587
rect 35253 54547 35311 54553
rect 40144 54528 40172 54624
rect 40681 54621 40693 54624
rect 40727 54621 40739 54655
rect 42794 54652 42800 54664
rect 42755 54624 42800 54652
rect 40681 54615 40739 54621
rect 42794 54612 42800 54624
rect 42852 54652 42858 54664
rect 43257 54655 43315 54661
rect 43257 54652 43269 54655
rect 42852 54624 43269 54652
rect 42852 54612 42858 54624
rect 43257 54621 43269 54624
rect 43303 54621 43315 54655
rect 45462 54652 45468 54664
rect 45423 54624 45468 54652
rect 43257 54615 43315 54621
rect 45462 54612 45468 54624
rect 45520 54612 45526 54664
rect 47029 54655 47087 54661
rect 47029 54621 47041 54655
rect 47075 54652 47087 54655
rect 47578 54652 47584 54664
rect 47075 54624 47584 54652
rect 47075 54621 47087 54624
rect 47029 54615 47087 54621
rect 47578 54612 47584 54624
rect 47636 54612 47642 54664
rect 48958 54612 48964 54664
rect 49016 54652 49022 54664
rect 49237 54655 49295 54661
rect 49237 54652 49249 54655
rect 49016 54624 49249 54652
rect 49016 54612 49022 54624
rect 49237 54621 49249 54624
rect 49283 54621 49295 54655
rect 49237 54615 49295 54621
rect 51169 54655 51227 54661
rect 51169 54621 51181 54655
rect 51215 54652 51227 54655
rect 51626 54652 51632 54664
rect 51215 54624 51632 54652
rect 51215 54621 51227 54624
rect 51169 54615 51227 54621
rect 51626 54612 51632 54624
rect 51684 54612 51690 54664
rect 52917 54655 52975 54661
rect 52917 54621 52929 54655
rect 52963 54652 52975 54655
rect 53377 54655 53435 54661
rect 53377 54652 53389 54655
rect 52963 54624 53389 54652
rect 52963 54621 52975 54624
rect 52917 54615 52975 54621
rect 53377 54621 53389 54624
rect 53423 54652 53435 54655
rect 53466 54652 53472 54664
rect 53423 54624 53472 54652
rect 53423 54621 53435 54624
rect 53377 54615 53435 54621
rect 53466 54612 53472 54624
rect 53524 54612 53530 54664
rect 24026 54516 24032 54528
rect 22066 54488 24032 54516
rect 24026 54476 24032 54488
rect 24084 54476 24090 54528
rect 30098 54476 30104 54528
rect 30156 54516 30162 54528
rect 30469 54519 30527 54525
rect 30469 54516 30481 54519
rect 30156 54488 30481 54516
rect 30156 54476 30162 54488
rect 30469 54485 30481 54488
rect 30515 54485 30527 54519
rect 30469 54479 30527 54485
rect 30742 54476 30748 54528
rect 30800 54516 30806 54528
rect 31021 54519 31079 54525
rect 31021 54516 31033 54519
rect 30800 54488 31033 54516
rect 30800 54476 30806 54488
rect 31021 54485 31033 54488
rect 31067 54485 31079 54519
rect 31021 54479 31079 54485
rect 32585 54519 32643 54525
rect 32585 54485 32597 54519
rect 32631 54516 32643 54519
rect 33042 54516 33048 54528
rect 32631 54488 33048 54516
rect 32631 54485 32643 54488
rect 32585 54479 32643 54485
rect 33042 54476 33048 54488
rect 33100 54476 33106 54528
rect 34790 54476 34796 54528
rect 34848 54516 34854 54528
rect 35161 54519 35219 54525
rect 35161 54516 35173 54519
rect 34848 54488 35173 54516
rect 34848 54476 34854 54488
rect 35161 54485 35173 54488
rect 35207 54485 35219 54519
rect 38838 54516 38844 54528
rect 38799 54488 38844 54516
rect 35161 54479 35219 54485
rect 38838 54476 38844 54488
rect 38896 54476 38902 54528
rect 40126 54516 40132 54528
rect 40087 54488 40132 54516
rect 40126 54476 40132 54488
rect 40184 54476 40190 54528
rect 42610 54516 42616 54528
rect 42571 54488 42616 54516
rect 42610 54476 42616 54488
rect 42668 54476 42674 54528
rect 49142 54516 49148 54528
rect 49103 54488 49148 54516
rect 49142 54476 49148 54488
rect 49200 54476 49206 54528
rect 53561 54519 53619 54525
rect 53561 54485 53573 54519
rect 53607 54516 53619 54519
rect 53650 54516 53656 54528
rect 53607 54488 53656 54516
rect 53607 54485 53619 54488
rect 53561 54479 53619 54485
rect 53650 54476 53656 54488
rect 53708 54476 53714 54528
rect 1104 54426 54372 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 54372 54426
rect 1104 54352 54372 54374
rect 2593 54315 2651 54321
rect 2593 54281 2605 54315
rect 2639 54312 2651 54315
rect 2774 54312 2780 54324
rect 2639 54284 2780 54312
rect 2639 54281 2651 54284
rect 2593 54275 2651 54281
rect 2774 54272 2780 54284
rect 2832 54272 2838 54324
rect 3878 54312 3884 54324
rect 3839 54284 3884 54312
rect 3878 54272 3884 54284
rect 3936 54272 3942 54324
rect 6638 54272 6644 54324
rect 6696 54312 6702 54324
rect 6733 54315 6791 54321
rect 6733 54312 6745 54315
rect 6696 54284 6745 54312
rect 6696 54272 6702 54284
rect 6733 54281 6745 54284
rect 6779 54281 6791 54315
rect 6733 54275 6791 54281
rect 10962 54272 10968 54324
rect 11020 54312 11026 54324
rect 11517 54315 11575 54321
rect 11517 54312 11529 54315
rect 11020 54284 11529 54312
rect 11020 54272 11026 54284
rect 11517 54281 11529 54284
rect 11563 54281 11575 54315
rect 11517 54275 11575 54281
rect 22097 54315 22155 54321
rect 22097 54281 22109 54315
rect 22143 54312 22155 54315
rect 22278 54312 22284 54324
rect 22143 54284 22284 54312
rect 22143 54281 22155 54284
rect 22097 54275 22155 54281
rect 22278 54272 22284 54284
rect 22336 54272 22342 54324
rect 23198 54312 23204 54324
rect 23159 54284 23204 54312
rect 23198 54272 23204 54284
rect 23256 54272 23262 54324
rect 24670 54272 24676 54324
rect 24728 54312 24734 54324
rect 31386 54312 31392 54324
rect 24728 54284 31392 54312
rect 24728 54272 24734 54284
rect 31386 54272 31392 54284
rect 31444 54272 31450 54324
rect 34514 54272 34520 54324
rect 34572 54312 34578 54324
rect 34885 54315 34943 54321
rect 34885 54312 34897 54315
rect 34572 54284 34897 54312
rect 34572 54272 34578 54284
rect 34885 54281 34897 54284
rect 34931 54281 34943 54315
rect 40126 54312 40132 54324
rect 34885 54275 34943 54281
rect 35866 54284 40132 54312
rect 1302 54204 1308 54256
rect 1360 54244 1366 54256
rect 1857 54247 1915 54253
rect 1857 54244 1869 54247
rect 1360 54216 1869 54244
rect 1360 54204 1366 54216
rect 1857 54213 1869 54216
rect 1903 54213 1915 54247
rect 1857 54207 1915 54213
rect 22186 54204 22192 54256
rect 22244 54244 22250 54256
rect 30377 54247 30435 54253
rect 30377 54244 30389 54247
rect 22244 54216 30389 54244
rect 22244 54204 22250 54216
rect 30377 54213 30389 54216
rect 30423 54244 30435 54247
rect 30558 54244 30564 54256
rect 30423 54216 30564 54244
rect 30423 54213 30435 54216
rect 30377 54207 30435 54213
rect 30558 54204 30564 54216
rect 30616 54204 30622 54256
rect 31202 54204 31208 54256
rect 31260 54244 31266 54256
rect 35866 54244 35894 54284
rect 40126 54272 40132 54284
rect 40184 54272 40190 54324
rect 45094 54312 45100 54324
rect 45055 54284 45100 54312
rect 45094 54272 45100 54284
rect 45152 54272 45158 54324
rect 31260 54216 35894 54244
rect 52917 54247 52975 54253
rect 31260 54204 31266 54216
rect 52917 54213 52929 54247
rect 52963 54244 52975 54247
rect 53558 54244 53564 54256
rect 52963 54216 53564 54244
rect 52963 54213 52975 54216
rect 52917 54207 52975 54213
rect 53558 54204 53564 54216
rect 53616 54204 53622 54256
rect 28097 54179 28155 54185
rect 28097 54145 28109 54179
rect 28143 54176 28155 54179
rect 28258 54176 28264 54188
rect 28143 54148 28264 54176
rect 28143 54145 28155 54148
rect 28097 54139 28155 54145
rect 28258 54136 28264 54148
rect 28316 54136 28322 54188
rect 29365 54179 29423 54185
rect 29365 54145 29377 54179
rect 29411 54145 29423 54179
rect 29365 54139 29423 54145
rect 15102 54068 15108 54120
rect 15160 54108 15166 54120
rect 28353 54111 28411 54117
rect 15160 54080 27016 54108
rect 15160 54068 15166 54080
rect 2041 54043 2099 54049
rect 2041 54009 2053 54043
rect 2087 54040 2099 54043
rect 2130 54040 2136 54052
rect 2087 54012 2136 54040
rect 2087 54009 2099 54012
rect 2041 54003 2099 54009
rect 2130 54000 2136 54012
rect 2188 54000 2194 54052
rect 26988 53984 27016 54080
rect 28353 54077 28365 54111
rect 28399 54077 28411 54111
rect 29380 54108 29408 54139
rect 29454 54136 29460 54188
rect 29512 54176 29518 54188
rect 29549 54179 29607 54185
rect 29549 54176 29561 54179
rect 29512 54148 29561 54176
rect 29512 54136 29518 54148
rect 29549 54145 29561 54148
rect 29595 54145 29607 54179
rect 30576 54176 30604 54204
rect 31389 54179 31447 54185
rect 31389 54176 31401 54179
rect 30576 54148 31401 54176
rect 29549 54139 29607 54145
rect 31389 54145 31401 54148
rect 31435 54145 31447 54179
rect 31389 54139 31447 54145
rect 32585 54179 32643 54185
rect 32585 54145 32597 54179
rect 32631 54176 32643 54179
rect 32674 54176 32680 54188
rect 32631 54148 32680 54176
rect 32631 54145 32643 54148
rect 32585 54139 32643 54145
rect 30098 54108 30104 54120
rect 29380 54080 30104 54108
rect 28353 54071 28411 54077
rect 24854 53932 24860 53984
rect 24912 53972 24918 53984
rect 25958 53972 25964 53984
rect 24912 53944 25964 53972
rect 24912 53932 24918 53944
rect 25958 53932 25964 53944
rect 26016 53932 26022 53984
rect 26970 53972 26976 53984
rect 26931 53944 26976 53972
rect 26970 53932 26976 53944
rect 27028 53932 27034 53984
rect 28074 53932 28080 53984
rect 28132 53972 28138 53984
rect 28368 53972 28396 54071
rect 30098 54068 30104 54080
rect 30156 54068 30162 54120
rect 31938 54068 31944 54120
rect 31996 54108 32002 54120
rect 32398 54108 32404 54120
rect 31996 54080 32404 54108
rect 31996 54068 32002 54080
rect 32398 54068 32404 54080
rect 32456 54068 32462 54120
rect 32600 54108 32628 54139
rect 32674 54136 32680 54148
rect 32732 54136 32738 54188
rect 33042 54136 33048 54188
rect 33100 54176 33106 54188
rect 33229 54179 33287 54185
rect 33229 54176 33241 54179
rect 33100 54148 33241 54176
rect 33100 54136 33106 54148
rect 33229 54145 33241 54148
rect 33275 54145 33287 54179
rect 33229 54139 33287 54145
rect 33318 54136 33324 54188
rect 33376 54176 33382 54188
rect 33413 54179 33471 54185
rect 33413 54176 33425 54179
rect 33376 54148 33425 54176
rect 33376 54136 33382 54148
rect 33413 54145 33425 54148
rect 33459 54145 33471 54179
rect 33413 54139 33471 54145
rect 32600 54080 33364 54108
rect 33336 54040 33364 54080
rect 42610 54040 42616 54052
rect 33336 54012 42616 54040
rect 42610 54000 42616 54012
rect 42668 54000 42674 54052
rect 53374 54040 53380 54052
rect 53335 54012 53380 54040
rect 53374 54000 53380 54012
rect 53432 54000 53438 54052
rect 28902 53972 28908 53984
rect 28132 53944 28396 53972
rect 28863 53944 28908 53972
rect 28132 53932 28138 53944
rect 28902 53932 28908 53944
rect 28960 53932 28966 53984
rect 29457 53975 29515 53981
rect 29457 53941 29469 53975
rect 29503 53972 29515 53975
rect 29546 53972 29552 53984
rect 29503 53944 29552 53972
rect 29503 53941 29515 53944
rect 29457 53935 29515 53941
rect 29546 53932 29552 53944
rect 29604 53932 29610 53984
rect 30742 53932 30748 53984
rect 30800 53972 30806 53984
rect 30837 53975 30895 53981
rect 30837 53972 30849 53975
rect 30800 53944 30849 53972
rect 30800 53932 30806 53944
rect 30837 53941 30849 53944
rect 30883 53941 30895 53975
rect 30837 53935 30895 53941
rect 32214 53932 32220 53984
rect 32272 53972 32278 53984
rect 32769 53975 32827 53981
rect 32769 53972 32781 53975
rect 32272 53944 32781 53972
rect 32272 53932 32278 53944
rect 32769 53941 32781 53944
rect 32815 53972 32827 53975
rect 33226 53972 33232 53984
rect 32815 53944 33232 53972
rect 32815 53941 32827 53944
rect 32769 53935 32827 53941
rect 33226 53932 33232 53944
rect 33284 53932 33290 53984
rect 33410 53972 33416 53984
rect 33371 53944 33416 53972
rect 33410 53932 33416 53944
rect 33468 53932 33474 53984
rect 36078 53972 36084 53984
rect 36039 53944 36084 53972
rect 36078 53932 36084 53944
rect 36136 53932 36142 53984
rect 1104 53882 54372 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 54372 53882
rect 1104 53808 54372 53830
rect 1302 53728 1308 53780
rect 1360 53768 1366 53780
rect 1581 53771 1639 53777
rect 1581 53768 1593 53771
rect 1360 53740 1593 53768
rect 1360 53728 1366 53740
rect 1581 53737 1593 53740
rect 1627 53737 1639 53771
rect 31294 53768 31300 53780
rect 1581 53731 1639 53737
rect 29932 53740 31300 53768
rect 29454 53592 29460 53644
rect 29512 53632 29518 53644
rect 29549 53635 29607 53641
rect 29549 53632 29561 53635
rect 29512 53604 29561 53632
rect 29512 53592 29518 53604
rect 29549 53601 29561 53604
rect 29595 53601 29607 53635
rect 29549 53595 29607 53601
rect 26881 53567 26939 53573
rect 26881 53533 26893 53567
rect 26927 53564 26939 53567
rect 28074 53564 28080 53576
rect 26927 53536 28080 53564
rect 26927 53533 26939 53536
rect 26881 53527 26939 53533
rect 28074 53524 28080 53536
rect 28132 53524 28138 53576
rect 29932 53573 29960 53740
rect 31294 53728 31300 53740
rect 31352 53768 31358 53780
rect 33410 53768 33416 53780
rect 31352 53740 33416 53768
rect 31352 53728 31358 53740
rect 31386 53700 31392 53712
rect 31347 53672 31392 53700
rect 31386 53660 31392 53672
rect 31444 53660 31450 53712
rect 33244 53709 33272 53740
rect 33410 53728 33416 53740
rect 33468 53768 33474 53780
rect 34422 53768 34428 53780
rect 33468 53740 34428 53768
rect 33468 53728 33474 53740
rect 34422 53728 34428 53740
rect 34480 53728 34486 53780
rect 36170 53768 36176 53780
rect 35866 53740 36176 53768
rect 33229 53703 33287 53709
rect 33229 53669 33241 53703
rect 33275 53669 33287 53703
rect 33229 53663 33287 53669
rect 33318 53660 33324 53712
rect 33376 53700 33382 53712
rect 35866 53700 35894 53740
rect 36170 53728 36176 53740
rect 36228 53728 36234 53780
rect 33376 53672 35894 53700
rect 33376 53660 33382 53672
rect 30006 53592 30012 53644
rect 30064 53632 30070 53644
rect 30064 53604 30109 53632
rect 30064 53592 30070 53604
rect 28813 53567 28871 53573
rect 28813 53533 28825 53567
rect 28859 53533 28871 53567
rect 28813 53527 28871 53533
rect 28997 53567 29055 53573
rect 28997 53533 29009 53567
rect 29043 53564 29055 53567
rect 29917 53567 29975 53573
rect 29043 53536 29592 53564
rect 29043 53533 29055 53536
rect 28997 53527 29055 53533
rect 27154 53505 27160 53508
rect 27148 53459 27160 53505
rect 27212 53496 27218 53508
rect 28828 53496 28856 53527
rect 29564 53508 29592 53536
rect 29917 53533 29929 53567
rect 29963 53533 29975 53567
rect 30558 53564 30564 53576
rect 30519 53536 30564 53564
rect 29917 53527 29975 53533
rect 30558 53524 30564 53536
rect 30616 53524 30622 53576
rect 30742 53564 30748 53576
rect 30703 53536 30748 53564
rect 30742 53524 30748 53536
rect 30800 53524 30806 53576
rect 32122 53524 32128 53576
rect 32180 53564 32186 53576
rect 32769 53567 32827 53573
rect 32769 53564 32781 53567
rect 32180 53536 32781 53564
rect 32180 53524 32186 53536
rect 32769 53533 32781 53536
rect 32815 53533 32827 53567
rect 32769 53527 32827 53533
rect 29362 53496 29368 53508
rect 27212 53468 27248 53496
rect 28828 53468 29368 53496
rect 27154 53456 27160 53459
rect 27212 53456 27218 53468
rect 29362 53456 29368 53468
rect 29420 53456 29426 53508
rect 29546 53456 29552 53508
rect 29604 53456 29610 53508
rect 30653 53499 30711 53505
rect 30653 53465 30665 53499
rect 30699 53496 30711 53499
rect 32030 53496 32036 53508
rect 30699 53468 32036 53496
rect 30699 53465 30711 53468
rect 30653 53459 30711 53465
rect 32030 53456 32036 53468
rect 32088 53456 32094 53508
rect 32524 53499 32582 53505
rect 32524 53465 32536 53499
rect 32570 53496 32582 53499
rect 32950 53496 32956 53508
rect 32570 53468 32956 53496
rect 32570 53465 32582 53468
rect 32524 53459 32582 53465
rect 32950 53456 32956 53468
rect 33008 53456 33014 53508
rect 33597 53499 33655 53505
rect 33597 53465 33609 53499
rect 33643 53496 33655 53499
rect 34514 53496 34520 53508
rect 33643 53468 34520 53496
rect 33643 53465 33655 53468
rect 33597 53459 33655 53465
rect 34514 53456 34520 53468
rect 34572 53456 34578 53508
rect 52917 53499 52975 53505
rect 52917 53465 52929 53499
rect 52963 53496 52975 53499
rect 53558 53496 53564 53508
rect 52963 53468 53564 53496
rect 52963 53465 52975 53468
rect 52917 53459 52975 53465
rect 53558 53456 53564 53468
rect 53616 53456 53622 53508
rect 24486 53428 24492 53440
rect 24447 53400 24492 53428
rect 24486 53388 24492 53400
rect 24544 53388 24550 53440
rect 28166 53388 28172 53440
rect 28224 53428 28230 53440
rect 28261 53431 28319 53437
rect 28261 53428 28273 53431
rect 28224 53400 28273 53428
rect 28224 53388 28230 53400
rect 28261 53397 28273 53400
rect 28307 53397 28319 53431
rect 28810 53428 28816 53440
rect 28771 53400 28816 53428
rect 28261 53391 28319 53397
rect 28810 53388 28816 53400
rect 28868 53388 28874 53440
rect 31662 53388 31668 53440
rect 31720 53428 31726 53440
rect 33413 53431 33471 53437
rect 33413 53428 33425 53431
rect 31720 53400 33425 53428
rect 31720 53388 31726 53400
rect 33413 53397 33425 53400
rect 33459 53397 33471 53431
rect 33413 53391 33471 53397
rect 33502 53388 33508 53440
rect 33560 53428 33566 53440
rect 33778 53428 33784 53440
rect 33560 53400 33605 53428
rect 33739 53400 33784 53428
rect 33560 53388 33566 53400
rect 33778 53388 33784 53400
rect 33836 53388 33842 53440
rect 52454 53388 52460 53440
rect 52512 53428 52518 53440
rect 53469 53431 53527 53437
rect 53469 53428 53481 53431
rect 52512 53400 53481 53428
rect 52512 53388 52518 53400
rect 53469 53397 53481 53400
rect 53515 53397 53527 53431
rect 53469 53391 53527 53397
rect 1104 53338 54372 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 54372 53338
rect 1104 53264 54372 53286
rect 1394 53224 1400 53236
rect 1355 53196 1400 53224
rect 1394 53184 1400 53196
rect 1452 53184 1458 53236
rect 24486 53184 24492 53236
rect 24544 53224 24550 53236
rect 24949 53227 25007 53233
rect 24949 53224 24961 53227
rect 24544 53196 24961 53224
rect 24544 53184 24550 53196
rect 24949 53193 24961 53196
rect 24995 53224 25007 53227
rect 24995 53196 29684 53224
rect 24995 53193 25007 53196
rect 24949 53187 25007 53193
rect 24504 53156 24532 53184
rect 23860 53128 24532 53156
rect 29656 53156 29684 53196
rect 31386 53184 31392 53236
rect 31444 53224 31450 53236
rect 33318 53224 33324 53236
rect 31444 53196 33324 53224
rect 31444 53184 31450 53196
rect 33318 53184 33324 53196
rect 33376 53184 33382 53236
rect 33502 53184 33508 53236
rect 33560 53224 33566 53236
rect 33689 53227 33747 53233
rect 33689 53224 33701 53227
rect 33560 53196 33701 53224
rect 33560 53184 33566 53196
rect 33689 53193 33701 53196
rect 33735 53224 33747 53227
rect 34146 53224 34152 53236
rect 33735 53196 34152 53224
rect 33735 53193 33747 53196
rect 33689 53187 33747 53193
rect 34146 53184 34152 53196
rect 34204 53184 34210 53236
rect 34422 53224 34428 53236
rect 34383 53196 34428 53224
rect 34422 53184 34428 53196
rect 34480 53184 34486 53236
rect 45462 53156 45468 53168
rect 29656 53128 45468 53156
rect 23860 53097 23888 53128
rect 45462 53116 45468 53128
rect 45520 53116 45526 53168
rect 23845 53091 23903 53097
rect 23845 53057 23857 53091
rect 23891 53057 23903 53091
rect 24026 53088 24032 53100
rect 23987 53060 24032 53088
rect 23845 53051 23903 53057
rect 24026 53048 24032 53060
rect 24084 53048 24090 53100
rect 27893 53091 27951 53097
rect 27893 53057 27905 53091
rect 27939 53088 27951 53091
rect 28810 53088 28816 53100
rect 27939 53060 28816 53088
rect 27939 53057 27951 53060
rect 27893 53051 27951 53057
rect 28810 53048 28816 53060
rect 28868 53048 28874 53100
rect 31205 53091 31263 53097
rect 31205 53057 31217 53091
rect 31251 53088 31263 53091
rect 31662 53088 31668 53100
rect 31251 53060 31668 53088
rect 31251 53057 31263 53060
rect 31205 53051 31263 53057
rect 31662 53048 31668 53060
rect 31720 53048 31726 53100
rect 32030 53048 32036 53100
rect 32088 53088 32094 53100
rect 32125 53091 32183 53097
rect 32125 53088 32137 53091
rect 32088 53060 32137 53088
rect 32088 53048 32094 53060
rect 32125 53057 32137 53060
rect 32171 53057 32183 53091
rect 32125 53051 32183 53057
rect 33413 53091 33471 53097
rect 33413 53057 33425 53091
rect 33459 53088 33471 53091
rect 34238 53088 34244 53100
rect 33459 53060 34244 53088
rect 33459 53057 33471 53060
rect 33413 53051 33471 53057
rect 34238 53048 34244 53060
rect 34296 53048 34302 53100
rect 34330 53048 34336 53100
rect 34388 53088 34394 53100
rect 34609 53091 34667 53097
rect 34388 53060 34433 53088
rect 34388 53048 34394 53060
rect 34609 53057 34621 53091
rect 34655 53057 34667 53091
rect 34609 53051 34667 53057
rect 52917 53091 52975 53097
rect 52917 53057 52929 53091
rect 52963 53088 52975 53091
rect 53653 53091 53711 53097
rect 53653 53088 53665 53091
rect 52963 53060 53665 53088
rect 52963 53057 52975 53060
rect 52917 53051 52975 53057
rect 53653 53057 53665 53060
rect 53699 53088 53711 53091
rect 55398 53088 55404 53100
rect 53699 53060 55404 53088
rect 53699 53057 53711 53060
rect 53653 53051 53711 53057
rect 27982 53020 27988 53032
rect 27943 52992 27988 53020
rect 27982 52980 27988 52992
rect 28040 52980 28046 53032
rect 28074 52980 28080 53032
rect 28132 53020 28138 53032
rect 28721 53023 28779 53029
rect 28721 53020 28733 53023
rect 28132 52992 28733 53020
rect 28132 52980 28138 52992
rect 28721 52989 28733 52992
rect 28767 52989 28779 53023
rect 28994 53020 29000 53032
rect 28955 52992 29000 53020
rect 28721 52983 28779 52989
rect 28994 52980 29000 52992
rect 29052 52980 29058 53032
rect 31297 53023 31355 53029
rect 31297 52989 31309 53023
rect 31343 53020 31355 53023
rect 31478 53020 31484 53032
rect 31343 52992 31484 53020
rect 31343 52989 31355 52992
rect 31297 52983 31355 52989
rect 31478 52980 31484 52992
rect 31536 52980 31542 53032
rect 33502 53020 33508 53032
rect 33463 52992 33508 53020
rect 33502 52980 33508 52992
rect 33560 52980 33566 53032
rect 33781 53023 33839 53029
rect 33781 52989 33793 53023
rect 33827 52989 33839 53023
rect 33781 52983 33839 52989
rect 33873 53023 33931 53029
rect 33873 52989 33885 53023
rect 33919 53020 33931 53023
rect 34514 53020 34520 53032
rect 33919 52992 34520 53020
rect 33919 52989 33931 52992
rect 33873 52983 33931 52989
rect 30834 52952 30840 52964
rect 30795 52924 30840 52952
rect 30834 52912 30840 52924
rect 30892 52912 30898 52964
rect 32585 52955 32643 52961
rect 32585 52921 32597 52955
rect 32631 52952 32643 52955
rect 33796 52952 33824 52983
rect 34514 52980 34520 52992
rect 34572 52980 34578 53032
rect 34624 52952 34652 53051
rect 55398 53048 55404 53060
rect 55456 53048 55462 53100
rect 32631 52924 34652 52952
rect 32631 52921 32643 52924
rect 32585 52915 32643 52921
rect 23842 52884 23848 52896
rect 23803 52856 23848 52884
rect 23842 52844 23848 52856
rect 23900 52844 23906 52896
rect 26234 52884 26240 52896
rect 26147 52856 26240 52884
rect 26234 52844 26240 52856
rect 26292 52884 26298 52896
rect 26973 52887 27031 52893
rect 26973 52884 26985 52887
rect 26292 52856 26985 52884
rect 26292 52844 26298 52856
rect 26973 52853 26985 52856
rect 27019 52853 27031 52887
rect 26973 52847 27031 52853
rect 28261 52887 28319 52893
rect 28261 52853 28273 52887
rect 28307 52884 28319 52887
rect 28718 52884 28724 52896
rect 28307 52856 28724 52884
rect 28307 52853 28319 52856
rect 28261 52847 28319 52853
rect 28718 52844 28724 52856
rect 28776 52844 28782 52896
rect 30098 52884 30104 52896
rect 30059 52856 30104 52884
rect 30098 52844 30104 52856
rect 30156 52844 30162 52896
rect 32214 52884 32220 52896
rect 32175 52856 32220 52884
rect 32214 52844 32220 52856
rect 32272 52844 32278 52896
rect 33229 52887 33287 52893
rect 33229 52853 33241 52887
rect 33275 52884 33287 52887
rect 33502 52884 33508 52896
rect 33275 52856 33508 52884
rect 33275 52853 33287 52856
rect 33229 52847 33287 52853
rect 33502 52844 33508 52856
rect 33560 52844 33566 52896
rect 33686 52844 33692 52896
rect 33744 52884 33750 52896
rect 34793 52887 34851 52893
rect 34793 52884 34805 52887
rect 33744 52856 34805 52884
rect 33744 52844 33750 52856
rect 34793 52853 34805 52856
rect 34839 52853 34851 52887
rect 34793 52847 34851 52853
rect 35345 52887 35403 52893
rect 35345 52853 35357 52887
rect 35391 52884 35403 52887
rect 35618 52884 35624 52896
rect 35391 52856 35624 52884
rect 35391 52853 35403 52856
rect 35345 52847 35403 52853
rect 35618 52844 35624 52856
rect 35676 52844 35682 52896
rect 53282 52844 53288 52896
rect 53340 52884 53346 52896
rect 53469 52887 53527 52893
rect 53469 52884 53481 52887
rect 53340 52856 53481 52884
rect 53340 52844 53346 52856
rect 53469 52853 53481 52856
rect 53515 52853 53527 52887
rect 53469 52847 53527 52853
rect 1104 52794 54372 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 54372 52794
rect 1104 52720 54372 52742
rect 28994 52680 29000 52692
rect 28955 52652 29000 52680
rect 28994 52640 29000 52652
rect 29052 52640 29058 52692
rect 31481 52683 31539 52689
rect 31481 52649 31493 52683
rect 31527 52680 31539 52683
rect 31662 52680 31668 52692
rect 31527 52652 31668 52680
rect 31527 52649 31539 52652
rect 31481 52643 31539 52649
rect 31662 52640 31668 52652
rect 31720 52640 31726 52692
rect 34238 52640 34244 52692
rect 34296 52680 34302 52692
rect 35342 52680 35348 52692
rect 34296 52652 35348 52680
rect 34296 52640 34302 52652
rect 35342 52640 35348 52652
rect 35400 52640 35406 52692
rect 1581 52615 1639 52621
rect 1581 52581 1593 52615
rect 1627 52612 1639 52615
rect 1946 52612 1952 52624
rect 1627 52584 1952 52612
rect 1627 52581 1639 52584
rect 1581 52575 1639 52581
rect 1946 52572 1952 52584
rect 2004 52572 2010 52624
rect 24026 52572 24032 52624
rect 24084 52612 24090 52624
rect 27982 52612 27988 52624
rect 24084 52584 24808 52612
rect 24084 52572 24090 52584
rect 24780 52553 24808 52584
rect 26620 52584 27568 52612
rect 27895 52584 27988 52612
rect 24397 52547 24455 52553
rect 24397 52544 24409 52547
rect 23676 52516 24409 52544
rect 1394 52476 1400 52488
rect 1355 52448 1400 52476
rect 1394 52436 1400 52448
rect 1452 52436 1458 52488
rect 23474 52436 23480 52488
rect 23532 52476 23538 52488
rect 23676 52485 23704 52516
rect 24397 52513 24409 52516
rect 24443 52513 24455 52547
rect 24397 52507 24455 52513
rect 24765 52547 24823 52553
rect 24765 52513 24777 52547
rect 24811 52513 24823 52547
rect 25590 52544 25596 52556
rect 25551 52516 25596 52544
rect 24765 52507 24823 52513
rect 25590 52504 25596 52516
rect 25648 52504 25654 52556
rect 26053 52547 26111 52553
rect 26053 52513 26065 52547
rect 26099 52513 26111 52547
rect 26053 52507 26111 52513
rect 23661 52479 23719 52485
rect 23661 52476 23673 52479
rect 23532 52448 23673 52476
rect 23532 52436 23538 52448
rect 23661 52445 23673 52448
rect 23707 52445 23719 52479
rect 23842 52476 23848 52488
rect 23803 52448 23848 52476
rect 23661 52439 23719 52445
rect 23842 52436 23848 52448
rect 23900 52436 23906 52488
rect 24486 52436 24492 52488
rect 24544 52476 24550 52488
rect 24581 52479 24639 52485
rect 24581 52476 24593 52479
rect 24544 52448 24593 52476
rect 24544 52436 24550 52448
rect 24581 52445 24593 52448
rect 24627 52445 24639 52479
rect 24581 52439 24639 52445
rect 25685 52479 25743 52485
rect 25685 52445 25697 52479
rect 25731 52445 25743 52479
rect 26068 52476 26096 52507
rect 26142 52504 26148 52556
rect 26200 52544 26206 52556
rect 26620 52553 26648 52584
rect 26605 52547 26663 52553
rect 26605 52544 26617 52547
rect 26200 52516 26617 52544
rect 26200 52504 26206 52516
rect 26605 52513 26617 52516
rect 26651 52513 26663 52547
rect 26605 52507 26663 52513
rect 27540 52485 27568 52584
rect 27982 52572 27988 52584
rect 28040 52612 28046 52624
rect 32493 52615 32551 52621
rect 28040 52584 30052 52612
rect 28040 52572 28046 52584
rect 29546 52544 29552 52556
rect 29507 52516 29552 52544
rect 29546 52504 29552 52516
rect 29604 52504 29610 52556
rect 30024 52553 30052 52584
rect 32493 52581 32505 52615
rect 32539 52612 32551 52615
rect 32539 52584 35020 52612
rect 32539 52581 32551 52584
rect 32493 52575 32551 52581
rect 30009 52547 30067 52553
rect 30009 52513 30021 52547
rect 30055 52513 30067 52547
rect 30009 52507 30067 52513
rect 31849 52547 31907 52553
rect 31849 52513 31861 52547
rect 31895 52544 31907 52547
rect 32030 52544 32036 52556
rect 31895 52516 32036 52544
rect 31895 52513 31907 52516
rect 31849 52507 31907 52513
rect 32030 52504 32036 52516
rect 32088 52504 32094 52556
rect 33042 52544 33048 52556
rect 32416 52516 33048 52544
rect 26697 52479 26755 52485
rect 26697 52476 26709 52479
rect 26068 52448 26709 52476
rect 25685 52439 25743 52445
rect 26697 52445 26709 52448
rect 26743 52476 26755 52479
rect 27525 52479 27583 52485
rect 26743 52448 27476 52476
rect 26743 52445 26755 52448
rect 26697 52439 26755 52445
rect 25700 52408 25728 52439
rect 26234 52408 26240 52420
rect 25700 52380 26240 52408
rect 26234 52368 26240 52380
rect 26292 52368 26298 52420
rect 27448 52408 27476 52448
rect 27525 52445 27537 52479
rect 27571 52445 27583 52479
rect 27525 52439 27583 52445
rect 27617 52479 27675 52485
rect 27617 52445 27629 52479
rect 27663 52445 27675 52479
rect 27617 52439 27675 52445
rect 27632 52408 27660 52439
rect 27706 52436 27712 52488
rect 27764 52476 27770 52488
rect 27801 52479 27859 52485
rect 27801 52476 27813 52479
rect 27764 52448 27813 52476
rect 27764 52436 27770 52448
rect 27801 52445 27813 52448
rect 27847 52445 27859 52479
rect 28718 52476 28724 52488
rect 28679 52448 28724 52476
rect 27801 52439 27859 52445
rect 28718 52436 28724 52448
rect 28776 52436 28782 52488
rect 28810 52436 28816 52488
rect 28868 52476 28874 52488
rect 28868 52448 28913 52476
rect 28868 52436 28874 52448
rect 29362 52436 29368 52488
rect 29420 52476 29426 52488
rect 29822 52476 29828 52488
rect 29420 52448 29828 52476
rect 29420 52436 29426 52448
rect 29822 52436 29828 52448
rect 29880 52476 29886 52488
rect 29917 52479 29975 52485
rect 29917 52476 29929 52479
rect 29880 52448 29929 52476
rect 29880 52436 29886 52448
rect 29917 52445 29929 52448
rect 29963 52445 29975 52479
rect 29917 52439 29975 52445
rect 30193 52479 30251 52485
rect 30193 52445 30205 52479
rect 30239 52476 30251 52479
rect 30282 52476 30288 52488
rect 30239 52448 30288 52476
rect 30239 52445 30251 52448
rect 30193 52439 30251 52445
rect 30282 52436 30288 52448
rect 30340 52436 30346 52488
rect 30558 52436 30564 52488
rect 30616 52476 30622 52488
rect 32416 52485 32444 52516
rect 33042 52504 33048 52516
rect 33100 52504 33106 52556
rect 33321 52547 33379 52553
rect 33321 52513 33333 52547
rect 33367 52544 33379 52547
rect 33594 52544 33600 52556
rect 33367 52516 33600 52544
rect 33367 52513 33379 52516
rect 33321 52507 33379 52513
rect 33594 52504 33600 52516
rect 33652 52504 33658 52556
rect 34992 52553 35020 52584
rect 34977 52547 35035 52553
rect 34977 52513 34989 52547
rect 35023 52513 35035 52547
rect 34977 52507 35035 52513
rect 30653 52479 30711 52485
rect 30653 52476 30665 52479
rect 30616 52448 30665 52476
rect 30616 52436 30622 52448
rect 30653 52445 30665 52448
rect 30699 52445 30711 52479
rect 30653 52439 30711 52445
rect 31021 52479 31079 52485
rect 31021 52445 31033 52479
rect 31067 52476 31079 52479
rect 31665 52479 31723 52485
rect 31665 52476 31677 52479
rect 31067 52448 31677 52476
rect 31067 52445 31079 52448
rect 31021 52439 31079 52445
rect 31665 52445 31677 52448
rect 31711 52476 31723 52479
rect 32401 52479 32459 52485
rect 32401 52476 32413 52479
rect 31711 52448 32413 52476
rect 31711 52445 31723 52448
rect 31665 52439 31723 52445
rect 32401 52445 32413 52448
rect 32447 52445 32459 52479
rect 32401 52439 32459 52445
rect 32585 52479 32643 52485
rect 32585 52445 32597 52479
rect 32631 52476 32643 52479
rect 33870 52476 33876 52488
rect 32631 52448 33088 52476
rect 33810 52448 33876 52476
rect 32631 52445 32643 52448
rect 32585 52439 32643 52445
rect 28994 52408 29000 52420
rect 27448 52380 27660 52408
rect 28955 52380 29000 52408
rect 28994 52368 29000 52380
rect 29052 52368 29058 52420
rect 30742 52368 30748 52420
rect 30800 52408 30806 52420
rect 30837 52411 30895 52417
rect 30837 52408 30849 52411
rect 30800 52380 30849 52408
rect 30800 52368 30806 52380
rect 30837 52377 30849 52380
rect 30883 52377 30895 52411
rect 33060 52408 33088 52448
rect 33870 52436 33876 52448
rect 33928 52476 33934 52488
rect 34146 52476 34152 52488
rect 33928 52448 34008 52476
rect 34059 52448 34152 52476
rect 33928 52436 33934 52448
rect 33060 52380 33180 52408
rect 30837 52371 30895 52377
rect 23753 52343 23811 52349
rect 23753 52309 23765 52343
rect 23799 52340 23811 52343
rect 23842 52340 23848 52352
rect 23799 52312 23848 52340
rect 23799 52309 23811 52312
rect 23753 52303 23811 52309
rect 23842 52300 23848 52312
rect 23900 52300 23906 52352
rect 27065 52343 27123 52349
rect 27065 52309 27077 52343
rect 27111 52340 27123 52343
rect 27338 52340 27344 52352
rect 27111 52312 27344 52340
rect 27111 52309 27123 52312
rect 27065 52303 27123 52309
rect 27338 52300 27344 52312
rect 27396 52300 27402 52352
rect 33152 52340 33180 52380
rect 33318 52368 33324 52420
rect 33376 52408 33382 52420
rect 33980 52408 34008 52448
rect 34146 52436 34152 52448
rect 34204 52476 34210 52488
rect 35069 52479 35127 52485
rect 35069 52476 35081 52479
rect 34204 52448 35081 52476
rect 34204 52436 34210 52448
rect 35069 52445 35081 52448
rect 35115 52445 35127 52479
rect 35069 52439 35127 52445
rect 35710 52408 35716 52420
rect 33376 52380 35716 52408
rect 33376 52368 33382 52380
rect 35710 52368 35716 52380
rect 35768 52368 35774 52420
rect 33686 52340 33692 52352
rect 33152 52312 33692 52340
rect 33686 52300 33692 52312
rect 33744 52300 33750 52352
rect 34606 52300 34612 52352
rect 34664 52340 34670 52352
rect 34701 52343 34759 52349
rect 34701 52340 34713 52343
rect 34664 52312 34713 52340
rect 34664 52300 34670 52312
rect 34701 52309 34713 52312
rect 34747 52309 34759 52343
rect 34701 52303 34759 52309
rect 35894 52300 35900 52352
rect 35952 52340 35958 52352
rect 36265 52343 36323 52349
rect 36265 52340 36277 52343
rect 35952 52312 36277 52340
rect 35952 52300 35958 52312
rect 36265 52309 36277 52312
rect 36311 52309 36323 52343
rect 36265 52303 36323 52309
rect 1104 52250 54372 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 54372 52250
rect 1104 52176 54372 52198
rect 1394 52136 1400 52148
rect 1355 52108 1400 52136
rect 1394 52096 1400 52108
rect 1452 52096 1458 52148
rect 25133 52139 25191 52145
rect 25133 52105 25145 52139
rect 25179 52136 25191 52139
rect 25590 52136 25596 52148
rect 25179 52108 25596 52136
rect 25179 52105 25191 52108
rect 25133 52099 25191 52105
rect 25590 52096 25596 52108
rect 25648 52096 25654 52148
rect 26421 52139 26479 52145
rect 26421 52105 26433 52139
rect 26467 52136 26479 52139
rect 27706 52136 27712 52148
rect 26467 52108 27712 52136
rect 26467 52105 26479 52108
rect 26421 52099 26479 52105
rect 27706 52096 27712 52108
rect 27764 52096 27770 52148
rect 29822 52136 29828 52148
rect 29783 52108 29828 52136
rect 29822 52096 29828 52108
rect 29880 52096 29886 52148
rect 31294 52136 31300 52148
rect 31255 52108 31300 52136
rect 31294 52096 31300 52108
rect 31352 52096 31358 52148
rect 33410 52096 33416 52148
rect 33468 52136 33474 52148
rect 35342 52136 35348 52148
rect 33468 52108 33548 52136
rect 35303 52108 35348 52136
rect 33468 52096 33474 52108
rect 23474 52068 23480 52080
rect 23400 52040 23480 52068
rect 23400 52009 23428 52040
rect 23474 52028 23480 52040
rect 23532 52028 23538 52080
rect 23750 52068 23756 52080
rect 23711 52040 23756 52068
rect 23750 52028 23756 52040
rect 23808 52028 23814 52080
rect 23385 52003 23443 52009
rect 23385 51969 23397 52003
rect 23431 51969 23443 52003
rect 23566 52000 23572 52012
rect 23527 51972 23572 52000
rect 23385 51963 23443 51969
rect 23566 51960 23572 51972
rect 23624 51960 23630 52012
rect 23658 51960 23664 52012
rect 23716 52000 23722 52012
rect 23716 51972 23761 52000
rect 23716 51960 23722 51972
rect 23842 51960 23848 52012
rect 23900 52000 23906 52012
rect 24765 52003 24823 52009
rect 24765 52000 24777 52003
rect 23900 51972 24777 52000
rect 23900 51960 23906 51972
rect 24765 51969 24777 51972
rect 24811 51969 24823 52003
rect 25608 52000 25636 52096
rect 29454 52068 29460 52080
rect 29415 52040 29460 52068
rect 29454 52028 29460 52040
rect 29512 52028 29518 52080
rect 29641 52071 29699 52077
rect 29641 52037 29653 52071
rect 29687 52068 29699 52071
rect 30098 52068 30104 52080
rect 29687 52040 30104 52068
rect 29687 52037 29699 52040
rect 29641 52031 29699 52037
rect 30098 52028 30104 52040
rect 30156 52068 30162 52080
rect 30377 52071 30435 52077
rect 30377 52068 30389 52071
rect 30156 52040 30389 52068
rect 30156 52028 30162 52040
rect 30377 52037 30389 52040
rect 30423 52068 30435 52071
rect 31481 52071 31539 52077
rect 30423 52040 31340 52068
rect 30423 52037 30435 52040
rect 30377 52031 30435 52037
rect 26237 52003 26295 52009
rect 26237 52000 26249 52003
rect 25608 51972 26249 52000
rect 24765 51963 24823 51969
rect 26237 51969 26249 51972
rect 26283 51969 26295 52003
rect 26237 51963 26295 51969
rect 27341 52003 27399 52009
rect 27341 51969 27353 52003
rect 27387 52000 27399 52003
rect 27982 52000 27988 52012
rect 27387 51972 27988 52000
rect 27387 51969 27399 51972
rect 27341 51963 27399 51969
rect 27982 51960 27988 51972
rect 28040 51960 28046 52012
rect 30006 52000 30012 52012
rect 28552 51972 30012 52000
rect 23198 51892 23204 51944
rect 23256 51932 23262 51944
rect 24673 51935 24731 51941
rect 24673 51932 24685 51935
rect 23256 51904 24685 51932
rect 23256 51892 23262 51904
rect 24673 51901 24685 51904
rect 24719 51901 24731 51935
rect 24673 51895 24731 51901
rect 26053 51935 26111 51941
rect 26053 51901 26065 51935
rect 26099 51901 26111 51935
rect 27614 51932 27620 51944
rect 27575 51904 27620 51932
rect 26053 51895 26111 51901
rect 26068 51864 26096 51895
rect 27614 51892 27620 51904
rect 27672 51892 27678 51944
rect 26234 51864 26240 51876
rect 26068 51836 26240 51864
rect 26234 51824 26240 51836
rect 26292 51824 26298 51876
rect 22830 51796 22836 51808
rect 22791 51768 22836 51796
rect 22830 51756 22836 51768
rect 22888 51756 22894 51808
rect 24029 51799 24087 51805
rect 24029 51765 24041 51799
rect 24075 51796 24087 51799
rect 28552 51796 28580 51972
rect 30006 51960 30012 51972
rect 30064 52000 30070 52012
rect 31205 52003 31263 52009
rect 31205 52000 31217 52003
rect 30064 51972 31217 52000
rect 30064 51960 30070 51972
rect 31205 51969 31217 51972
rect 31251 51969 31263 52003
rect 31312 52000 31340 52040
rect 31481 52037 31493 52071
rect 31527 52068 31539 52071
rect 32214 52068 32220 52080
rect 31527 52040 32220 52068
rect 31527 52037 31539 52040
rect 31481 52031 31539 52037
rect 32214 52028 32220 52040
rect 32272 52028 32278 52080
rect 33520 52077 33548 52108
rect 35342 52096 35348 52108
rect 35400 52096 35406 52148
rect 35710 52096 35716 52148
rect 35768 52136 35774 52148
rect 36265 52139 36323 52145
rect 36265 52136 36277 52139
rect 35768 52108 36277 52136
rect 35768 52096 35774 52108
rect 36265 52105 36277 52108
rect 36311 52105 36323 52139
rect 36265 52099 36323 52105
rect 33505 52071 33563 52077
rect 33505 52037 33517 52071
rect 33551 52037 33563 52071
rect 33505 52031 33563 52037
rect 33597 52071 33655 52077
rect 33597 52037 33609 52071
rect 33643 52068 33655 52071
rect 34146 52068 34152 52080
rect 33643 52040 34152 52068
rect 33643 52037 33655 52040
rect 33597 52031 33655 52037
rect 34146 52028 34152 52040
rect 34204 52028 34210 52080
rect 31754 52000 31760 52012
rect 31312 51972 31760 52000
rect 31205 51963 31263 51969
rect 31220 51932 31248 51963
rect 31754 51960 31760 51972
rect 31812 52000 31818 52012
rect 32125 52003 32183 52009
rect 32125 52000 32137 52003
rect 31812 51972 32137 52000
rect 31812 51960 31818 51972
rect 32125 51969 32137 51972
rect 32171 51969 32183 52003
rect 32125 51963 32183 51969
rect 33318 51960 33324 52012
rect 33376 52009 33382 52012
rect 33376 52003 33425 52009
rect 33376 51969 33379 52003
rect 33413 51969 33425 52003
rect 33376 51963 33425 51969
rect 33376 51960 33382 51963
rect 33686 51960 33692 52012
rect 33744 52000 33750 52012
rect 34514 52000 34520 52012
rect 33744 51972 33789 52000
rect 34475 51972 34520 52000
rect 33744 51960 33750 51972
rect 34514 51960 34520 51972
rect 34572 51960 34578 52012
rect 35526 52000 35532 52012
rect 35487 51972 35532 52000
rect 35526 51960 35532 51972
rect 35584 51960 35590 52012
rect 33134 51932 33140 51944
rect 31220 51904 33140 51932
rect 33134 51892 33140 51904
rect 33192 51892 33198 51944
rect 33229 51935 33287 51941
rect 33229 51901 33241 51935
rect 33275 51901 33287 51935
rect 33229 51895 33287 51901
rect 33873 51935 33931 51941
rect 33873 51901 33885 51935
rect 33919 51932 33931 51935
rect 34425 51935 34483 51941
rect 34425 51932 34437 51935
rect 33919 51904 34437 51932
rect 33919 51901 33931 51904
rect 33873 51895 33931 51901
rect 34425 51901 34437 51904
rect 34471 51901 34483 51935
rect 34425 51895 34483 51901
rect 31478 51864 31484 51876
rect 31439 51836 31484 51864
rect 31478 51824 31484 51836
rect 31536 51824 31542 51876
rect 33244 51864 33272 51895
rect 35342 51892 35348 51944
rect 35400 51932 35406 51944
rect 35713 51935 35771 51941
rect 35713 51932 35725 51935
rect 35400 51904 35725 51932
rect 35400 51892 35406 51904
rect 35713 51901 35725 51904
rect 35759 51901 35771 51935
rect 35713 51895 35771 51901
rect 35805 51935 35863 51941
rect 35805 51901 35817 51935
rect 35851 51932 35863 51935
rect 35894 51932 35900 51944
rect 35851 51904 35900 51932
rect 35851 51901 35863 51904
rect 35805 51895 35863 51901
rect 35894 51892 35900 51904
rect 35952 51892 35958 51944
rect 33594 51864 33600 51876
rect 33244 51836 33600 51864
rect 33594 51824 33600 51836
rect 33652 51864 33658 51876
rect 35618 51864 35624 51876
rect 33652 51836 35624 51864
rect 33652 51824 33658 51836
rect 35618 51824 35624 51836
rect 35676 51824 35682 51876
rect 28718 51796 28724 51808
rect 24075 51768 28580 51796
rect 28679 51768 28724 51796
rect 24075 51765 24087 51768
rect 24029 51759 24087 51765
rect 28718 51756 28724 51768
rect 28776 51756 28782 51808
rect 30742 51756 30748 51808
rect 30800 51796 30806 51808
rect 32769 51799 32827 51805
rect 32769 51796 32781 51799
rect 30800 51768 32781 51796
rect 30800 51756 30806 51768
rect 32769 51765 32781 51768
rect 32815 51765 32827 51799
rect 32769 51759 32827 51765
rect 34885 51799 34943 51805
rect 34885 51765 34897 51799
rect 34931 51796 34943 51799
rect 35434 51796 35440 51808
rect 34931 51768 35440 51796
rect 34931 51765 34943 51768
rect 34885 51759 34943 51765
rect 35434 51756 35440 51768
rect 35492 51756 35498 51808
rect 37274 51796 37280 51808
rect 37235 51768 37280 51796
rect 37274 51756 37280 51768
rect 37332 51756 37338 51808
rect 1104 51706 54372 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 54372 51706
rect 1104 51632 54372 51654
rect 22189 51595 22247 51601
rect 22189 51561 22201 51595
rect 22235 51592 22247 51595
rect 22646 51592 22652 51604
rect 22235 51564 22652 51592
rect 22235 51561 22247 51564
rect 22189 51555 22247 51561
rect 22646 51552 22652 51564
rect 22704 51592 22710 51604
rect 22830 51592 22836 51604
rect 22704 51564 22836 51592
rect 22704 51552 22710 51564
rect 22830 51552 22836 51564
rect 22888 51552 22894 51604
rect 23198 51592 23204 51604
rect 23159 51564 23204 51592
rect 23198 51552 23204 51564
rect 23256 51552 23262 51604
rect 26234 51592 26240 51604
rect 26195 51564 26240 51592
rect 26234 51552 26240 51564
rect 26292 51552 26298 51604
rect 27614 51592 27620 51604
rect 27575 51564 27620 51592
rect 27614 51552 27620 51564
rect 27672 51552 27678 51604
rect 28810 51552 28816 51604
rect 28868 51592 28874 51604
rect 32582 51592 32588 51604
rect 28868 51564 32588 51592
rect 28868 51552 28874 51564
rect 32582 51552 32588 51564
rect 32640 51552 32646 51604
rect 35253 51595 35311 51601
rect 35253 51561 35265 51595
rect 35299 51592 35311 51595
rect 35526 51592 35532 51604
rect 35299 51564 35532 51592
rect 35299 51561 35311 51564
rect 35253 51555 35311 51561
rect 35526 51552 35532 51564
rect 35584 51552 35590 51604
rect 23566 51484 23572 51536
rect 23624 51524 23630 51536
rect 23842 51524 23848 51536
rect 23624 51496 23848 51524
rect 23624 51484 23630 51496
rect 23842 51484 23848 51496
rect 23900 51484 23906 51536
rect 24854 51524 24860 51536
rect 24767 51496 24860 51524
rect 24854 51484 24860 51496
rect 24912 51524 24918 51536
rect 26970 51524 26976 51536
rect 24912 51496 26976 51524
rect 24912 51484 24918 51496
rect 26970 51484 26976 51496
rect 27028 51484 27034 51536
rect 35618 51484 35624 51536
rect 35676 51524 35682 51536
rect 36265 51527 36323 51533
rect 36265 51524 36277 51527
rect 35676 51496 36277 51524
rect 35676 51484 35682 51496
rect 36265 51493 36277 51496
rect 36311 51493 36323 51527
rect 36265 51487 36323 51493
rect 22741 51459 22799 51465
rect 22741 51425 22753 51459
rect 22787 51456 22799 51459
rect 24486 51456 24492 51468
rect 22787 51428 24492 51456
rect 22787 51425 22799 51428
rect 22741 51419 22799 51425
rect 24486 51416 24492 51428
rect 24544 51416 24550 51468
rect 26881 51459 26939 51465
rect 26881 51425 26893 51459
rect 26927 51456 26939 51459
rect 30742 51456 30748 51468
rect 26927 51428 27476 51456
rect 26927 51425 26939 51428
rect 26881 51419 26939 51425
rect 23477 51391 23535 51397
rect 23477 51357 23489 51391
rect 23523 51388 23535 51391
rect 23750 51388 23756 51400
rect 23523 51360 23756 51388
rect 23523 51357 23535 51360
rect 23477 51351 23535 51357
rect 23750 51348 23756 51360
rect 23808 51348 23814 51400
rect 24946 51348 24952 51400
rect 25004 51388 25010 51400
rect 25501 51391 25559 51397
rect 25501 51388 25513 51391
rect 25004 51360 25513 51388
rect 25004 51348 25010 51360
rect 25501 51357 25513 51360
rect 25547 51357 25559 51391
rect 25501 51351 25559 51357
rect 25590 51348 25596 51400
rect 25648 51388 25654 51400
rect 25685 51391 25743 51397
rect 25685 51388 25697 51391
rect 25648 51360 25697 51388
rect 25648 51348 25654 51360
rect 25685 51357 25697 51360
rect 25731 51357 25743 51391
rect 27338 51388 27344 51400
rect 27299 51360 27344 51388
rect 25685 51351 25743 51357
rect 27338 51348 27344 51360
rect 27396 51348 27402 51400
rect 27448 51397 27476 51428
rect 30668 51428 30748 51456
rect 27433 51391 27491 51397
rect 27433 51357 27445 51391
rect 27479 51388 27491 51391
rect 28810 51388 28816 51400
rect 27479 51360 28816 51388
rect 27479 51357 27491 51360
rect 27433 51351 27491 51357
rect 28810 51348 28816 51360
rect 28868 51348 28874 51400
rect 30668 51397 30696 51428
rect 30742 51416 30748 51428
rect 30800 51416 30806 51468
rect 33321 51459 33379 51465
rect 33321 51425 33333 51459
rect 33367 51456 33379 51459
rect 36446 51456 36452 51468
rect 33367 51428 36452 51456
rect 33367 51425 33379 51428
rect 33321 51419 33379 51425
rect 36446 51416 36452 51428
rect 36504 51416 36510 51468
rect 28997 51391 29055 51397
rect 28997 51357 29009 51391
rect 29043 51388 29055 51391
rect 30653 51391 30711 51397
rect 30653 51388 30665 51391
rect 29043 51360 30665 51388
rect 29043 51357 29055 51360
rect 28997 51351 29055 51357
rect 30653 51357 30665 51360
rect 30699 51357 30711 51391
rect 30834 51388 30840 51400
rect 30795 51360 30840 51388
rect 30653 51351 30711 51357
rect 30834 51348 30840 51360
rect 30892 51348 30898 51400
rect 31294 51388 31300 51400
rect 31255 51360 31300 51388
rect 31294 51348 31300 51360
rect 31352 51348 31358 51400
rect 31481 51391 31539 51397
rect 31481 51357 31493 51391
rect 31527 51357 31539 51391
rect 33502 51388 33508 51400
rect 33463 51360 33508 51388
rect 31481 51351 31539 51357
rect 22554 51280 22560 51332
rect 22612 51320 22618 51332
rect 23201 51323 23259 51329
rect 23201 51320 23213 51323
rect 22612 51292 23213 51320
rect 22612 51280 22618 51292
rect 23201 51289 23213 51292
rect 23247 51289 23259 51323
rect 23201 51283 23259 51289
rect 23385 51323 23443 51329
rect 23385 51289 23397 51323
rect 23431 51320 23443 51323
rect 23658 51320 23664 51332
rect 23431 51292 23664 51320
rect 23431 51289 23443 51292
rect 23385 51283 23443 51289
rect 23658 51280 23664 51292
rect 23716 51280 23722 51332
rect 27246 51280 27252 51332
rect 27304 51320 27310 51332
rect 27617 51323 27675 51329
rect 27617 51320 27629 51323
rect 27304 51292 27629 51320
rect 27304 51280 27310 51292
rect 27617 51289 27629 51292
rect 27663 51289 27675 51323
rect 29549 51323 29607 51329
rect 29549 51320 29561 51323
rect 27617 51283 27675 51289
rect 28092 51292 29561 51320
rect 25685 51255 25743 51261
rect 25685 51221 25697 51255
rect 25731 51252 25743 51255
rect 26142 51252 26148 51264
rect 25731 51224 26148 51252
rect 25731 51221 25743 51224
rect 25685 51215 25743 51221
rect 26142 51212 26148 51224
rect 26200 51212 26206 51264
rect 27522 51212 27528 51264
rect 27580 51252 27586 51264
rect 28092 51261 28120 51292
rect 29549 51289 29561 51292
rect 29595 51320 29607 51323
rect 30006 51320 30012 51332
rect 29595 51292 30012 51320
rect 29595 51289 29607 51292
rect 29549 51283 29607 51289
rect 30006 51280 30012 51292
rect 30064 51280 30070 51332
rect 30745 51323 30803 51329
rect 30745 51289 30757 51323
rect 30791 51320 30803 51323
rect 31496 51320 31524 51351
rect 33502 51348 33508 51360
rect 33560 51348 33566 51400
rect 33778 51388 33784 51400
rect 33739 51360 33784 51388
rect 33778 51348 33784 51360
rect 33836 51348 33842 51400
rect 34698 51388 34704 51400
rect 34659 51360 34704 51388
rect 34698 51348 34704 51360
rect 34756 51348 34762 51400
rect 35069 51391 35127 51397
rect 35069 51357 35081 51391
rect 35115 51388 35127 51391
rect 35710 51388 35716 51400
rect 35115 51360 35716 51388
rect 35115 51357 35127 51360
rect 35069 51351 35127 51357
rect 35710 51348 35716 51360
rect 35768 51348 35774 51400
rect 30791 51292 31524 51320
rect 30791 51289 30803 51292
rect 30745 51283 30803 51289
rect 33134 51280 33140 51332
rect 33192 51320 33198 51332
rect 33689 51323 33747 51329
rect 33689 51320 33701 51323
rect 33192 51292 33701 51320
rect 33192 51280 33198 51292
rect 33689 51289 33701 51292
rect 33735 51320 33747 51323
rect 34330 51320 34336 51332
rect 33735 51292 34336 51320
rect 33735 51289 33747 51292
rect 33689 51283 33747 51289
rect 34330 51280 34336 51292
rect 34388 51280 34394 51332
rect 34882 51320 34888 51332
rect 34843 51292 34888 51320
rect 34882 51280 34888 51292
rect 34940 51280 34946 51332
rect 34977 51323 35035 51329
rect 34977 51289 34989 51323
rect 35023 51289 35035 51323
rect 34977 51283 35035 51289
rect 28077 51255 28135 51261
rect 28077 51252 28089 51255
rect 27580 51224 28089 51252
rect 27580 51212 27586 51224
rect 28077 51221 28089 51224
rect 28123 51221 28135 51255
rect 28077 51215 28135 51221
rect 29822 51212 29828 51264
rect 29880 51252 29886 51264
rect 30101 51255 30159 51261
rect 30101 51252 30113 51255
rect 29880 51224 30113 51252
rect 29880 51212 29886 51224
rect 30101 51221 30113 51224
rect 30147 51221 30159 51255
rect 31386 51252 31392 51264
rect 31347 51224 31392 51252
rect 30101 51215 30159 51221
rect 31386 51212 31392 51224
rect 31444 51212 31450 51264
rect 31938 51252 31944 51264
rect 31899 51224 31944 51252
rect 31938 51212 31944 51224
rect 31996 51212 32002 51264
rect 32582 51252 32588 51264
rect 32543 51224 32588 51252
rect 32582 51212 32588 51224
rect 32640 51212 32646 51264
rect 34992 51252 35020 51283
rect 35526 51252 35532 51264
rect 34992 51224 35532 51252
rect 35526 51212 35532 51224
rect 35584 51252 35590 51264
rect 35713 51255 35771 51261
rect 35713 51252 35725 51255
rect 35584 51224 35725 51252
rect 35584 51212 35590 51224
rect 35713 51221 35725 51224
rect 35759 51221 35771 51255
rect 35713 51215 35771 51221
rect 36909 51255 36967 51261
rect 36909 51221 36921 51255
rect 36955 51252 36967 51255
rect 37182 51252 37188 51264
rect 36955 51224 37188 51252
rect 36955 51221 36967 51224
rect 36909 51215 36967 51221
rect 37182 51212 37188 51224
rect 37240 51212 37246 51264
rect 1104 51162 54372 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 54372 51162
rect 1104 51088 54372 51110
rect 23842 51048 23848 51060
rect 23803 51020 23848 51048
rect 23842 51008 23848 51020
rect 23900 51008 23906 51060
rect 26050 51008 26056 51060
rect 26108 51048 26114 51060
rect 26145 51051 26203 51057
rect 26145 51048 26157 51051
rect 26108 51020 26157 51048
rect 26108 51008 26114 51020
rect 26145 51017 26157 51020
rect 26191 51017 26203 51051
rect 26145 51011 26203 51017
rect 31113 51051 31171 51057
rect 31113 51017 31125 51051
rect 31159 51048 31171 51051
rect 31294 51048 31300 51060
rect 31159 51020 31300 51048
rect 31159 51017 31171 51020
rect 31113 51011 31171 51017
rect 31294 51008 31300 51020
rect 31352 51008 31358 51060
rect 31754 51008 31760 51060
rect 31812 51048 31818 51060
rect 32861 51051 32919 51057
rect 32861 51048 32873 51051
rect 31812 51020 32873 51048
rect 31812 51008 31818 51020
rect 32861 51017 32873 51020
rect 32907 51017 32919 51051
rect 32861 51011 32919 51017
rect 35621 51051 35679 51057
rect 35621 51017 35633 51051
rect 35667 51048 35679 51051
rect 35710 51048 35716 51060
rect 35667 51020 35716 51048
rect 35667 51017 35679 51020
rect 35621 51011 35679 51017
rect 35710 51008 35716 51020
rect 35768 51008 35774 51060
rect 24486 50980 24492 50992
rect 23492 50952 24492 50980
rect 1394 50912 1400 50924
rect 1355 50884 1400 50912
rect 1394 50872 1400 50884
rect 1452 50872 1458 50924
rect 22554 50912 22560 50924
rect 22515 50884 22560 50912
rect 22554 50872 22560 50884
rect 22612 50872 22618 50924
rect 22738 50912 22744 50924
rect 22699 50884 22744 50912
rect 22738 50872 22744 50884
rect 22796 50872 22802 50924
rect 23198 50912 23204 50924
rect 23159 50884 23204 50912
rect 23198 50872 23204 50884
rect 23256 50872 23262 50924
rect 23492 50921 23520 50952
rect 24486 50940 24492 50952
rect 24544 50940 24550 50992
rect 30006 50980 30012 50992
rect 29967 50952 30012 50980
rect 30006 50940 30012 50952
rect 30064 50940 30070 50992
rect 30193 50983 30251 50989
rect 30193 50949 30205 50983
rect 30239 50980 30251 50983
rect 30374 50980 30380 50992
rect 30239 50952 30380 50980
rect 30239 50949 30251 50952
rect 30193 50943 30251 50949
rect 30374 50940 30380 50952
rect 30432 50940 30438 50992
rect 23385 50915 23443 50921
rect 23385 50881 23397 50915
rect 23431 50881 23443 50915
rect 23385 50875 23443 50881
rect 23477 50915 23535 50921
rect 23477 50881 23489 50915
rect 23523 50881 23535 50915
rect 23477 50875 23535 50881
rect 23569 50915 23627 50921
rect 23569 50881 23581 50915
rect 23615 50912 23627 50915
rect 23934 50912 23940 50924
rect 23615 50884 23940 50912
rect 23615 50881 23627 50884
rect 23569 50875 23627 50881
rect 23400 50776 23428 50875
rect 23934 50872 23940 50884
rect 23992 50872 23998 50924
rect 25041 50915 25099 50921
rect 25041 50881 25053 50915
rect 25087 50912 25099 50915
rect 25130 50912 25136 50924
rect 25087 50884 25136 50912
rect 25087 50881 25099 50884
rect 25041 50875 25099 50881
rect 25130 50872 25136 50884
rect 25188 50912 25194 50924
rect 25590 50912 25596 50924
rect 25188 50884 25596 50912
rect 25188 50872 25194 50884
rect 25590 50872 25596 50884
rect 25648 50872 25654 50924
rect 25866 50912 25872 50924
rect 25827 50884 25872 50912
rect 25866 50872 25872 50884
rect 25924 50872 25930 50924
rect 30282 50912 30288 50924
rect 30243 50884 30288 50912
rect 30282 50872 30288 50884
rect 30340 50872 30346 50924
rect 30834 50872 30840 50924
rect 30892 50912 30898 50924
rect 30929 50915 30987 50921
rect 30929 50912 30941 50915
rect 30892 50884 30941 50912
rect 30892 50872 30898 50884
rect 30929 50881 30941 50884
rect 30975 50881 30987 50915
rect 32398 50912 32404 50924
rect 32359 50884 32404 50912
rect 30929 50875 30987 50881
rect 32398 50872 32404 50884
rect 32456 50872 32462 50924
rect 34882 50912 34888 50924
rect 34795 50884 34888 50912
rect 34882 50872 34888 50884
rect 34940 50912 34946 50924
rect 35894 50912 35900 50924
rect 34940 50884 35900 50912
rect 34940 50872 34946 50884
rect 35894 50872 35900 50884
rect 35952 50872 35958 50924
rect 52917 50915 52975 50921
rect 52917 50881 52929 50915
rect 52963 50912 52975 50915
rect 53558 50912 53564 50924
rect 52963 50884 53564 50912
rect 52963 50881 52975 50884
rect 52917 50875 52975 50881
rect 53558 50872 53564 50884
rect 53616 50872 53622 50924
rect 24946 50844 24952 50856
rect 24907 50816 24952 50844
rect 24946 50804 24952 50816
rect 25004 50804 25010 50856
rect 26142 50844 26148 50856
rect 26103 50816 26148 50844
rect 26142 50804 26148 50816
rect 26200 50804 26206 50856
rect 30742 50844 30748 50856
rect 30703 50816 30748 50844
rect 30742 50804 30748 50816
rect 30800 50804 30806 50856
rect 32125 50847 32183 50853
rect 32125 50813 32137 50847
rect 32171 50844 32183 50847
rect 32490 50844 32496 50856
rect 32171 50816 32496 50844
rect 32171 50813 32183 50816
rect 32125 50807 32183 50813
rect 32490 50804 32496 50816
rect 32548 50804 32554 50856
rect 34514 50844 34520 50856
rect 34475 50816 34520 50844
rect 34514 50804 34520 50816
rect 34572 50804 34578 50856
rect 34698 50804 34704 50856
rect 34756 50844 34762 50856
rect 34977 50847 35035 50853
rect 34977 50844 34989 50847
rect 34756 50816 34989 50844
rect 34756 50804 34762 50816
rect 34977 50813 34989 50816
rect 35023 50844 35035 50847
rect 35342 50844 35348 50856
rect 35023 50816 35348 50844
rect 35023 50813 35035 50816
rect 34977 50807 35035 50813
rect 35342 50804 35348 50816
rect 35400 50804 35406 50856
rect 22664 50748 23428 50776
rect 25409 50779 25467 50785
rect 1581 50711 1639 50717
rect 1581 50677 1593 50711
rect 1627 50708 1639 50711
rect 1762 50708 1768 50720
rect 1627 50680 1768 50708
rect 1627 50677 1639 50680
rect 1581 50671 1639 50677
rect 1762 50668 1768 50680
rect 1820 50668 1826 50720
rect 22002 50708 22008 50720
rect 21963 50680 22008 50708
rect 22002 50668 22008 50680
rect 22060 50708 22066 50720
rect 22664 50708 22692 50748
rect 25409 50745 25421 50779
rect 25455 50776 25467 50779
rect 25774 50776 25780 50788
rect 25455 50748 25780 50776
rect 25455 50745 25467 50748
rect 25409 50739 25467 50745
rect 25774 50736 25780 50748
rect 25832 50776 25838 50788
rect 25961 50779 26019 50785
rect 25961 50776 25973 50779
rect 25832 50748 25973 50776
rect 25832 50736 25838 50748
rect 25961 50745 25973 50748
rect 26007 50745 26019 50779
rect 28445 50779 28503 50785
rect 28445 50776 28457 50779
rect 25961 50739 26019 50745
rect 27080 50748 28457 50776
rect 22060 50680 22692 50708
rect 22741 50711 22799 50717
rect 22060 50668 22066 50680
rect 22741 50677 22753 50711
rect 22787 50708 22799 50711
rect 23474 50708 23480 50720
rect 22787 50680 23480 50708
rect 22787 50677 22799 50680
rect 22741 50671 22799 50677
rect 23474 50668 23480 50680
rect 23532 50708 23538 50720
rect 23750 50708 23756 50720
rect 23532 50680 23756 50708
rect 23532 50668 23538 50680
rect 23750 50668 23756 50680
rect 23808 50668 23814 50720
rect 24026 50668 24032 50720
rect 24084 50708 24090 50720
rect 24305 50711 24363 50717
rect 24305 50708 24317 50711
rect 24084 50680 24317 50708
rect 24084 50668 24090 50680
rect 24305 50677 24317 50680
rect 24351 50677 24363 50711
rect 24305 50671 24363 50677
rect 26234 50668 26240 50720
rect 26292 50708 26298 50720
rect 26878 50708 26884 50720
rect 26292 50680 26884 50708
rect 26292 50668 26298 50680
rect 26878 50668 26884 50680
rect 26936 50708 26942 50720
rect 27080 50717 27108 50748
rect 28445 50745 28457 50748
rect 28491 50776 28503 50779
rect 28718 50776 28724 50788
rect 28491 50748 28724 50776
rect 28491 50745 28503 50748
rect 28445 50739 28503 50745
rect 28718 50736 28724 50748
rect 28776 50736 28782 50788
rect 35894 50736 35900 50788
rect 35952 50776 35958 50788
rect 36173 50779 36231 50785
rect 36173 50776 36185 50779
rect 35952 50748 36185 50776
rect 35952 50736 35958 50748
rect 36173 50745 36185 50748
rect 36219 50776 36231 50779
rect 37182 50776 37188 50788
rect 36219 50748 37188 50776
rect 36219 50745 36231 50748
rect 36173 50739 36231 50745
rect 37182 50736 37188 50748
rect 37240 50736 37246 50788
rect 27065 50711 27123 50717
rect 27065 50708 27077 50711
rect 26936 50680 27077 50708
rect 26936 50668 26942 50680
rect 27065 50677 27077 50680
rect 27111 50677 27123 50711
rect 27065 50671 27123 50677
rect 27985 50711 28043 50717
rect 27985 50677 27997 50711
rect 28031 50708 28043 50711
rect 28902 50708 28908 50720
rect 28031 50680 28908 50708
rect 28031 50677 28043 50680
rect 27985 50671 28043 50677
rect 28902 50668 28908 50680
rect 28960 50668 28966 50720
rect 29270 50668 29276 50720
rect 29328 50708 29334 50720
rect 29457 50711 29515 50717
rect 29457 50708 29469 50711
rect 29328 50680 29469 50708
rect 29328 50668 29334 50680
rect 29457 50677 29469 50680
rect 29503 50677 29515 50711
rect 29457 50671 29515 50677
rect 30009 50711 30067 50717
rect 30009 50677 30021 50711
rect 30055 50708 30067 50711
rect 30098 50708 30104 50720
rect 30055 50680 30104 50708
rect 30055 50677 30067 50680
rect 30009 50671 30067 50677
rect 30098 50668 30104 50680
rect 30156 50668 30162 50720
rect 32214 50708 32220 50720
rect 32175 50680 32220 50708
rect 32214 50668 32220 50680
rect 32272 50668 32278 50720
rect 32306 50668 32312 50720
rect 32364 50708 32370 50720
rect 33689 50711 33747 50717
rect 32364 50680 32409 50708
rect 32364 50668 32370 50680
rect 33689 50677 33701 50711
rect 33735 50708 33747 50711
rect 33778 50708 33784 50720
rect 33735 50680 33784 50708
rect 33735 50677 33747 50680
rect 33689 50671 33747 50677
rect 33778 50668 33784 50680
rect 33836 50668 33842 50720
rect 36725 50711 36783 50717
rect 36725 50677 36737 50711
rect 36771 50708 36783 50711
rect 37274 50708 37280 50720
rect 36771 50680 37280 50708
rect 36771 50677 36783 50680
rect 36725 50671 36783 50677
rect 37274 50668 37280 50680
rect 37332 50668 37338 50720
rect 53466 50708 53472 50720
rect 53427 50680 53472 50708
rect 53466 50668 53472 50680
rect 53524 50668 53530 50720
rect 1104 50618 54372 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 54372 50618
rect 1104 50544 54372 50566
rect 22554 50464 22560 50516
rect 22612 50504 22618 50516
rect 22833 50507 22891 50513
rect 22833 50504 22845 50507
rect 22612 50476 22845 50504
rect 22612 50464 22618 50476
rect 22833 50473 22845 50476
rect 22879 50473 22891 50507
rect 22833 50467 22891 50473
rect 23845 50507 23903 50513
rect 23845 50473 23857 50507
rect 23891 50504 23903 50507
rect 24946 50504 24952 50516
rect 23891 50476 24952 50504
rect 23891 50473 23903 50476
rect 23845 50467 23903 50473
rect 24946 50464 24952 50476
rect 25004 50464 25010 50516
rect 27154 50504 27160 50516
rect 27115 50476 27160 50504
rect 27154 50464 27160 50476
rect 27212 50464 27218 50516
rect 30282 50504 30288 50516
rect 30243 50476 30288 50504
rect 30282 50464 30288 50476
rect 30340 50504 30346 50516
rect 30340 50476 31524 50504
rect 30340 50464 30346 50476
rect 1394 50436 1400 50448
rect 1355 50408 1400 50436
rect 1394 50396 1400 50408
rect 1452 50396 1458 50448
rect 23474 50396 23480 50448
rect 23532 50396 23538 50448
rect 23385 50371 23443 50377
rect 23385 50337 23397 50371
rect 23431 50368 23443 50371
rect 23492 50368 23520 50396
rect 25774 50368 25780 50380
rect 23431 50340 23520 50368
rect 25735 50340 25780 50368
rect 23431 50337 23443 50340
rect 23385 50331 23443 50337
rect 25774 50328 25780 50340
rect 25832 50328 25838 50380
rect 26237 50371 26295 50377
rect 26237 50337 26249 50371
rect 26283 50368 26295 50371
rect 26510 50368 26516 50380
rect 26283 50340 26516 50368
rect 26283 50337 26295 50340
rect 26237 50331 26295 50337
rect 26510 50328 26516 50340
rect 26568 50328 26574 50380
rect 27522 50368 27528 50380
rect 26712 50340 27528 50368
rect 26712 50312 26740 50340
rect 27522 50328 27528 50340
rect 27580 50328 27586 50380
rect 28169 50371 28227 50377
rect 28169 50337 28181 50371
rect 28215 50368 28227 50371
rect 29270 50368 29276 50380
rect 28215 50340 29276 50368
rect 28215 50337 28227 50340
rect 28169 50331 28227 50337
rect 29270 50328 29276 50340
rect 29328 50328 29334 50380
rect 30374 50368 30380 50380
rect 30287 50340 30380 50368
rect 30374 50328 30380 50340
rect 30432 50368 30438 50380
rect 31018 50368 31024 50380
rect 30432 50340 31024 50368
rect 30432 50328 30438 50340
rect 31018 50328 31024 50340
rect 31076 50328 31082 50380
rect 31294 50368 31300 50380
rect 31128 50340 31300 50368
rect 20901 50303 20959 50309
rect 20901 50269 20913 50303
rect 20947 50300 20959 50303
rect 22002 50300 22008 50312
rect 20947 50272 22008 50300
rect 20947 50269 20959 50272
rect 20901 50263 20959 50269
rect 22002 50260 22008 50272
rect 22060 50300 22066 50312
rect 22465 50303 22523 50309
rect 22465 50300 22477 50303
rect 22060 50272 22477 50300
rect 22060 50260 22066 50272
rect 22465 50269 22477 50272
rect 22511 50269 22523 50303
rect 22465 50263 22523 50269
rect 22646 50260 22652 50312
rect 22704 50300 22710 50312
rect 23198 50300 23204 50312
rect 22704 50272 23204 50300
rect 22704 50260 22710 50272
rect 23198 50260 23204 50272
rect 23256 50260 23262 50312
rect 23477 50303 23535 50309
rect 23477 50269 23489 50303
rect 23523 50269 23535 50303
rect 25866 50300 25872 50312
rect 25827 50272 25872 50300
rect 23477 50263 23535 50269
rect 23492 50232 23520 50263
rect 25866 50260 25872 50272
rect 25924 50260 25930 50312
rect 26694 50300 26700 50312
rect 26655 50272 26700 50300
rect 26694 50260 26700 50272
rect 26752 50260 26758 50312
rect 26786 50260 26792 50312
rect 26844 50300 26850 50312
rect 26844 50272 26889 50300
rect 26844 50260 26850 50272
rect 26970 50260 26976 50312
rect 27028 50300 27034 50312
rect 30098 50300 30104 50312
rect 27028 50272 27073 50300
rect 30059 50272 30104 50300
rect 27028 50260 27034 50272
rect 30098 50260 30104 50272
rect 30156 50260 30162 50312
rect 31128 50309 31156 50340
rect 31294 50328 31300 50340
rect 31352 50328 31358 50380
rect 31113 50303 31171 50309
rect 31113 50269 31125 50303
rect 31159 50269 31171 50303
rect 31113 50263 31171 50269
rect 31205 50303 31263 50309
rect 31205 50269 31217 50303
rect 31251 50269 31263 50303
rect 31386 50300 31392 50312
rect 31347 50272 31392 50300
rect 31205 50263 31263 50269
rect 23566 50232 23572 50244
rect 23492 50204 23572 50232
rect 23566 50192 23572 50204
rect 23624 50192 23630 50244
rect 24854 50232 24860 50244
rect 24815 50204 24860 50232
rect 24854 50192 24860 50204
rect 24912 50192 24918 50244
rect 25041 50235 25099 50241
rect 25041 50201 25053 50235
rect 25087 50232 25099 50235
rect 25498 50232 25504 50244
rect 25087 50204 25504 50232
rect 25087 50201 25099 50204
rect 25041 50195 25099 50201
rect 21453 50167 21511 50173
rect 21453 50133 21465 50167
rect 21499 50164 21511 50167
rect 21634 50164 21640 50176
rect 21499 50136 21640 50164
rect 21499 50133 21511 50136
rect 21453 50127 21511 50133
rect 21634 50124 21640 50136
rect 21692 50124 21698 50176
rect 22005 50167 22063 50173
rect 22005 50133 22017 50167
rect 22051 50164 22063 50167
rect 24026 50164 24032 50176
rect 22051 50136 24032 50164
rect 22051 50133 22063 50136
rect 22005 50127 22063 50133
rect 24026 50124 24032 50136
rect 24084 50124 24090 50176
rect 24670 50124 24676 50176
rect 24728 50164 24734 50176
rect 25056 50164 25084 50195
rect 25498 50192 25504 50204
rect 25556 50232 25562 50244
rect 28166 50232 28172 50244
rect 25556 50204 28172 50232
rect 25556 50192 25562 50204
rect 28166 50192 28172 50204
rect 28224 50192 28230 50244
rect 31220 50232 31248 50263
rect 31386 50260 31392 50272
rect 31444 50260 31450 50312
rect 31496 50309 31524 50476
rect 32398 50464 32404 50516
rect 32456 50504 32462 50516
rect 32677 50507 32735 50513
rect 32677 50504 32689 50507
rect 32456 50476 32689 50504
rect 32456 50464 32462 50476
rect 32677 50473 32689 50476
rect 32723 50504 32735 50507
rect 34057 50507 34115 50513
rect 34057 50504 34069 50507
rect 32723 50476 34069 50504
rect 32723 50473 32735 50476
rect 32677 50467 32735 50473
rect 34057 50473 34069 50476
rect 34103 50473 34115 50507
rect 34057 50467 34115 50473
rect 37182 50464 37188 50516
rect 37240 50504 37246 50516
rect 53466 50504 53472 50516
rect 37240 50476 53472 50504
rect 37240 50464 37246 50476
rect 53466 50464 53472 50476
rect 53524 50464 53530 50516
rect 31665 50439 31723 50445
rect 31665 50405 31677 50439
rect 31711 50436 31723 50439
rect 33318 50436 33324 50448
rect 31711 50408 33324 50436
rect 31711 50405 31723 50408
rect 31665 50399 31723 50405
rect 33318 50396 33324 50408
rect 33376 50396 33382 50448
rect 34606 50368 34612 50380
rect 33336 50340 34612 50368
rect 31481 50303 31539 50309
rect 31481 50269 31493 50303
rect 31527 50269 31539 50303
rect 31481 50263 31539 50269
rect 32306 50260 32312 50312
rect 32364 50260 32370 50312
rect 32490 50300 32496 50312
rect 32451 50272 32496 50300
rect 32490 50260 32496 50272
rect 32548 50260 32554 50312
rect 33336 50309 33364 50340
rect 34606 50328 34612 50340
rect 34664 50328 34670 50380
rect 32677 50303 32735 50309
rect 32677 50269 32689 50303
rect 32723 50300 32735 50303
rect 33137 50303 33195 50309
rect 33137 50300 33149 50303
rect 32723 50272 33149 50300
rect 32723 50269 32735 50272
rect 32677 50263 32735 50269
rect 33137 50269 33149 50272
rect 33183 50269 33195 50303
rect 33137 50263 33195 50269
rect 33321 50303 33379 50309
rect 33321 50269 33333 50303
rect 33367 50269 33379 50303
rect 33321 50263 33379 50269
rect 33505 50303 33563 50309
rect 33505 50269 33517 50303
rect 33551 50300 33563 50303
rect 33778 50300 33784 50312
rect 33551 50272 33784 50300
rect 33551 50269 33563 50272
rect 33505 50263 33563 50269
rect 32324 50232 32352 50260
rect 32692 50232 32720 50263
rect 33778 50260 33784 50272
rect 33836 50260 33842 50312
rect 34146 50300 34152 50312
rect 34107 50272 34152 50300
rect 34146 50260 34152 50272
rect 34204 50260 34210 50312
rect 31220 50204 32720 50232
rect 34330 50192 34336 50244
rect 34388 50232 34394 50244
rect 53374 50232 53380 50244
rect 34388 50204 53380 50232
rect 34388 50192 34394 50204
rect 53374 50192 53380 50204
rect 53432 50192 53438 50244
rect 24728 50136 25084 50164
rect 25225 50167 25283 50173
rect 24728 50124 24734 50136
rect 25225 50133 25237 50167
rect 25271 50164 25283 50167
rect 26234 50164 26240 50176
rect 25271 50136 26240 50164
rect 25271 50133 25283 50136
rect 25225 50127 25283 50133
rect 26234 50124 26240 50136
rect 26292 50124 26298 50176
rect 28902 50164 28908 50176
rect 28863 50136 28908 50164
rect 28902 50124 28908 50136
rect 28960 50124 28966 50176
rect 29914 50164 29920 50176
rect 29875 50136 29920 50164
rect 29914 50124 29920 50136
rect 29972 50124 29978 50176
rect 31018 50124 31024 50176
rect 31076 50164 31082 50176
rect 31386 50164 31392 50176
rect 31076 50136 31392 50164
rect 31076 50124 31082 50136
rect 31386 50124 31392 50136
rect 31444 50124 31450 50176
rect 32309 50167 32367 50173
rect 32309 50133 32321 50167
rect 32355 50164 32367 50167
rect 32398 50164 32404 50176
rect 32355 50136 32404 50164
rect 32355 50133 32367 50136
rect 32309 50127 32367 50133
rect 32398 50124 32404 50136
rect 32456 50124 32462 50176
rect 34422 50124 34428 50176
rect 34480 50164 34486 50176
rect 34701 50167 34759 50173
rect 34701 50164 34713 50167
rect 34480 50136 34713 50164
rect 34480 50124 34486 50136
rect 34701 50133 34713 50136
rect 34747 50164 34759 50167
rect 35253 50167 35311 50173
rect 35253 50164 35265 50167
rect 34747 50136 35265 50164
rect 34747 50133 34759 50136
rect 34701 50127 34759 50133
rect 35253 50133 35265 50136
rect 35299 50133 35311 50167
rect 35253 50127 35311 50133
rect 35342 50124 35348 50176
rect 35400 50164 35406 50176
rect 35897 50167 35955 50173
rect 35897 50164 35909 50167
rect 35400 50136 35909 50164
rect 35400 50124 35406 50136
rect 35897 50133 35909 50136
rect 35943 50164 35955 50167
rect 37274 50164 37280 50176
rect 35943 50136 37280 50164
rect 35943 50133 35955 50136
rect 35897 50127 35955 50133
rect 37274 50124 37280 50136
rect 37332 50124 37338 50176
rect 1104 50074 54372 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 54372 50074
rect 1104 50000 54372 50022
rect 22738 49960 22744 49972
rect 22699 49932 22744 49960
rect 22738 49920 22744 49932
rect 22796 49920 22802 49972
rect 24486 49920 24492 49972
rect 24544 49960 24550 49972
rect 26421 49963 26479 49969
rect 24544 49932 24900 49960
rect 24544 49920 24550 49932
rect 21269 49895 21327 49901
rect 21269 49861 21281 49895
rect 21315 49892 21327 49895
rect 22189 49895 22247 49901
rect 22189 49892 22201 49895
rect 21315 49864 22201 49892
rect 21315 49861 21327 49864
rect 21269 49855 21327 49861
rect 22189 49861 22201 49864
rect 22235 49892 22247 49895
rect 24762 49892 24768 49904
rect 22235 49864 23704 49892
rect 22235 49861 22247 49864
rect 22189 49855 22247 49861
rect 21634 49784 21640 49836
rect 21692 49824 21698 49836
rect 22646 49824 22652 49836
rect 21692 49796 22652 49824
rect 21692 49784 21698 49796
rect 22646 49784 22652 49796
rect 22704 49784 22710 49836
rect 23676 49833 23704 49864
rect 24320 49864 24768 49892
rect 24320 49836 24348 49864
rect 24762 49852 24768 49864
rect 24820 49852 24826 49904
rect 24872 49892 24900 49932
rect 26421 49929 26433 49963
rect 26467 49960 26479 49963
rect 26786 49960 26792 49972
rect 26467 49932 26792 49960
rect 26467 49929 26479 49932
rect 26421 49923 26479 49929
rect 26786 49920 26792 49932
rect 26844 49920 26850 49972
rect 31389 49963 31447 49969
rect 26896 49932 31340 49960
rect 26896 49892 26924 49932
rect 31018 49892 31024 49904
rect 24872 49864 26924 49892
rect 30979 49864 31024 49892
rect 31018 49852 31024 49864
rect 31076 49852 31082 49904
rect 31312 49892 31340 49932
rect 31389 49929 31401 49963
rect 31435 49960 31447 49963
rect 32490 49960 32496 49972
rect 31435 49932 32496 49960
rect 31435 49929 31447 49932
rect 31389 49923 31447 49929
rect 32490 49920 32496 49932
rect 32548 49920 32554 49972
rect 34146 49920 34152 49972
rect 34204 49960 34210 49972
rect 34241 49963 34299 49969
rect 34241 49960 34253 49963
rect 34204 49932 34253 49960
rect 34204 49920 34210 49932
rect 34241 49929 34253 49932
rect 34287 49929 34299 49963
rect 34241 49923 34299 49929
rect 35161 49963 35219 49969
rect 35161 49929 35173 49963
rect 35207 49960 35219 49963
rect 52454 49960 52460 49972
rect 35207 49932 52460 49960
rect 35207 49929 35219 49932
rect 35161 49923 35219 49929
rect 31312 49864 32260 49892
rect 22833 49827 22891 49833
rect 22833 49793 22845 49827
rect 22879 49793 22891 49827
rect 22833 49787 22891 49793
rect 23661 49827 23719 49833
rect 23661 49793 23673 49827
rect 23707 49793 23719 49827
rect 23661 49787 23719 49793
rect 23845 49827 23903 49833
rect 23845 49793 23857 49827
rect 23891 49824 23903 49827
rect 24026 49824 24032 49836
rect 23891 49796 24032 49824
rect 23891 49793 23903 49796
rect 23845 49787 23903 49793
rect 22002 49716 22008 49768
rect 22060 49756 22066 49768
rect 22848 49756 22876 49787
rect 22060 49728 22876 49756
rect 23676 49756 23704 49787
rect 24026 49784 24032 49796
rect 24084 49784 24090 49836
rect 24302 49824 24308 49836
rect 24263 49796 24308 49824
rect 24302 49784 24308 49796
rect 24360 49784 24366 49836
rect 24486 49824 24492 49836
rect 24447 49796 24492 49824
rect 24486 49784 24492 49796
rect 24544 49784 24550 49836
rect 24854 49784 24860 49836
rect 24912 49824 24918 49836
rect 25317 49827 25375 49833
rect 25317 49824 25329 49827
rect 24912 49796 25329 49824
rect 24912 49784 24918 49796
rect 25317 49793 25329 49796
rect 25363 49793 25375 49827
rect 25498 49824 25504 49836
rect 25459 49796 25504 49824
rect 25317 49787 25375 49793
rect 25498 49784 25504 49796
rect 25556 49784 25562 49836
rect 26234 49824 26240 49836
rect 26195 49796 26240 49824
rect 26234 49784 26240 49796
rect 26292 49784 26298 49836
rect 29730 49824 29736 49836
rect 29788 49833 29794 49836
rect 29700 49796 29736 49824
rect 29730 49784 29736 49796
rect 29788 49787 29800 49833
rect 29788 49784 29794 49787
rect 30282 49784 30288 49836
rect 30340 49824 30346 49836
rect 30929 49827 30987 49833
rect 30929 49824 30941 49827
rect 30340 49796 30941 49824
rect 30340 49784 30346 49796
rect 30929 49793 30941 49796
rect 30975 49793 30987 49827
rect 30929 49787 30987 49793
rect 31205 49827 31263 49833
rect 31205 49793 31217 49827
rect 31251 49824 31263 49827
rect 31294 49824 31300 49836
rect 31251 49796 31300 49824
rect 31251 49793 31263 49796
rect 31205 49787 31263 49793
rect 31294 49784 31300 49796
rect 31352 49784 31358 49836
rect 32122 49824 32128 49836
rect 32083 49796 32128 49824
rect 32122 49784 32128 49796
rect 32180 49784 32186 49836
rect 32232 49824 32260 49864
rect 33778 49852 33784 49904
rect 33836 49892 33842 49904
rect 34422 49892 34428 49904
rect 33836 49864 34428 49892
rect 33836 49852 33842 49864
rect 34422 49852 34428 49864
rect 34480 49852 34486 49904
rect 34606 49892 34612 49904
rect 34567 49864 34612 49892
rect 34606 49852 34612 49864
rect 34664 49852 34670 49904
rect 34330 49824 34336 49836
rect 32232 49796 34336 49824
rect 34330 49784 34336 49796
rect 34388 49784 34394 49836
rect 24504 49756 24532 49784
rect 23676 49728 24532 49756
rect 25409 49759 25467 49765
rect 22060 49716 22066 49728
rect 23860 49700 23888 49728
rect 25409 49725 25421 49759
rect 25455 49756 25467 49759
rect 25866 49756 25872 49768
rect 25455 49728 25872 49756
rect 25455 49725 25467 49728
rect 25409 49719 25467 49725
rect 25866 49716 25872 49728
rect 25924 49756 25930 49768
rect 26053 49759 26111 49765
rect 26053 49756 26065 49759
rect 25924 49728 26065 49756
rect 25924 49716 25930 49728
rect 26053 49725 26065 49728
rect 26099 49725 26111 49759
rect 26053 49719 26111 49725
rect 27065 49759 27123 49765
rect 27065 49725 27077 49759
rect 27111 49756 27123 49759
rect 27614 49756 27620 49768
rect 27111 49728 27620 49756
rect 27111 49725 27123 49728
rect 27065 49719 27123 49725
rect 27614 49716 27620 49728
rect 27672 49716 27678 49768
rect 28074 49756 28080 49768
rect 28035 49728 28080 49756
rect 28074 49716 28080 49728
rect 28132 49716 28138 49768
rect 30006 49716 30012 49768
rect 30064 49756 30070 49768
rect 32140 49756 32168 49784
rect 30064 49728 32168 49756
rect 32401 49759 32459 49765
rect 30064 49716 30070 49728
rect 32401 49725 32413 49759
rect 32447 49756 32459 49759
rect 32582 49756 32588 49768
rect 32447 49728 32588 49756
rect 32447 49725 32459 49728
rect 32401 49719 32459 49725
rect 32582 49716 32588 49728
rect 32640 49716 32646 49768
rect 33042 49716 33048 49768
rect 33100 49756 33106 49768
rect 35176 49756 35204 49923
rect 52454 49920 52460 49932
rect 52512 49920 52518 49972
rect 33100 49728 35204 49756
rect 33100 49716 33106 49728
rect 36906 49716 36912 49768
rect 36964 49756 36970 49768
rect 37274 49756 37280 49768
rect 36964 49728 37280 49756
rect 36964 49716 36970 49728
rect 37274 49716 37280 49728
rect 37332 49716 37338 49768
rect 23842 49648 23848 49700
rect 23900 49648 23906 49700
rect 23474 49580 23480 49632
rect 23532 49620 23538 49632
rect 23753 49623 23811 49629
rect 23753 49620 23765 49623
rect 23532 49592 23765 49620
rect 23532 49580 23538 49592
rect 23753 49589 23765 49592
rect 23799 49589 23811 49623
rect 23753 49583 23811 49589
rect 24397 49623 24455 49629
rect 24397 49589 24409 49623
rect 24443 49620 24455 49623
rect 24486 49620 24492 49632
rect 24443 49592 24492 49620
rect 24443 49589 24455 49592
rect 24397 49583 24455 49589
rect 24486 49580 24492 49592
rect 24544 49580 24550 49632
rect 28629 49623 28687 49629
rect 28629 49589 28641 49623
rect 28675 49620 28687 49623
rect 29362 49620 29368 49632
rect 28675 49592 29368 49620
rect 28675 49589 28687 49592
rect 28629 49583 28687 49589
rect 29362 49580 29368 49592
rect 29420 49620 29426 49632
rect 30742 49620 30748 49632
rect 29420 49592 30748 49620
rect 29420 49580 29426 49592
rect 30742 49580 30748 49592
rect 30800 49580 30806 49632
rect 33689 49623 33747 49629
rect 33689 49589 33701 49623
rect 33735 49620 33747 49623
rect 33778 49620 33784 49632
rect 33735 49592 33784 49620
rect 33735 49589 33747 49592
rect 33689 49583 33747 49589
rect 33778 49580 33784 49592
rect 33836 49580 33842 49632
rect 35526 49580 35532 49632
rect 35584 49620 35590 49632
rect 35621 49623 35679 49629
rect 35621 49620 35633 49623
rect 35584 49592 35633 49620
rect 35584 49580 35590 49592
rect 35621 49589 35633 49592
rect 35667 49589 35679 49623
rect 35621 49583 35679 49589
rect 35894 49580 35900 49632
rect 35952 49620 35958 49632
rect 36170 49620 36176 49632
rect 35952 49592 36176 49620
rect 35952 49580 35958 49592
rect 36170 49580 36176 49592
rect 36228 49580 36234 49632
rect 1104 49530 54372 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 54372 49530
rect 1104 49456 54372 49478
rect 22281 49419 22339 49425
rect 22281 49385 22293 49419
rect 22327 49416 22339 49419
rect 25406 49416 25412 49428
rect 22327 49388 25412 49416
rect 22327 49385 22339 49388
rect 22281 49379 22339 49385
rect 25406 49376 25412 49388
rect 25464 49376 25470 49428
rect 29549 49419 29607 49425
rect 29549 49385 29561 49419
rect 29595 49416 29607 49419
rect 29730 49416 29736 49428
rect 29595 49388 29736 49416
rect 29595 49385 29607 49388
rect 29549 49379 29607 49385
rect 29730 49376 29736 49388
rect 29788 49376 29794 49428
rect 32582 49376 32588 49428
rect 32640 49416 32646 49428
rect 32677 49419 32735 49425
rect 32677 49416 32689 49419
rect 32640 49388 32689 49416
rect 32640 49376 32646 49388
rect 32677 49385 32689 49388
rect 32723 49385 32735 49419
rect 32677 49379 32735 49385
rect 36817 49419 36875 49425
rect 36817 49385 36829 49419
rect 36863 49416 36875 49419
rect 37182 49416 37188 49428
rect 36863 49388 37188 49416
rect 36863 49385 36875 49388
rect 36817 49379 36875 49385
rect 23845 49351 23903 49357
rect 23845 49317 23857 49351
rect 23891 49348 23903 49351
rect 24854 49348 24860 49360
rect 23891 49320 24860 49348
rect 23891 49317 23903 49320
rect 23845 49311 23903 49317
rect 24854 49308 24860 49320
rect 24912 49308 24918 49360
rect 29914 49308 29920 49360
rect 29972 49308 29978 49360
rect 31938 49348 31944 49360
rect 31726 49320 31944 49348
rect 23569 49283 23627 49289
rect 23569 49249 23581 49283
rect 23615 49280 23627 49283
rect 23658 49280 23664 49292
rect 23615 49252 23664 49280
rect 23615 49249 23627 49252
rect 23569 49243 23627 49249
rect 23658 49240 23664 49252
rect 23716 49240 23722 49292
rect 23934 49240 23940 49292
rect 23992 49280 23998 49292
rect 29932 49280 29960 49308
rect 30009 49283 30067 49289
rect 30009 49280 30021 49283
rect 23992 49252 26188 49280
rect 29932 49252 30021 49280
rect 23992 49240 23998 49252
rect 23474 49212 23480 49224
rect 23435 49184 23480 49212
rect 23474 49172 23480 49184
rect 23532 49172 23538 49224
rect 24394 49212 24400 49224
rect 24355 49184 24400 49212
rect 24394 49172 24400 49184
rect 24452 49172 24458 49224
rect 24486 49172 24492 49224
rect 24544 49212 24550 49224
rect 24673 49215 24731 49221
rect 24544 49184 24589 49212
rect 24544 49172 24550 49184
rect 24673 49181 24685 49215
rect 24719 49181 24731 49215
rect 25498 49212 25504 49224
rect 25459 49184 25504 49212
rect 24673 49175 24731 49181
rect 23750 49104 23756 49156
rect 23808 49144 23814 49156
rect 24688 49144 24716 49175
rect 25498 49172 25504 49184
rect 25556 49172 25562 49224
rect 26160 49221 26188 49252
rect 30009 49249 30021 49252
rect 30055 49249 30067 49283
rect 31726 49280 31754 49320
rect 31938 49308 31944 49320
rect 31996 49348 32002 49360
rect 33042 49348 33048 49360
rect 31996 49320 33048 49348
rect 31996 49308 32002 49320
rect 33042 49308 33048 49320
rect 33100 49308 33106 49360
rect 32490 49280 32496 49292
rect 30009 49243 30067 49249
rect 31312 49252 31754 49280
rect 32451 49252 32496 49280
rect 25961 49215 26019 49221
rect 25961 49181 25973 49215
rect 26007 49181 26019 49215
rect 25961 49175 26019 49181
rect 26145 49215 26203 49221
rect 26145 49181 26157 49215
rect 26191 49212 26203 49215
rect 26789 49215 26847 49221
rect 26789 49212 26801 49215
rect 26191 49184 26801 49212
rect 26191 49181 26203 49184
rect 26145 49175 26203 49181
rect 26789 49181 26801 49184
rect 26835 49181 26847 49215
rect 26789 49175 26847 49181
rect 25038 49144 25044 49156
rect 23808 49116 24716 49144
rect 24780 49116 25044 49144
rect 23808 49104 23814 49116
rect 21729 49079 21787 49085
rect 21729 49045 21741 49079
rect 21775 49076 21787 49079
rect 22002 49076 22008 49088
rect 21775 49048 22008 49076
rect 21775 49045 21787 49048
rect 21729 49039 21787 49045
rect 22002 49036 22008 49048
rect 22060 49036 22066 49088
rect 22833 49079 22891 49085
rect 22833 49045 22845 49079
rect 22879 49076 22891 49079
rect 24780 49076 24808 49116
rect 25038 49104 25044 49116
rect 25096 49104 25102 49156
rect 25976 49144 26004 49175
rect 27890 49172 27896 49224
rect 27948 49212 27954 49224
rect 27985 49215 28043 49221
rect 27985 49212 27997 49215
rect 27948 49184 27997 49212
rect 27948 49172 27954 49184
rect 27985 49181 27997 49184
rect 28031 49181 28043 49215
rect 27985 49175 28043 49181
rect 28169 49215 28227 49221
rect 28169 49181 28181 49215
rect 28215 49212 28227 49215
rect 28534 49212 28540 49224
rect 28215 49184 28540 49212
rect 28215 49181 28227 49184
rect 28169 49175 28227 49181
rect 26605 49147 26663 49153
rect 26605 49144 26617 49147
rect 25976 49116 26617 49144
rect 26605 49113 26617 49116
rect 26651 49113 26663 49147
rect 26605 49107 26663 49113
rect 22879 49048 24808 49076
rect 24857 49079 24915 49085
rect 22879 49045 22891 49048
rect 22833 49039 22891 49045
rect 24857 49045 24869 49079
rect 24903 49076 24915 49079
rect 25314 49076 25320 49088
rect 24903 49048 25320 49076
rect 24903 49045 24915 49048
rect 24857 49039 24915 49045
rect 25314 49036 25320 49048
rect 25372 49036 25378 49088
rect 25409 49079 25467 49085
rect 25409 49045 25421 49079
rect 25455 49076 25467 49079
rect 26050 49076 26056 49088
rect 25455 49048 26056 49076
rect 25455 49045 25467 49048
rect 25409 49039 25467 49045
rect 26050 49036 26056 49048
rect 26108 49036 26114 49088
rect 26145 49079 26203 49085
rect 26145 49045 26157 49079
rect 26191 49076 26203 49079
rect 26234 49076 26240 49088
rect 26191 49048 26240 49076
rect 26191 49045 26203 49048
rect 26145 49039 26203 49045
rect 26234 49036 26240 49048
rect 26292 49036 26298 49088
rect 26620 49076 26648 49107
rect 26878 49104 26884 49156
rect 26936 49144 26942 49156
rect 26973 49147 27031 49153
rect 26973 49144 26985 49147
rect 26936 49116 26985 49144
rect 26936 49104 26942 49116
rect 26973 49113 26985 49116
rect 27019 49144 27031 49147
rect 28184 49144 28212 49175
rect 28534 49172 28540 49184
rect 28592 49172 28598 49224
rect 28813 49215 28871 49221
rect 28813 49181 28825 49215
rect 28859 49181 28871 49215
rect 28813 49175 28871 49181
rect 28997 49215 29055 49221
rect 28997 49181 29009 49215
rect 29043 49212 29055 49215
rect 29546 49212 29552 49224
rect 29043 49184 29552 49212
rect 29043 49181 29055 49184
rect 28997 49175 29055 49181
rect 27019 49116 28212 49144
rect 28828 49144 28856 49175
rect 29546 49172 29552 49184
rect 29604 49172 29610 49224
rect 29730 49212 29736 49224
rect 29691 49184 29736 49212
rect 29730 49172 29736 49184
rect 29788 49172 29794 49224
rect 29822 49172 29828 49224
rect 29880 49212 29886 49224
rect 31312 49221 31340 49252
rect 32490 49240 32496 49252
rect 32548 49240 32554 49292
rect 32582 49240 32588 49292
rect 32640 49280 32646 49292
rect 33413 49283 33471 49289
rect 33413 49280 33425 49283
rect 32640 49252 33425 49280
rect 32640 49240 32646 49252
rect 33413 49249 33425 49252
rect 33459 49249 33471 49283
rect 35250 49280 35256 49292
rect 33413 49243 33471 49249
rect 33796 49252 35256 49280
rect 29917 49215 29975 49221
rect 29917 49212 29929 49215
rect 29880 49184 29929 49212
rect 29880 49172 29886 49184
rect 29917 49181 29929 49184
rect 29963 49181 29975 49215
rect 29917 49175 29975 49181
rect 30653 49215 30711 49221
rect 30653 49181 30665 49215
rect 30699 49212 30711 49215
rect 31297 49215 31355 49221
rect 31297 49212 31309 49215
rect 30699 49184 31309 49212
rect 30699 49181 30711 49184
rect 30653 49175 30711 49181
rect 31297 49181 31309 49184
rect 31343 49181 31355 49215
rect 31297 49175 31355 49181
rect 31481 49215 31539 49221
rect 31481 49181 31493 49215
rect 31527 49212 31539 49215
rect 31754 49212 31760 49224
rect 31527 49184 31760 49212
rect 31527 49181 31539 49184
rect 31481 49175 31539 49181
rect 30469 49147 30527 49153
rect 30469 49144 30481 49147
rect 28828 49116 30481 49144
rect 27019 49113 27031 49116
rect 26973 49107 27031 49113
rect 30469 49113 30481 49116
rect 30515 49113 30527 49147
rect 30469 49107 30527 49113
rect 30837 49147 30895 49153
rect 30837 49113 30849 49147
rect 30883 49144 30895 49147
rect 31496 49144 31524 49175
rect 31754 49172 31760 49184
rect 31812 49172 31818 49224
rect 32214 49172 32220 49224
rect 32272 49212 32278 49224
rect 32309 49215 32367 49221
rect 32309 49212 32321 49215
rect 32272 49184 32321 49212
rect 32272 49172 32278 49184
rect 32309 49181 32321 49184
rect 32355 49181 32367 49215
rect 32309 49175 32367 49181
rect 32398 49172 32404 49224
rect 32456 49212 32462 49224
rect 32674 49212 32680 49224
rect 32456 49184 32501 49212
rect 32635 49184 32680 49212
rect 32456 49172 32462 49184
rect 32674 49172 32680 49184
rect 32732 49172 32738 49224
rect 33226 49172 33232 49224
rect 33284 49212 33290 49224
rect 33321 49215 33379 49221
rect 33321 49212 33333 49215
rect 33284 49184 33333 49212
rect 33284 49172 33290 49184
rect 33321 49181 33333 49184
rect 33367 49181 33379 49215
rect 33502 49212 33508 49224
rect 33463 49184 33508 49212
rect 33321 49175 33379 49181
rect 33502 49172 33508 49184
rect 33560 49172 33566 49224
rect 33594 49172 33600 49224
rect 33652 49212 33658 49224
rect 33796 49221 33824 49252
rect 35250 49240 35256 49252
rect 35308 49280 35314 49292
rect 35621 49283 35679 49289
rect 35621 49280 35633 49283
rect 35308 49252 35633 49280
rect 35308 49240 35314 49252
rect 35621 49249 35633 49252
rect 35667 49249 35679 49283
rect 35621 49243 35679 49249
rect 33781 49215 33839 49221
rect 33652 49184 33697 49212
rect 33652 49172 33658 49184
rect 33781 49181 33793 49215
rect 33827 49181 33839 49215
rect 33781 49175 33839 49181
rect 34885 49215 34943 49221
rect 34885 49181 34897 49215
rect 34931 49212 34943 49215
rect 35529 49215 35587 49221
rect 35529 49212 35541 49215
rect 34931 49184 35541 49212
rect 34931 49181 34943 49184
rect 34885 49175 34943 49181
rect 35529 49181 35541 49184
rect 35575 49181 35587 49215
rect 35529 49175 35587 49181
rect 35713 49215 35771 49221
rect 35713 49181 35725 49215
rect 35759 49212 35771 49215
rect 35894 49212 35900 49224
rect 35759 49184 35900 49212
rect 35759 49181 35771 49184
rect 35713 49175 35771 49181
rect 30883 49116 31524 49144
rect 30883 49113 30895 49116
rect 30837 49107 30895 49113
rect 32490 49104 32496 49156
rect 32548 49144 32554 49156
rect 34330 49144 34336 49156
rect 32548 49116 34336 49144
rect 32548 49104 32554 49116
rect 34330 49104 34336 49116
rect 34388 49104 34394 49156
rect 35069 49147 35127 49153
rect 35069 49113 35081 49147
rect 35115 49113 35127 49147
rect 35544 49144 35572 49175
rect 35894 49172 35900 49184
rect 35952 49172 35958 49224
rect 36832 49144 36860 49379
rect 37182 49376 37188 49388
rect 37240 49416 37246 49428
rect 37277 49419 37335 49425
rect 37277 49416 37289 49419
rect 37240 49388 37289 49416
rect 37240 49376 37246 49388
rect 37277 49385 37289 49388
rect 37323 49385 37335 49419
rect 37277 49379 37335 49385
rect 35544 49116 36860 49144
rect 35069 49107 35127 49113
rect 26786 49076 26792 49088
rect 26620 49048 26792 49076
rect 26786 49036 26792 49048
rect 26844 49036 26850 49088
rect 27525 49079 27583 49085
rect 27525 49045 27537 49079
rect 27571 49076 27583 49079
rect 28074 49076 28080 49088
rect 27571 49048 28080 49076
rect 27571 49045 27583 49048
rect 27525 49039 27583 49045
rect 28074 49036 28080 49048
rect 28132 49036 28138 49088
rect 28169 49079 28227 49085
rect 28169 49045 28181 49079
rect 28215 49076 28227 49079
rect 28442 49076 28448 49088
rect 28215 49048 28448 49076
rect 28215 49045 28227 49048
rect 28169 49039 28227 49045
rect 28442 49036 28448 49048
rect 28500 49036 28506 49088
rect 28810 49076 28816 49088
rect 28771 49048 28816 49076
rect 28810 49036 28816 49048
rect 28868 49036 28874 49088
rect 29546 49036 29552 49088
rect 29604 49076 29610 49088
rect 31110 49076 31116 49088
rect 29604 49048 31116 49076
rect 29604 49036 29610 49048
rect 31110 49036 31116 49048
rect 31168 49076 31174 49088
rect 31297 49079 31355 49085
rect 31297 49076 31309 49079
rect 31168 49048 31309 49076
rect 31168 49036 31174 49048
rect 31297 49045 31309 49048
rect 31343 49045 31355 49079
rect 31297 49039 31355 49045
rect 33137 49079 33195 49085
rect 33137 49045 33149 49079
rect 33183 49076 33195 49079
rect 33410 49076 33416 49088
rect 33183 49048 33416 49076
rect 33183 49045 33195 49048
rect 33137 49039 33195 49045
rect 33410 49036 33416 49048
rect 33468 49036 33474 49088
rect 34606 49036 34612 49088
rect 34664 49076 34670 49088
rect 34701 49079 34759 49085
rect 34701 49076 34713 49079
rect 34664 49048 34713 49076
rect 34664 49036 34670 49048
rect 34701 49045 34713 49048
rect 34747 49045 34759 49079
rect 35084 49076 35112 49107
rect 35894 49076 35900 49088
rect 35084 49048 35900 49076
rect 34701 49039 34759 49045
rect 35894 49036 35900 49048
rect 35952 49076 35958 49088
rect 36173 49079 36231 49085
rect 36173 49076 36185 49079
rect 35952 49048 36185 49076
rect 35952 49036 35958 49048
rect 36173 49045 36185 49048
rect 36219 49045 36231 49079
rect 36173 49039 36231 49045
rect 1104 48986 54372 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 54372 48986
rect 1104 48912 54372 48934
rect 23477 48875 23535 48881
rect 23477 48841 23489 48875
rect 23523 48872 23535 48875
rect 23566 48872 23572 48884
rect 23523 48844 23572 48872
rect 23523 48841 23535 48844
rect 23477 48835 23535 48841
rect 23566 48832 23572 48844
rect 23624 48832 23630 48884
rect 25317 48875 25375 48881
rect 25317 48841 25329 48875
rect 25363 48872 25375 48875
rect 28258 48872 28264 48884
rect 25363 48844 28264 48872
rect 25363 48841 25375 48844
rect 25317 48835 25375 48841
rect 28258 48832 28264 48844
rect 28316 48832 28322 48884
rect 33594 48832 33600 48884
rect 33652 48872 33658 48884
rect 34333 48875 34391 48881
rect 34333 48872 34345 48875
rect 33652 48844 34345 48872
rect 33652 48832 33658 48844
rect 34333 48841 34345 48844
rect 34379 48841 34391 48875
rect 34333 48835 34391 48841
rect 24486 48764 24492 48816
rect 24544 48804 24550 48816
rect 24544 48776 25084 48804
rect 24544 48764 24550 48776
rect 21269 48739 21327 48745
rect 21269 48705 21281 48739
rect 21315 48736 21327 48739
rect 22465 48739 22523 48745
rect 22465 48736 22477 48739
rect 21315 48708 22477 48736
rect 21315 48705 21327 48708
rect 21269 48699 21327 48705
rect 22465 48705 22477 48708
rect 22511 48736 22523 48739
rect 23842 48736 23848 48748
rect 22511 48708 23848 48736
rect 22511 48705 22523 48708
rect 22465 48699 22523 48705
rect 23842 48696 23848 48708
rect 23900 48696 23906 48748
rect 24673 48739 24731 48745
rect 24673 48705 24685 48739
rect 24719 48705 24731 48739
rect 24854 48736 24860 48748
rect 24815 48708 24860 48736
rect 24673 48699 24731 48705
rect 23658 48668 23664 48680
rect 23619 48640 23664 48668
rect 23658 48628 23664 48640
rect 23716 48628 23722 48680
rect 23753 48671 23811 48677
rect 23753 48637 23765 48671
rect 23799 48637 23811 48671
rect 23753 48631 23811 48637
rect 21913 48603 21971 48609
rect 21913 48569 21925 48603
rect 21959 48600 21971 48603
rect 22922 48600 22928 48612
rect 21959 48572 22928 48600
rect 21959 48569 21971 48572
rect 21913 48563 21971 48569
rect 22922 48560 22928 48572
rect 22980 48560 22986 48612
rect 23566 48560 23572 48612
rect 23624 48600 23630 48612
rect 23768 48600 23796 48631
rect 23934 48628 23940 48680
rect 23992 48668 23998 48680
rect 23992 48640 24037 48668
rect 23992 48628 23998 48640
rect 24026 48600 24032 48612
rect 23624 48572 24032 48600
rect 23624 48560 23630 48572
rect 24026 48560 24032 48572
rect 24084 48560 24090 48612
rect 24688 48600 24716 48699
rect 24854 48696 24860 48708
rect 24912 48696 24918 48748
rect 25056 48745 25084 48776
rect 25130 48764 25136 48816
rect 25188 48804 25194 48816
rect 25188 48776 27200 48804
rect 25188 48764 25194 48776
rect 24949 48739 25007 48745
rect 24949 48705 24961 48739
rect 24995 48705 25007 48739
rect 24949 48699 25007 48705
rect 25041 48739 25099 48745
rect 25041 48705 25053 48739
rect 25087 48705 25099 48739
rect 26234 48736 26240 48748
rect 26147 48708 26240 48736
rect 25041 48699 25099 48705
rect 24964 48668 24992 48699
rect 26234 48696 26240 48708
rect 26292 48696 26298 48748
rect 26421 48739 26479 48745
rect 26421 48705 26433 48739
rect 26467 48736 26479 48739
rect 26878 48736 26884 48748
rect 26467 48708 26884 48736
rect 26467 48705 26479 48708
rect 26421 48699 26479 48705
rect 26878 48696 26884 48708
rect 26936 48696 26942 48748
rect 27172 48745 27200 48776
rect 29270 48764 29276 48816
rect 29328 48804 29334 48816
rect 33505 48807 33563 48813
rect 29328 48776 32812 48804
rect 29328 48764 29334 48776
rect 27157 48739 27215 48745
rect 27157 48705 27169 48739
rect 27203 48705 27215 48739
rect 27157 48699 27215 48705
rect 28350 48696 28356 48748
rect 28408 48736 28414 48748
rect 28537 48739 28595 48745
rect 28537 48736 28549 48739
rect 28408 48708 28549 48736
rect 28408 48696 28414 48708
rect 28537 48705 28549 48708
rect 28583 48736 28595 48739
rect 28810 48736 28816 48748
rect 28583 48708 28816 48736
rect 28583 48705 28595 48708
rect 28537 48699 28595 48705
rect 28810 48696 28816 48708
rect 28868 48696 28874 48748
rect 29546 48696 29552 48748
rect 29604 48736 29610 48748
rect 30101 48739 30159 48745
rect 30101 48736 30113 48739
rect 29604 48708 30113 48736
rect 29604 48696 29610 48708
rect 30101 48705 30113 48708
rect 30147 48705 30159 48739
rect 30101 48699 30159 48705
rect 30190 48696 30196 48748
rect 30248 48736 30254 48748
rect 30377 48739 30435 48745
rect 30248 48708 30293 48736
rect 30248 48696 30254 48708
rect 30377 48705 30389 48739
rect 30423 48705 30435 48739
rect 30834 48736 30840 48748
rect 30795 48708 30840 48736
rect 30377 48699 30435 48705
rect 25406 48668 25412 48680
rect 24964 48640 25412 48668
rect 25406 48628 25412 48640
rect 25464 48628 25470 48680
rect 26252 48668 26280 48696
rect 26602 48668 26608 48680
rect 26252 48640 26608 48668
rect 26602 48628 26608 48640
rect 26660 48628 26666 48680
rect 26786 48628 26792 48680
rect 26844 48668 26850 48680
rect 27249 48671 27307 48677
rect 27249 48668 27261 48671
rect 26844 48640 27261 48668
rect 26844 48628 26850 48640
rect 27249 48637 27261 48640
rect 27295 48668 27307 48671
rect 27706 48668 27712 48680
rect 27295 48640 27712 48668
rect 27295 48637 27307 48640
rect 27249 48631 27307 48637
rect 27706 48628 27712 48640
rect 27764 48628 27770 48680
rect 28442 48668 28448 48680
rect 28403 48640 28448 48668
rect 28442 48628 28448 48640
rect 28500 48628 28506 48680
rect 29730 48668 29736 48680
rect 28552 48640 29736 48668
rect 25038 48600 25044 48612
rect 24688 48572 25044 48600
rect 25038 48560 25044 48572
rect 25096 48600 25102 48612
rect 27522 48600 27528 48612
rect 25096 48572 26464 48600
rect 27483 48572 27528 48600
rect 25096 48560 25102 48572
rect 26326 48532 26332 48544
rect 26287 48504 26332 48532
rect 26326 48492 26332 48504
rect 26384 48492 26390 48544
rect 26436 48532 26464 48572
rect 27522 48560 27528 48572
rect 27580 48560 27586 48612
rect 28552 48532 28580 48640
rect 29730 48628 29736 48640
rect 29788 48628 29794 48680
rect 30392 48668 30420 48699
rect 30834 48696 30840 48708
rect 30892 48696 30898 48748
rect 31018 48736 31024 48748
rect 30979 48708 31024 48736
rect 31018 48696 31024 48708
rect 31076 48696 31082 48748
rect 30392 48640 30972 48668
rect 28905 48603 28963 48609
rect 28905 48569 28917 48603
rect 28951 48600 28963 48603
rect 29178 48600 29184 48612
rect 28951 48572 29184 48600
rect 28951 48569 28963 48572
rect 28905 48563 28963 48569
rect 29178 48560 29184 48572
rect 29236 48560 29242 48612
rect 30944 48544 30972 48640
rect 31294 48560 31300 48612
rect 31352 48600 31358 48612
rect 32677 48603 32735 48609
rect 32677 48600 32689 48603
rect 31352 48572 32689 48600
rect 31352 48560 31358 48572
rect 32677 48569 32689 48572
rect 32723 48569 32735 48603
rect 32677 48563 32735 48569
rect 29362 48532 29368 48544
rect 26436 48504 28580 48532
rect 29323 48504 29368 48532
rect 29362 48492 29368 48504
rect 29420 48492 29426 48544
rect 29914 48492 29920 48544
rect 29972 48532 29978 48544
rect 30101 48535 30159 48541
rect 30101 48532 30113 48535
rect 29972 48504 30113 48532
rect 29972 48492 29978 48504
rect 30101 48501 30113 48504
rect 30147 48501 30159 48535
rect 30926 48532 30932 48544
rect 30887 48504 30932 48532
rect 30101 48495 30159 48501
rect 30926 48492 30932 48504
rect 30984 48492 30990 48544
rect 31478 48532 31484 48544
rect 31439 48504 31484 48532
rect 31478 48492 31484 48504
rect 31536 48492 31542 48544
rect 32217 48535 32275 48541
rect 32217 48501 32229 48535
rect 32263 48532 32275 48535
rect 32784 48532 32812 48776
rect 33505 48773 33517 48807
rect 33551 48804 33563 48807
rect 33778 48804 33784 48816
rect 33551 48776 33784 48804
rect 33551 48773 33563 48776
rect 33505 48767 33563 48773
rect 33778 48764 33784 48776
rect 33836 48804 33842 48816
rect 34238 48804 34244 48816
rect 33836 48776 34244 48804
rect 33836 48764 33842 48776
rect 34238 48764 34244 48776
rect 34296 48804 34302 48816
rect 34425 48807 34483 48813
rect 34425 48804 34437 48807
rect 34296 48776 34437 48804
rect 34296 48764 34302 48776
rect 34425 48773 34437 48776
rect 34471 48773 34483 48807
rect 34606 48804 34612 48816
rect 34567 48776 34612 48804
rect 34425 48767 34483 48773
rect 34606 48764 34612 48776
rect 34664 48764 34670 48816
rect 33689 48739 33747 48745
rect 33689 48705 33701 48739
rect 33735 48736 33747 48739
rect 34333 48739 34391 48745
rect 34333 48736 34345 48739
rect 33735 48708 34345 48736
rect 33735 48705 33747 48708
rect 33689 48699 33747 48705
rect 34333 48705 34345 48708
rect 34379 48705 34391 48739
rect 34624 48736 34652 48764
rect 35069 48739 35127 48745
rect 35069 48736 35081 48739
rect 34624 48708 35081 48736
rect 34333 48699 34391 48705
rect 35069 48705 35081 48708
rect 35115 48705 35127 48739
rect 35250 48736 35256 48748
rect 35211 48708 35256 48736
rect 35069 48699 35127 48705
rect 34348 48668 34376 48699
rect 35250 48696 35256 48708
rect 35308 48696 35314 48748
rect 52917 48739 52975 48745
rect 52917 48705 52929 48739
rect 52963 48736 52975 48739
rect 53558 48736 53564 48748
rect 52963 48708 53564 48736
rect 52963 48705 52975 48708
rect 52917 48699 52975 48705
rect 53558 48696 53564 48708
rect 53616 48696 53622 48748
rect 35526 48668 35532 48680
rect 34348 48640 35532 48668
rect 35526 48628 35532 48640
rect 35584 48628 35590 48680
rect 33502 48560 33508 48612
rect 33560 48600 33566 48612
rect 35161 48603 35219 48609
rect 35161 48600 35173 48603
rect 33560 48572 35173 48600
rect 33560 48560 33566 48572
rect 35161 48569 35173 48572
rect 35207 48569 35219 48603
rect 35161 48563 35219 48569
rect 53098 48560 53104 48612
rect 53156 48600 53162 48612
rect 53377 48603 53435 48609
rect 53377 48600 53389 48603
rect 53156 48572 53389 48600
rect 53156 48560 53162 48572
rect 53377 48569 53389 48572
rect 53423 48569 53435 48603
rect 53377 48563 53435 48569
rect 33594 48532 33600 48544
rect 32263 48504 33600 48532
rect 32263 48501 32275 48504
rect 32217 48495 32275 48501
rect 33594 48492 33600 48504
rect 33652 48492 33658 48544
rect 33873 48535 33931 48541
rect 33873 48501 33885 48535
rect 33919 48532 33931 48535
rect 34790 48532 34796 48544
rect 33919 48504 34796 48532
rect 33919 48501 33931 48504
rect 33873 48495 33931 48501
rect 34790 48492 34796 48504
rect 34848 48492 34854 48544
rect 35526 48492 35532 48544
rect 35584 48532 35590 48544
rect 35713 48535 35771 48541
rect 35713 48532 35725 48535
rect 35584 48504 35725 48532
rect 35584 48492 35590 48504
rect 35713 48501 35725 48504
rect 35759 48532 35771 48535
rect 35802 48532 35808 48544
rect 35759 48504 35808 48532
rect 35759 48501 35771 48504
rect 35713 48495 35771 48501
rect 35802 48492 35808 48504
rect 35860 48492 35866 48544
rect 36357 48535 36415 48541
rect 36357 48501 36369 48535
rect 36403 48532 36415 48535
rect 36538 48532 36544 48544
rect 36403 48504 36544 48532
rect 36403 48501 36415 48504
rect 36357 48495 36415 48501
rect 36538 48492 36544 48504
rect 36596 48492 36602 48544
rect 1104 48442 54372 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 54372 48442
rect 1104 48368 54372 48390
rect 24854 48288 24860 48340
rect 24912 48328 24918 48340
rect 24949 48331 25007 48337
rect 24949 48328 24961 48331
rect 24912 48300 24961 48328
rect 24912 48288 24918 48300
rect 24949 48297 24961 48300
rect 24995 48297 25007 48331
rect 24949 48291 25007 48297
rect 29733 48331 29791 48337
rect 29733 48297 29745 48331
rect 29779 48328 29791 48331
rect 29822 48328 29828 48340
rect 29779 48300 29828 48328
rect 29779 48297 29791 48300
rect 29733 48291 29791 48297
rect 29822 48288 29828 48300
rect 29880 48288 29886 48340
rect 30098 48288 30104 48340
rect 30156 48328 30162 48340
rect 31478 48328 31484 48340
rect 30156 48300 31484 48328
rect 30156 48288 30162 48300
rect 31478 48288 31484 48300
rect 31536 48288 31542 48340
rect 21821 48263 21879 48269
rect 21821 48229 21833 48263
rect 21867 48260 21879 48263
rect 23845 48263 23903 48269
rect 21867 48232 22094 48260
rect 21867 48229 21879 48232
rect 21821 48223 21879 48229
rect 22066 48192 22094 48232
rect 23845 48229 23857 48263
rect 23891 48260 23903 48263
rect 24026 48260 24032 48272
rect 23891 48232 24032 48260
rect 23891 48229 23903 48232
rect 23845 48223 23903 48229
rect 24026 48220 24032 48232
rect 24084 48260 24090 48272
rect 25038 48260 25044 48272
rect 24084 48232 25044 48260
rect 24084 48220 24090 48232
rect 25038 48220 25044 48232
rect 25096 48220 25102 48272
rect 26697 48263 26755 48269
rect 26697 48229 26709 48263
rect 26743 48229 26755 48263
rect 26697 48223 26755 48229
rect 27157 48263 27215 48269
rect 27157 48229 27169 48263
rect 27203 48260 27215 48263
rect 27246 48260 27252 48272
rect 27203 48232 27252 48260
rect 27203 48229 27215 48232
rect 27157 48223 27215 48229
rect 24302 48192 24308 48204
rect 22066 48164 24308 48192
rect 24302 48152 24308 48164
rect 24360 48192 24366 48204
rect 26418 48192 26424 48204
rect 24360 48164 24808 48192
rect 26379 48164 26424 48192
rect 24360 48152 24366 48164
rect 1673 48127 1731 48133
rect 1673 48093 1685 48127
rect 1719 48093 1731 48127
rect 1673 48087 1731 48093
rect 1688 48056 1716 48087
rect 20162 48084 20168 48136
rect 20220 48124 20226 48136
rect 21177 48127 21235 48133
rect 21177 48124 21189 48127
rect 20220 48096 21189 48124
rect 20220 48084 20226 48096
rect 21177 48093 21189 48096
rect 21223 48093 21235 48127
rect 21177 48087 21235 48093
rect 22922 48084 22928 48136
rect 22980 48124 22986 48136
rect 24780 48133 24808 48164
rect 26418 48152 26424 48164
rect 26476 48152 26482 48204
rect 24489 48127 24547 48133
rect 24489 48124 24501 48127
rect 22980 48096 24501 48124
rect 22980 48084 22986 48096
rect 24489 48093 24501 48096
rect 24535 48124 24547 48127
rect 24765 48127 24823 48133
rect 24535 48096 24716 48124
rect 24535 48093 24547 48096
rect 24489 48087 24547 48093
rect 2222 48056 2228 48068
rect 1688 48028 2228 48056
rect 2222 48016 2228 48028
rect 2280 48016 2286 48068
rect 23842 48016 23848 48068
rect 23900 48056 23906 48068
rect 24581 48059 24639 48065
rect 24581 48056 24593 48059
rect 23900 48028 24593 48056
rect 23900 48016 23906 48028
rect 24581 48025 24593 48028
rect 24627 48025 24639 48059
rect 24688 48056 24716 48096
rect 24765 48093 24777 48127
rect 24811 48093 24823 48127
rect 24765 48087 24823 48093
rect 24854 48084 24860 48136
rect 24912 48124 24918 48136
rect 25409 48127 25467 48133
rect 25409 48124 25421 48127
rect 24912 48096 25421 48124
rect 24912 48084 24918 48096
rect 25409 48093 25421 48096
rect 25455 48093 25467 48127
rect 25409 48087 25467 48093
rect 25593 48127 25651 48133
rect 25593 48093 25605 48127
rect 25639 48093 25651 48127
rect 26326 48124 26332 48136
rect 26287 48096 26332 48124
rect 25593 48087 25651 48093
rect 25608 48056 25636 48087
rect 26326 48084 26332 48096
rect 26384 48084 26390 48136
rect 26712 48124 26740 48223
rect 27246 48220 27252 48232
rect 27304 48220 27310 48272
rect 28997 48263 29055 48269
rect 28997 48229 29009 48263
rect 29043 48260 29055 48263
rect 30190 48260 30196 48272
rect 29043 48232 30196 48260
rect 29043 48229 29055 48232
rect 28997 48223 29055 48229
rect 30190 48220 30196 48232
rect 30248 48260 30254 48272
rect 30248 48232 31248 48260
rect 30248 48220 30254 48232
rect 28902 48192 28908 48204
rect 27723 48164 28908 48192
rect 27295 48127 27353 48133
rect 27295 48124 27307 48127
rect 26712 48096 27307 48124
rect 27295 48093 27307 48096
rect 27341 48093 27353 48127
rect 27522 48124 27528 48136
rect 27483 48096 27528 48124
rect 27295 48087 27353 48093
rect 27522 48084 27528 48096
rect 27580 48084 27586 48136
rect 27723 48133 27751 48164
rect 28902 48152 28908 48164
rect 28960 48152 28966 48204
rect 29914 48192 29920 48204
rect 29875 48164 29920 48192
rect 29914 48152 29920 48164
rect 29972 48152 29978 48204
rect 30009 48195 30067 48201
rect 30009 48161 30021 48195
rect 30055 48192 30067 48195
rect 30745 48195 30803 48201
rect 30745 48192 30757 48195
rect 30055 48164 30757 48192
rect 30055 48161 30067 48164
rect 30009 48155 30067 48161
rect 30745 48161 30757 48164
rect 30791 48161 30803 48195
rect 30745 48155 30803 48161
rect 27708 48127 27766 48133
rect 27708 48093 27720 48127
rect 27754 48093 27766 48127
rect 27708 48087 27766 48093
rect 27801 48127 27859 48133
rect 27801 48093 27813 48127
rect 27847 48124 27859 48127
rect 28166 48124 28172 48136
rect 27847 48096 28172 48124
rect 27847 48093 27859 48096
rect 27801 48087 27859 48093
rect 28166 48084 28172 48096
rect 28224 48084 28230 48136
rect 28350 48124 28356 48136
rect 28311 48096 28356 48124
rect 28350 48084 28356 48096
rect 28408 48084 28414 48136
rect 28534 48124 28540 48136
rect 28495 48096 28540 48124
rect 28534 48084 28540 48096
rect 28592 48084 28598 48136
rect 28626 48084 28632 48136
rect 28684 48124 28690 48136
rect 29270 48124 29276 48136
rect 28684 48096 28729 48124
rect 28966 48096 29276 48124
rect 28684 48084 28690 48096
rect 27433 48059 27491 48065
rect 27433 48056 27445 48059
rect 24688 48028 27445 48056
rect 24581 48019 24639 48025
rect 27433 48025 27445 48028
rect 27479 48056 27491 48059
rect 28966 48056 28994 48096
rect 29270 48084 29276 48096
rect 29328 48124 29334 48136
rect 30101 48127 30159 48133
rect 30101 48124 30113 48127
rect 29328 48096 30113 48124
rect 29328 48084 29334 48096
rect 30101 48093 30113 48096
rect 30147 48093 30159 48127
rect 30101 48087 30159 48093
rect 30193 48127 30251 48133
rect 30193 48093 30205 48127
rect 30239 48124 30251 48127
rect 30282 48124 30288 48136
rect 30239 48096 30288 48124
rect 30239 48093 30251 48096
rect 30193 48087 30251 48093
rect 30282 48084 30288 48096
rect 30340 48084 30346 48136
rect 30926 48124 30932 48136
rect 30839 48096 30932 48124
rect 30926 48084 30932 48096
rect 30984 48084 30990 48136
rect 31110 48124 31116 48136
rect 31071 48096 31116 48124
rect 31110 48084 31116 48096
rect 31168 48084 31174 48136
rect 31220 48133 31248 48232
rect 32214 48220 32220 48272
rect 32272 48260 32278 48272
rect 36081 48263 36139 48269
rect 36081 48260 36093 48263
rect 32272 48232 36093 48260
rect 32272 48220 32278 48232
rect 36081 48229 36093 48232
rect 36127 48229 36139 48263
rect 36081 48223 36139 48229
rect 32398 48192 32404 48204
rect 32232 48164 32404 48192
rect 32232 48133 32260 48164
rect 32398 48152 32404 48164
rect 32456 48152 32462 48204
rect 32677 48195 32735 48201
rect 32677 48161 32689 48195
rect 32723 48192 32735 48195
rect 33597 48195 33655 48201
rect 33597 48192 33609 48195
rect 32723 48164 33609 48192
rect 32723 48161 32735 48164
rect 32677 48155 32735 48161
rect 33597 48161 33609 48164
rect 33643 48192 33655 48195
rect 34793 48195 34851 48201
rect 34793 48192 34805 48195
rect 33643 48164 34805 48192
rect 33643 48161 33655 48164
rect 33597 48155 33655 48161
rect 34793 48161 34805 48164
rect 34839 48161 34851 48195
rect 34793 48155 34851 48161
rect 34977 48195 35035 48201
rect 34977 48161 34989 48195
rect 35023 48192 35035 48195
rect 35342 48192 35348 48204
rect 35023 48164 35348 48192
rect 35023 48161 35035 48164
rect 34977 48155 35035 48161
rect 35342 48152 35348 48164
rect 35400 48192 35406 48204
rect 35529 48195 35587 48201
rect 35529 48192 35541 48195
rect 35400 48164 35541 48192
rect 35400 48152 35406 48164
rect 35529 48161 35541 48164
rect 35575 48161 35587 48195
rect 35529 48155 35587 48161
rect 35802 48152 35808 48204
rect 35860 48192 35866 48204
rect 37277 48195 37335 48201
rect 37277 48192 37289 48195
rect 35860 48164 37289 48192
rect 35860 48152 35866 48164
rect 37277 48161 37289 48164
rect 37323 48161 37335 48195
rect 37277 48155 37335 48161
rect 31205 48127 31263 48133
rect 31205 48093 31217 48127
rect 31251 48124 31263 48127
rect 32217 48127 32275 48133
rect 32217 48124 32229 48127
rect 31251 48096 32229 48124
rect 31251 48093 31263 48096
rect 31205 48087 31263 48093
rect 32217 48093 32229 48096
rect 32263 48093 32275 48127
rect 32217 48087 32275 48093
rect 32309 48127 32367 48133
rect 32309 48093 32321 48127
rect 32355 48093 32367 48127
rect 32309 48087 32367 48093
rect 32493 48127 32551 48133
rect 32493 48093 32505 48127
rect 32539 48124 32551 48127
rect 32582 48124 32588 48136
rect 32539 48096 32588 48124
rect 32539 48093 32551 48096
rect 32493 48087 32551 48093
rect 27479 48028 28994 48056
rect 30944 48056 30972 48084
rect 32324 48056 32352 48087
rect 32582 48084 32588 48096
rect 32640 48084 32646 48136
rect 33226 48084 33232 48136
rect 33284 48124 33290 48136
rect 33505 48127 33563 48133
rect 33505 48124 33517 48127
rect 33284 48096 33517 48124
rect 33284 48084 33290 48096
rect 33505 48093 33517 48096
rect 33551 48124 33563 48127
rect 34422 48124 34428 48136
rect 33551 48096 34428 48124
rect 33551 48093 33563 48096
rect 33505 48087 33563 48093
rect 34422 48084 34428 48096
rect 34480 48124 34486 48136
rect 34701 48127 34759 48133
rect 34701 48124 34713 48127
rect 34480 48096 34713 48124
rect 34480 48084 34486 48096
rect 34701 48093 34713 48096
rect 34747 48093 34759 48127
rect 34701 48087 34759 48093
rect 35437 48127 35495 48133
rect 35437 48093 35449 48127
rect 35483 48124 35495 48127
rect 35621 48127 35679 48133
rect 35483 48096 35572 48124
rect 35483 48093 35495 48096
rect 35437 48087 35495 48093
rect 35544 48068 35572 48096
rect 35621 48093 35633 48127
rect 35667 48124 35679 48127
rect 36538 48124 36544 48136
rect 35667 48096 36544 48124
rect 35667 48093 35679 48096
rect 35621 48087 35679 48093
rect 33042 48056 33048 48068
rect 30944 48028 33048 48056
rect 27479 48025 27491 48028
rect 27433 48019 27491 48025
rect 33042 48016 33048 48028
rect 33100 48016 33106 48068
rect 34238 48016 34244 48068
rect 34296 48056 34302 48068
rect 34296 48028 35112 48056
rect 34296 48016 34302 48028
rect 1486 47988 1492 48000
rect 1447 47960 1492 47988
rect 1486 47948 1492 47960
rect 1544 47948 1550 48000
rect 20714 47988 20720 48000
rect 20675 47960 20720 47988
rect 20714 47948 20720 47960
rect 20772 47948 20778 48000
rect 22002 47948 22008 48000
rect 22060 47988 22066 48000
rect 22281 47991 22339 47997
rect 22281 47988 22293 47991
rect 22060 47960 22293 47988
rect 22060 47948 22066 47960
rect 22281 47957 22293 47960
rect 22327 47957 22339 47991
rect 22281 47951 22339 47957
rect 22925 47991 22983 47997
rect 22925 47957 22937 47991
rect 22971 47988 22983 47991
rect 23106 47988 23112 48000
rect 22971 47960 23112 47988
rect 22971 47957 22983 47960
rect 22925 47951 22983 47957
rect 23106 47948 23112 47960
rect 23164 47948 23170 48000
rect 25593 47991 25651 47997
rect 25593 47957 25605 47991
rect 25639 47988 25651 47991
rect 26234 47988 26240 48000
rect 25639 47960 26240 47988
rect 25639 47957 25651 47960
rect 25593 47951 25651 47957
rect 26234 47948 26240 47960
rect 26292 47948 26298 48000
rect 29914 47948 29920 48000
rect 29972 47988 29978 48000
rect 31665 47991 31723 47997
rect 31665 47988 31677 47991
rect 29972 47960 31677 47988
rect 29972 47948 29978 47960
rect 31665 47957 31677 47960
rect 31711 47988 31723 47991
rect 31754 47988 31760 48000
rect 31711 47960 31760 47988
rect 31711 47957 31723 47960
rect 31665 47951 31723 47957
rect 31754 47948 31760 47960
rect 31812 47948 31818 48000
rect 33134 47988 33140 48000
rect 33095 47960 33140 47988
rect 33134 47948 33140 47960
rect 33192 47948 33198 48000
rect 34606 47948 34612 48000
rect 34664 47988 34670 48000
rect 34977 47991 35035 47997
rect 34977 47988 34989 47991
rect 34664 47960 34989 47988
rect 34664 47948 34670 47960
rect 34977 47957 34989 47960
rect 35023 47957 35035 47991
rect 35084 47988 35112 48028
rect 35526 48016 35532 48068
rect 35584 48016 35590 48068
rect 35636 47988 35664 48087
rect 36538 48084 36544 48096
rect 36596 48084 36602 48136
rect 35084 47960 35664 47988
rect 34977 47951 35035 47957
rect 36538 47948 36544 48000
rect 36596 47988 36602 48000
rect 36633 47991 36691 47997
rect 36633 47988 36645 47991
rect 36596 47960 36645 47988
rect 36596 47948 36602 47960
rect 36633 47957 36645 47960
rect 36679 47957 36691 47991
rect 36633 47951 36691 47957
rect 1104 47898 54372 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 54372 47898
rect 1104 47824 54372 47846
rect 23477 47787 23535 47793
rect 23477 47753 23489 47787
rect 23523 47784 23535 47787
rect 23934 47784 23940 47796
rect 23523 47756 23940 47784
rect 23523 47753 23535 47756
rect 23477 47747 23535 47753
rect 23934 47744 23940 47756
rect 23992 47744 23998 47796
rect 24026 47744 24032 47796
rect 24084 47784 24090 47796
rect 24581 47787 24639 47793
rect 24084 47756 24129 47784
rect 24084 47744 24090 47756
rect 24581 47753 24593 47787
rect 24627 47784 24639 47787
rect 25682 47784 25688 47796
rect 24627 47756 25688 47784
rect 24627 47753 24639 47756
rect 24581 47747 24639 47753
rect 25682 47744 25688 47756
rect 25740 47784 25746 47796
rect 26418 47784 26424 47796
rect 25740 47756 26188 47784
rect 26379 47756 26424 47784
rect 25740 47744 25746 47756
rect 21542 47676 21548 47728
rect 21600 47716 21606 47728
rect 22002 47716 22008 47728
rect 21600 47688 22008 47716
rect 21600 47676 21606 47688
rect 22002 47676 22008 47688
rect 22060 47716 22066 47728
rect 25317 47719 25375 47725
rect 25317 47716 25329 47719
rect 22060 47688 25329 47716
rect 22060 47676 22066 47688
rect 20162 47608 20168 47660
rect 20220 47648 20226 47660
rect 22278 47648 22284 47660
rect 20220 47620 22284 47648
rect 20220 47608 20226 47620
rect 22278 47608 22284 47620
rect 22336 47608 22342 47660
rect 24504 47657 24532 47688
rect 25317 47685 25329 47688
rect 25363 47685 25375 47719
rect 25498 47716 25504 47728
rect 25459 47688 25504 47716
rect 25317 47679 25375 47685
rect 25498 47676 25504 47688
rect 25556 47676 25562 47728
rect 26160 47716 26188 47756
rect 26418 47744 26424 47756
rect 26476 47744 26482 47796
rect 28994 47784 29000 47796
rect 28955 47756 29000 47784
rect 28994 47744 29000 47756
rect 29052 47744 29058 47796
rect 30561 47787 30619 47793
rect 30561 47753 30573 47787
rect 30607 47784 30619 47787
rect 30834 47784 30840 47796
rect 30607 47756 30840 47784
rect 30607 47753 30619 47756
rect 30561 47747 30619 47753
rect 30834 47744 30840 47756
rect 30892 47744 30898 47796
rect 31205 47787 31263 47793
rect 31205 47753 31217 47787
rect 31251 47784 31263 47787
rect 32582 47784 32588 47796
rect 31251 47756 32588 47784
rect 31251 47753 31263 47756
rect 31205 47747 31263 47753
rect 32582 47744 32588 47756
rect 32640 47744 32646 47796
rect 34422 47744 34428 47796
rect 34480 47784 34486 47796
rect 35253 47787 35311 47793
rect 35253 47784 35265 47787
rect 34480 47756 35265 47784
rect 34480 47744 34486 47756
rect 35253 47753 35265 47756
rect 35299 47753 35311 47787
rect 35253 47747 35311 47753
rect 27709 47719 27767 47725
rect 26160 47688 27568 47716
rect 23293 47651 23351 47657
rect 23293 47648 23305 47651
rect 22388 47620 23305 47648
rect 20714 47540 20720 47592
rect 20772 47580 20778 47592
rect 22388 47589 22416 47620
rect 23293 47617 23305 47620
rect 23339 47617 23351 47651
rect 23293 47611 23351 47617
rect 24489 47651 24547 47657
rect 24489 47617 24501 47651
rect 24535 47617 24547 47651
rect 24489 47611 24547 47617
rect 24673 47651 24731 47657
rect 24673 47617 24685 47651
rect 24719 47648 24731 47651
rect 25130 47648 25136 47660
rect 24719 47620 25136 47648
rect 24719 47617 24731 47620
rect 24673 47611 24731 47617
rect 25130 47608 25136 47620
rect 25188 47608 25194 47660
rect 26050 47648 26056 47660
rect 26011 47620 26056 47648
rect 26050 47608 26056 47620
rect 26108 47608 26114 47660
rect 26160 47648 26188 47688
rect 26237 47651 26295 47657
rect 26237 47648 26249 47651
rect 26160 47620 26249 47648
rect 26237 47617 26249 47620
rect 26283 47617 26295 47651
rect 26973 47651 27031 47657
rect 26973 47648 26985 47651
rect 26237 47611 26295 47617
rect 26436 47620 26985 47648
rect 22373 47583 22431 47589
rect 22373 47580 22385 47583
rect 20772 47552 22385 47580
rect 20772 47540 20778 47552
rect 22373 47549 22385 47552
rect 22419 47549 22431 47583
rect 23109 47583 23167 47589
rect 23109 47580 23121 47583
rect 22373 47543 22431 47549
rect 22480 47552 23121 47580
rect 22278 47472 22284 47524
rect 22336 47512 22342 47524
rect 22480 47512 22508 47552
rect 23109 47549 23121 47552
rect 23155 47580 23167 47583
rect 23382 47580 23388 47592
rect 23155 47552 23388 47580
rect 23155 47549 23167 47552
rect 23109 47543 23167 47549
rect 23382 47540 23388 47552
rect 23440 47540 23446 47592
rect 25314 47540 25320 47592
rect 25372 47580 25378 47592
rect 25866 47580 25872 47592
rect 25372 47552 25872 47580
rect 25372 47540 25378 47552
rect 25866 47540 25872 47552
rect 25924 47580 25930 47592
rect 25961 47583 26019 47589
rect 25961 47580 25973 47583
rect 25924 47552 25973 47580
rect 25924 47540 25930 47552
rect 25961 47549 25973 47552
rect 26007 47549 26019 47583
rect 25961 47543 26019 47549
rect 22336 47484 22508 47512
rect 22649 47515 22707 47521
rect 22336 47472 22342 47484
rect 22649 47481 22661 47515
rect 22695 47512 22707 47515
rect 23658 47512 23664 47524
rect 22695 47484 23664 47512
rect 22695 47481 22707 47484
rect 22649 47475 22707 47481
rect 23658 47472 23664 47484
rect 23716 47472 23722 47524
rect 25976 47512 26004 47543
rect 26436 47512 26464 47620
rect 26973 47617 26985 47620
rect 27019 47648 27031 47651
rect 27154 47648 27160 47660
rect 27019 47620 27160 47648
rect 27019 47617 27031 47620
rect 26973 47611 27031 47617
rect 27154 47608 27160 47620
rect 27212 47608 27218 47660
rect 27249 47651 27307 47657
rect 27249 47617 27261 47651
rect 27295 47617 27307 47651
rect 27249 47611 27307 47617
rect 27264 47580 27292 47611
rect 27430 47608 27436 47660
rect 27488 47648 27494 47660
rect 27540 47657 27568 47688
rect 27709 47685 27721 47719
rect 27755 47716 27767 47719
rect 27890 47716 27896 47728
rect 27755 47688 27896 47716
rect 27755 47685 27767 47688
rect 27709 47679 27767 47685
rect 27890 47676 27896 47688
rect 27948 47716 27954 47728
rect 28626 47716 28632 47728
rect 27948 47688 28632 47716
rect 27948 47676 27954 47688
rect 28626 47676 28632 47688
rect 28684 47676 28690 47728
rect 29270 47716 29276 47728
rect 29231 47688 29276 47716
rect 29270 47676 29276 47688
rect 29328 47676 29334 47728
rect 31294 47676 31300 47728
rect 31352 47716 31358 47728
rect 33778 47716 33784 47728
rect 31352 47688 33784 47716
rect 31352 47676 31358 47688
rect 29178 47657 29184 47660
rect 27525 47651 27583 47657
rect 27525 47648 27537 47651
rect 27488 47620 27537 47648
rect 27488 47608 27494 47620
rect 27525 47617 27537 47620
rect 27571 47617 27583 47651
rect 29176 47648 29184 47657
rect 29139 47620 29184 47648
rect 27525 47611 27583 47617
rect 29176 47611 29184 47620
rect 29178 47608 29184 47611
rect 29236 47608 29242 47660
rect 29362 47608 29368 47660
rect 29420 47648 29426 47660
rect 29548 47651 29606 47657
rect 29420 47620 29465 47648
rect 29420 47608 29426 47620
rect 29548 47617 29560 47651
rect 29594 47617 29606 47651
rect 29548 47611 29606 47617
rect 29641 47651 29699 47657
rect 29641 47617 29653 47651
rect 29687 47648 29699 47651
rect 30558 47648 30564 47660
rect 29687 47620 30564 47648
rect 29687 47617 29699 47620
rect 29641 47611 29699 47617
rect 25976 47484 26464 47512
rect 26528 47552 27292 47580
rect 20162 47444 20168 47456
rect 20123 47416 20168 47444
rect 20162 47404 20168 47416
rect 20220 47404 20226 47456
rect 20714 47444 20720 47456
rect 20675 47416 20720 47444
rect 20714 47404 20720 47416
rect 20772 47404 20778 47456
rect 21269 47447 21327 47453
rect 21269 47413 21281 47447
rect 21315 47444 21327 47447
rect 21542 47444 21548 47456
rect 21315 47416 21548 47444
rect 21315 47413 21327 47416
rect 21269 47407 21327 47413
rect 21542 47404 21548 47416
rect 21600 47404 21606 47456
rect 26050 47404 26056 47456
rect 26108 47444 26114 47456
rect 26528 47444 26556 47552
rect 28902 47540 28908 47592
rect 28960 47580 28966 47592
rect 29563 47580 29591 47611
rect 30558 47608 30564 47620
rect 30616 47608 30622 47660
rect 31018 47648 31024 47660
rect 30979 47620 31024 47648
rect 31018 47608 31024 47620
rect 31076 47648 31082 47660
rect 31076 47620 31754 47648
rect 31076 47608 31082 47620
rect 28960 47552 29591 47580
rect 30929 47583 30987 47589
rect 28960 47540 28966 47552
rect 30929 47549 30941 47583
rect 30975 47580 30987 47583
rect 31110 47580 31116 47592
rect 30975 47552 31116 47580
rect 30975 47549 30987 47552
rect 30929 47543 30987 47549
rect 31110 47540 31116 47552
rect 31168 47540 31174 47592
rect 31726 47580 31754 47620
rect 32030 47608 32036 47660
rect 32088 47654 32094 47660
rect 32324 47657 32352 47688
rect 33778 47676 33784 47688
rect 33836 47676 33842 47728
rect 32125 47654 32183 47657
rect 32088 47651 32183 47654
rect 32088 47626 32137 47651
rect 32088 47608 32094 47626
rect 32125 47617 32137 47626
rect 32171 47617 32183 47651
rect 32125 47611 32183 47617
rect 32309 47651 32367 47657
rect 32309 47617 32321 47651
rect 32355 47617 32367 47651
rect 32309 47611 32367 47617
rect 32398 47608 32404 47660
rect 32456 47648 32462 47660
rect 32953 47651 33011 47657
rect 32953 47648 32965 47651
rect 32456 47620 32965 47648
rect 32456 47608 32462 47620
rect 32953 47617 32965 47620
rect 32999 47617 33011 47651
rect 32953 47611 33011 47617
rect 33042 47608 33048 47660
rect 33100 47648 33106 47660
rect 33137 47651 33195 47657
rect 33137 47648 33149 47651
rect 33100 47620 33149 47648
rect 33100 47608 33106 47620
rect 33137 47617 33149 47620
rect 33183 47617 33195 47651
rect 33137 47611 33195 47617
rect 33226 47608 33232 47660
rect 33284 47648 33290 47660
rect 33410 47648 33416 47660
rect 33284 47620 33329 47648
rect 33371 47620 33416 47648
rect 33284 47608 33290 47620
rect 33410 47608 33416 47620
rect 33468 47608 33474 47660
rect 34517 47651 34575 47657
rect 34517 47648 34529 47651
rect 33520 47620 34529 47648
rect 33520 47592 33548 47620
rect 34517 47617 34529 47620
rect 34563 47617 34575 47651
rect 34517 47611 34575 47617
rect 34790 47608 34796 47660
rect 34848 47648 34854 47660
rect 35161 47651 35219 47657
rect 35161 47648 35173 47651
rect 34848 47620 35173 47648
rect 34848 47608 34854 47620
rect 35161 47617 35173 47620
rect 35207 47617 35219 47651
rect 35342 47648 35348 47660
rect 35303 47620 35348 47648
rect 35161 47611 35219 47617
rect 35342 47608 35348 47620
rect 35400 47608 35406 47660
rect 32217 47583 32275 47589
rect 32217 47580 32229 47583
rect 31726 47552 32229 47580
rect 32217 47549 32229 47552
rect 32263 47549 32275 47583
rect 32217 47543 32275 47549
rect 33321 47583 33379 47589
rect 33321 47549 33333 47583
rect 33367 47580 33379 47583
rect 33502 47580 33508 47592
rect 33367 47552 33508 47580
rect 33367 47549 33379 47552
rect 33321 47543 33379 47549
rect 33502 47540 33508 47552
rect 33560 47540 33566 47592
rect 34606 47580 34612 47592
rect 34567 47552 34612 47580
rect 34606 47540 34612 47552
rect 34664 47540 34670 47592
rect 26602 47472 26608 47524
rect 26660 47512 26666 47524
rect 27801 47515 27859 47521
rect 27801 47512 27813 47515
rect 26660 47484 27813 47512
rect 26660 47472 26666 47484
rect 27801 47481 27813 47484
rect 27847 47481 27859 47515
rect 27801 47475 27859 47481
rect 33226 47472 33232 47524
rect 33284 47512 33290 47524
rect 34149 47515 34207 47521
rect 34149 47512 34161 47515
rect 33284 47484 34161 47512
rect 33284 47472 33290 47484
rect 34149 47481 34161 47484
rect 34195 47481 34207 47515
rect 34149 47475 34207 47481
rect 35342 47472 35348 47524
rect 35400 47512 35406 47524
rect 36357 47515 36415 47521
rect 36357 47512 36369 47515
rect 35400 47484 36369 47512
rect 35400 47472 35406 47484
rect 36357 47481 36369 47484
rect 36403 47481 36415 47515
rect 36357 47475 36415 47481
rect 28534 47444 28540 47456
rect 26108 47416 26556 47444
rect 28495 47416 28540 47444
rect 26108 47404 26114 47416
rect 28534 47404 28540 47416
rect 28592 47404 28598 47456
rect 33686 47444 33692 47456
rect 33647 47416 33692 47444
rect 33686 47404 33692 47416
rect 33744 47404 33750 47456
rect 35802 47444 35808 47456
rect 35763 47416 35808 47444
rect 35802 47404 35808 47416
rect 35860 47404 35866 47456
rect 37369 47447 37427 47453
rect 37369 47413 37381 47447
rect 37415 47444 37427 47447
rect 37458 47444 37464 47456
rect 37415 47416 37464 47444
rect 37415 47413 37427 47416
rect 37369 47407 37427 47413
rect 37458 47404 37464 47416
rect 37516 47404 37522 47456
rect 1104 47354 54372 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 54372 47354
rect 1104 47280 54372 47302
rect 24670 47200 24676 47252
rect 24728 47240 24734 47252
rect 26418 47240 26424 47252
rect 24728 47212 26424 47240
rect 24728 47200 24734 47212
rect 26418 47200 26424 47212
rect 26476 47200 26482 47252
rect 26697 47243 26755 47249
rect 26697 47209 26709 47243
rect 26743 47240 26755 47243
rect 26970 47240 26976 47252
rect 26743 47212 26976 47240
rect 26743 47209 26755 47212
rect 26697 47203 26755 47209
rect 26970 47200 26976 47212
rect 27028 47200 27034 47252
rect 28629 47243 28687 47249
rect 27080 47212 27292 47240
rect 23569 47175 23627 47181
rect 23569 47141 23581 47175
rect 23615 47172 23627 47175
rect 24394 47172 24400 47184
rect 23615 47144 24400 47172
rect 23615 47141 23627 47144
rect 23569 47135 23627 47141
rect 24394 47132 24400 47144
rect 24452 47132 24458 47184
rect 25222 47132 25228 47184
rect 25280 47132 25286 47184
rect 25498 47132 25504 47184
rect 25556 47172 25562 47184
rect 27080 47172 27108 47212
rect 25556 47144 27108 47172
rect 27157 47175 27215 47181
rect 25556 47132 25562 47144
rect 27157 47141 27169 47175
rect 27203 47141 27215 47175
rect 27157 47135 27215 47141
rect 23293 47107 23351 47113
rect 23293 47073 23305 47107
rect 23339 47104 23351 47107
rect 23382 47104 23388 47116
rect 23339 47076 23388 47104
rect 23339 47073 23351 47076
rect 23293 47067 23351 47073
rect 23382 47064 23388 47076
rect 23440 47064 23446 47116
rect 24489 47107 24547 47113
rect 24489 47073 24501 47107
rect 24535 47104 24547 47107
rect 24578 47104 24584 47116
rect 24535 47076 24584 47104
rect 24535 47073 24547 47076
rect 24489 47067 24547 47073
rect 24578 47064 24584 47076
rect 24636 47064 24642 47116
rect 20162 46996 20168 47048
rect 20220 47036 20226 47048
rect 20257 47039 20315 47045
rect 20257 47036 20269 47039
rect 20220 47008 20269 47036
rect 20220 46996 20226 47008
rect 20257 47005 20269 47008
rect 20303 47036 20315 47039
rect 23201 47039 23259 47045
rect 20303 47008 20668 47036
rect 20303 47005 20315 47008
rect 20257 46999 20315 47005
rect 20640 46980 20668 47008
rect 23201 47005 23213 47039
rect 23247 47036 23259 47039
rect 23566 47036 23572 47048
rect 23247 47008 23572 47036
rect 23247 47005 23259 47008
rect 23201 46999 23259 47005
rect 23566 46996 23572 47008
rect 23624 47036 23630 47048
rect 24670 47036 24676 47048
rect 23624 47008 24676 47036
rect 23624 46996 23630 47008
rect 24670 46996 24676 47008
rect 24728 46996 24734 47048
rect 24946 47036 24952 47048
rect 24907 47008 24952 47036
rect 24946 46996 24952 47008
rect 25004 46996 25010 47048
rect 25038 46996 25044 47048
rect 25096 47036 25102 47048
rect 25240 47045 25268 47132
rect 27172 47104 27200 47135
rect 25332 47076 27200 47104
rect 25332 47045 25360 47076
rect 25133 47039 25191 47045
rect 25133 47036 25145 47039
rect 25096 47008 25145 47036
rect 25096 46996 25102 47008
rect 25133 47005 25145 47008
rect 25179 47005 25191 47039
rect 25133 46999 25191 47005
rect 25225 47039 25283 47045
rect 25225 47005 25237 47039
rect 25271 47005 25283 47039
rect 25225 46999 25283 47005
rect 25317 47039 25375 47045
rect 25317 47005 25329 47039
rect 25363 47005 25375 47039
rect 25774 47036 25780 47048
rect 25317 46999 25375 47005
rect 25516 47008 25780 47036
rect 20622 46928 20628 46980
rect 20680 46968 20686 46980
rect 20717 46971 20775 46977
rect 20717 46968 20729 46971
rect 20680 46940 20729 46968
rect 20680 46928 20686 46940
rect 20717 46937 20729 46940
rect 20763 46937 20775 46971
rect 20717 46931 20775 46937
rect 21361 46971 21419 46977
rect 21361 46937 21373 46971
rect 21407 46968 21419 46971
rect 22462 46968 22468 46980
rect 21407 46940 22468 46968
rect 21407 46937 21419 46940
rect 21361 46931 21419 46937
rect 22462 46928 22468 46940
rect 22520 46928 22526 46980
rect 24964 46968 24992 46996
rect 25516 46968 25544 47008
rect 25774 46996 25780 47008
rect 25832 47036 25838 47048
rect 26053 47039 26111 47045
rect 26053 47036 26065 47039
rect 25832 47008 26065 47036
rect 25832 46996 25838 47008
rect 26053 47005 26065 47008
rect 26099 47005 26111 47039
rect 26234 47036 26240 47048
rect 26195 47008 26240 47036
rect 26053 46999 26111 47005
rect 26234 46996 26240 47008
rect 26292 46996 26298 47048
rect 26329 47039 26387 47045
rect 26329 47005 26341 47039
rect 26375 47005 26387 47039
rect 26329 46999 26387 47005
rect 24964 46940 25544 46968
rect 25593 46971 25651 46977
rect 25593 46937 25605 46971
rect 25639 46968 25651 46971
rect 25639 46940 26280 46968
rect 25639 46937 25651 46940
rect 25593 46931 25651 46937
rect 26252 46912 26280 46940
rect 19334 46860 19340 46912
rect 19392 46900 19398 46912
rect 19613 46903 19671 46909
rect 19613 46900 19625 46903
rect 19392 46872 19625 46900
rect 19392 46860 19398 46872
rect 19613 46869 19625 46872
rect 19659 46869 19671 46903
rect 21818 46900 21824 46912
rect 21779 46872 21824 46900
rect 19613 46863 19671 46869
rect 21818 46860 21824 46872
rect 21876 46860 21882 46912
rect 22370 46900 22376 46912
rect 22331 46872 22376 46900
rect 22370 46860 22376 46872
rect 22428 46860 22434 46912
rect 26234 46860 26240 46912
rect 26292 46860 26298 46912
rect 26344 46900 26372 46999
rect 26418 46996 26424 47048
rect 26476 47036 26482 47048
rect 27154 47036 27160 47048
rect 26476 47008 26521 47036
rect 27115 47008 27160 47036
rect 26476 46996 26482 47008
rect 27154 46996 27160 47008
rect 27212 46996 27218 47048
rect 27264 46968 27292 47212
rect 28629 47209 28641 47243
rect 28675 47240 28687 47243
rect 29362 47240 29368 47252
rect 28675 47212 29368 47240
rect 28675 47209 28687 47212
rect 28629 47203 28687 47209
rect 29362 47200 29368 47212
rect 29420 47200 29426 47252
rect 30282 47240 30288 47252
rect 30243 47212 30288 47240
rect 30282 47200 30288 47212
rect 30340 47200 30346 47252
rect 30745 47243 30803 47249
rect 30745 47209 30757 47243
rect 30791 47240 30803 47243
rect 30834 47240 30840 47252
rect 30791 47212 30840 47240
rect 30791 47209 30803 47212
rect 30745 47203 30803 47209
rect 30834 47200 30840 47212
rect 30892 47200 30898 47252
rect 32674 47200 32680 47252
rect 32732 47240 32738 47252
rect 32953 47243 33011 47249
rect 32953 47240 32965 47243
rect 32732 47212 32965 47240
rect 32732 47200 32738 47212
rect 32953 47209 32965 47212
rect 32999 47209 33011 47243
rect 32953 47203 33011 47209
rect 33060 47212 33275 47240
rect 28902 47132 28908 47184
rect 28960 47172 28966 47184
rect 33060 47172 33088 47212
rect 28960 47144 33088 47172
rect 33247 47172 33275 47212
rect 33778 47200 33784 47252
rect 33836 47240 33842 47252
rect 34149 47243 34207 47249
rect 34149 47240 34161 47243
rect 33836 47212 34161 47240
rect 33836 47200 33842 47212
rect 34149 47209 34161 47212
rect 34195 47240 34207 47243
rect 35802 47240 35808 47252
rect 34195 47212 35808 47240
rect 34195 47209 34207 47212
rect 34149 47203 34207 47209
rect 35802 47200 35808 47212
rect 35860 47200 35866 47252
rect 35342 47172 35348 47184
rect 33247 47144 33456 47172
rect 35303 47144 35348 47172
rect 28960 47132 28966 47144
rect 27706 47064 27712 47116
rect 27764 47104 27770 47116
rect 28169 47107 28227 47113
rect 28169 47104 28181 47107
rect 27764 47076 28181 47104
rect 27764 47064 27770 47076
rect 28169 47073 28181 47076
rect 28215 47104 28227 47107
rect 28534 47104 28540 47116
rect 28215 47076 28540 47104
rect 28215 47073 28227 47076
rect 28169 47067 28227 47073
rect 28534 47064 28540 47076
rect 28592 47104 28598 47116
rect 28994 47104 29000 47116
rect 28592 47076 29000 47104
rect 28592 47064 28598 47076
rect 28994 47064 29000 47076
rect 29052 47064 29058 47116
rect 29454 47064 29460 47116
rect 29512 47104 29518 47116
rect 29825 47107 29883 47113
rect 29825 47104 29837 47107
rect 29512 47076 29837 47104
rect 29512 47064 29518 47076
rect 29825 47073 29837 47076
rect 29871 47104 29883 47107
rect 30190 47104 30196 47116
rect 29871 47076 30196 47104
rect 29871 47073 29883 47076
rect 29825 47067 29883 47073
rect 30190 47064 30196 47076
rect 30248 47104 30254 47116
rect 32490 47104 32496 47116
rect 30248 47076 31156 47104
rect 32451 47076 32496 47104
rect 30248 47064 30254 47076
rect 27430 47036 27436 47048
rect 27391 47008 27436 47036
rect 27430 46996 27436 47008
rect 27488 46996 27494 47048
rect 28813 47039 28871 47045
rect 28813 47005 28825 47039
rect 28859 47036 28871 47039
rect 29546 47036 29552 47048
rect 28859 47008 29552 47036
rect 28859 47005 28871 47008
rect 28813 46999 28871 47005
rect 29546 46996 29552 47008
rect 29604 46996 29610 47048
rect 29917 47039 29975 47045
rect 29917 47005 29929 47039
rect 29963 47005 29975 47039
rect 29917 46999 29975 47005
rect 30101 47039 30159 47045
rect 30101 47005 30113 47039
rect 30147 47036 30159 47039
rect 30742 47036 30748 47048
rect 30147 47008 30748 47036
rect 30147 47005 30159 47008
rect 30101 46999 30159 47005
rect 27341 46971 27399 46977
rect 27341 46968 27353 46971
rect 27264 46940 27353 46968
rect 27341 46937 27353 46940
rect 27387 46937 27399 46971
rect 27614 46968 27620 46980
rect 27341 46931 27399 46937
rect 27448 46940 27620 46968
rect 27448 46900 27476 46940
rect 27614 46928 27620 46940
rect 27672 46968 27678 46980
rect 28442 46968 28448 46980
rect 27672 46940 28448 46968
rect 27672 46928 27678 46940
rect 28442 46928 28448 46940
rect 28500 46968 28506 46980
rect 28997 46971 29055 46977
rect 28500 46940 28948 46968
rect 28500 46928 28506 46940
rect 26344 46872 27476 46900
rect 28920 46900 28948 46940
rect 28997 46937 29009 46971
rect 29043 46968 29055 46971
rect 29178 46968 29184 46980
rect 29043 46940 29184 46968
rect 29043 46937 29055 46940
rect 28997 46931 29055 46937
rect 29178 46928 29184 46940
rect 29236 46968 29242 46980
rect 29932 46968 29960 46999
rect 30742 46996 30748 47008
rect 30800 46996 30806 47048
rect 31128 47045 31156 47076
rect 32490 47064 32496 47076
rect 32548 47064 32554 47116
rect 33226 47104 33232 47116
rect 33060 47076 33232 47104
rect 31113 47039 31171 47045
rect 31113 47005 31125 47039
rect 31159 47036 31171 47039
rect 31294 47036 31300 47048
rect 31159 47008 31300 47036
rect 31159 47005 31171 47008
rect 31113 46999 31171 47005
rect 31294 46996 31300 47008
rect 31352 46996 31358 47048
rect 32214 47036 32220 47048
rect 32175 47008 32220 47036
rect 32214 46996 32220 47008
rect 32272 46996 32278 47048
rect 32309 47039 32367 47045
rect 32309 47005 32321 47039
rect 32355 47036 32367 47039
rect 33060 47036 33088 47076
rect 33226 47064 33232 47076
rect 33284 47064 33290 47116
rect 33428 47104 33456 47144
rect 35342 47132 35348 47144
rect 35400 47132 35406 47184
rect 37182 47104 37188 47116
rect 33428 47076 37188 47104
rect 33134 47045 33140 47048
rect 32355 47008 33088 47036
rect 32355 47005 32367 47008
rect 32309 46999 32367 47005
rect 33132 46999 33140 47045
rect 33192 47036 33198 47048
rect 33428 47045 33456 47076
rect 37182 47064 37188 47076
rect 37240 47104 37246 47116
rect 37461 47107 37519 47113
rect 37461 47104 37473 47107
rect 37240 47076 37473 47104
rect 37240 47064 37246 47076
rect 37461 47073 37473 47076
rect 37507 47073 37519 47107
rect 37461 47067 37519 47073
rect 33612 47045 33666 47046
rect 33428 47039 33507 47045
rect 33192 47008 33232 47036
rect 33428 47008 33461 47039
rect 33134 46996 33140 46999
rect 33192 46996 33198 47008
rect 33449 47005 33461 47008
rect 33495 47005 33507 47039
rect 33449 46999 33507 47005
rect 33572 47039 33666 47045
rect 33572 47005 33584 47039
rect 33618 47036 33666 47039
rect 33962 47036 33968 47048
rect 33618 47008 33968 47036
rect 33618 47005 33630 47008
rect 33572 46999 33630 47005
rect 33962 46996 33968 47008
rect 34020 47036 34026 47048
rect 36909 47039 36967 47045
rect 36909 47036 36921 47039
rect 34020 47008 36921 47036
rect 34020 46996 34026 47008
rect 36909 47005 36921 47008
rect 36955 47005 36967 47039
rect 36909 46999 36967 47005
rect 29236 46940 29960 46968
rect 29236 46928 29242 46940
rect 30650 46928 30656 46980
rect 30708 46968 30714 46980
rect 30926 46968 30932 46980
rect 30708 46940 30932 46968
rect 30708 46928 30714 46940
rect 30926 46928 30932 46940
rect 30984 46928 30990 46980
rect 31662 46968 31668 46980
rect 31623 46940 31668 46968
rect 31662 46928 31668 46940
rect 31720 46928 31726 46980
rect 33226 46968 33232 46980
rect 33187 46940 33232 46968
rect 33226 46928 33232 46940
rect 33284 46928 33290 46980
rect 33318 46928 33324 46980
rect 33376 46968 33382 46980
rect 33376 46940 33421 46968
rect 33376 46928 33382 46940
rect 34054 46928 34060 46980
rect 34112 46968 34118 46980
rect 34701 46971 34759 46977
rect 34701 46968 34713 46971
rect 34112 46940 34713 46968
rect 34112 46928 34118 46940
rect 34701 46937 34713 46940
rect 34747 46937 34759 46971
rect 35897 46971 35955 46977
rect 35897 46968 35909 46971
rect 34701 46931 34759 46937
rect 34808 46940 35909 46968
rect 30834 46900 30840 46912
rect 28920 46872 30840 46900
rect 30834 46860 30840 46872
rect 30892 46860 30898 46912
rect 32493 46903 32551 46909
rect 32493 46869 32505 46903
rect 32539 46900 32551 46903
rect 33134 46900 33140 46912
rect 32539 46872 33140 46900
rect 32539 46869 32551 46872
rect 32493 46863 32551 46869
rect 33134 46860 33140 46872
rect 33192 46860 33198 46912
rect 34606 46860 34612 46912
rect 34664 46900 34670 46912
rect 34808 46900 34836 46940
rect 35897 46937 35909 46940
rect 35943 46937 35955 46971
rect 35897 46931 35955 46937
rect 34664 46872 34836 46900
rect 36449 46903 36507 46909
rect 34664 46860 34670 46872
rect 36449 46869 36461 46903
rect 36495 46900 36507 46903
rect 36538 46900 36544 46912
rect 36495 46872 36544 46900
rect 36495 46869 36507 46872
rect 36449 46863 36507 46869
rect 36538 46860 36544 46872
rect 36596 46860 36602 46912
rect 1104 46810 54372 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 54372 46810
rect 1104 46736 54372 46758
rect 21269 46699 21327 46705
rect 21269 46665 21281 46699
rect 21315 46696 21327 46699
rect 22094 46696 22100 46708
rect 21315 46668 22100 46696
rect 21315 46665 21327 46668
rect 21269 46659 21327 46665
rect 22094 46656 22100 46668
rect 22152 46696 22158 46708
rect 22370 46696 22376 46708
rect 22152 46668 22376 46696
rect 22152 46656 22158 46668
rect 22370 46656 22376 46668
rect 22428 46656 22434 46708
rect 23569 46699 23627 46705
rect 23569 46665 23581 46699
rect 23615 46696 23627 46699
rect 23750 46696 23756 46708
rect 23615 46668 23756 46696
rect 23615 46665 23627 46668
rect 23569 46659 23627 46665
rect 23750 46656 23756 46668
rect 23808 46656 23814 46708
rect 24581 46699 24639 46705
rect 24581 46665 24593 46699
rect 24627 46696 24639 46699
rect 24854 46696 24860 46708
rect 24627 46668 24860 46696
rect 24627 46665 24639 46668
rect 24581 46659 24639 46665
rect 24854 46656 24860 46668
rect 24912 46656 24918 46708
rect 25222 46656 25228 46708
rect 25280 46696 25286 46708
rect 25501 46699 25559 46705
rect 25501 46696 25513 46699
rect 25280 46668 25513 46696
rect 25280 46656 25286 46668
rect 25501 46665 25513 46668
rect 25547 46665 25559 46699
rect 29178 46696 29184 46708
rect 29139 46668 29184 46696
rect 25501 46659 25559 46665
rect 29178 46656 29184 46668
rect 29236 46656 29242 46708
rect 30009 46699 30067 46705
rect 30009 46665 30021 46699
rect 30055 46696 30067 46699
rect 30190 46696 30196 46708
rect 30055 46668 30196 46696
rect 30055 46665 30067 46668
rect 30009 46659 30067 46665
rect 30190 46656 30196 46668
rect 30248 46656 30254 46708
rect 30742 46696 30748 46708
rect 30703 46668 30748 46696
rect 30742 46656 30748 46668
rect 30800 46656 30806 46708
rect 31202 46656 31208 46708
rect 31260 46696 31266 46708
rect 31297 46699 31355 46705
rect 31297 46696 31309 46699
rect 31260 46668 31309 46696
rect 31260 46656 31266 46668
rect 31297 46665 31309 46668
rect 31343 46665 31355 46699
rect 31297 46659 31355 46665
rect 32677 46699 32735 46705
rect 32677 46665 32689 46699
rect 32723 46696 32735 46699
rect 33318 46696 33324 46708
rect 32723 46668 33324 46696
rect 32723 46665 32735 46668
rect 32677 46659 32735 46665
rect 33318 46656 33324 46668
rect 33376 46656 33382 46708
rect 34054 46696 34060 46708
rect 34015 46668 34060 46696
rect 34054 46656 34060 46668
rect 34112 46656 34118 46708
rect 26234 46588 26240 46640
rect 26292 46628 26298 46640
rect 26292 46600 27292 46628
rect 26292 46588 26298 46600
rect 23382 46560 23388 46572
rect 23343 46532 23388 46560
rect 23382 46520 23388 46532
rect 23440 46520 23446 46572
rect 23566 46560 23572 46572
rect 23527 46532 23572 46560
rect 23566 46520 23572 46532
rect 23624 46520 23630 46572
rect 24213 46563 24271 46569
rect 24213 46529 24225 46563
rect 24259 46560 24271 46563
rect 24394 46560 24400 46572
rect 24259 46532 24400 46560
rect 24259 46529 24271 46532
rect 24213 46523 24271 46529
rect 24394 46520 24400 46532
rect 24452 46520 24458 46572
rect 25682 46560 25688 46572
rect 25643 46532 25688 46560
rect 25682 46520 25688 46532
rect 25740 46520 25746 46572
rect 25866 46560 25872 46572
rect 25827 46532 25872 46560
rect 25866 46520 25872 46532
rect 25924 46520 25930 46572
rect 26510 46520 26516 46572
rect 26568 46560 26574 46572
rect 27264 46569 27292 46600
rect 27522 46588 27528 46640
rect 27580 46628 27586 46640
rect 28813 46631 28871 46637
rect 28813 46628 28825 46631
rect 27580 46600 28825 46628
rect 27580 46588 27586 46600
rect 28813 46597 28825 46600
rect 28859 46597 28871 46631
rect 28813 46591 28871 46597
rect 29029 46631 29087 46637
rect 29029 46597 29041 46631
rect 29075 46628 29087 46631
rect 29454 46628 29460 46640
rect 29075 46600 29460 46628
rect 29075 46597 29087 46600
rect 29029 46591 29087 46597
rect 26973 46563 27031 46569
rect 26973 46560 26985 46563
rect 26568 46532 26985 46560
rect 26568 46520 26574 46532
rect 26973 46529 26985 46532
rect 27019 46529 27031 46563
rect 26973 46523 27031 46529
rect 27249 46563 27307 46569
rect 27249 46529 27261 46563
rect 27295 46529 27307 46563
rect 28828 46560 28856 46591
rect 29454 46588 29460 46600
rect 29512 46628 29518 46640
rect 29914 46628 29920 46640
rect 29512 46600 29920 46628
rect 29512 46588 29518 46600
rect 29914 46588 29920 46600
rect 29972 46588 29978 46640
rect 32950 46588 32956 46640
rect 33008 46628 33014 46640
rect 33137 46631 33195 46637
rect 33137 46628 33149 46631
rect 33008 46600 33149 46628
rect 33008 46588 33014 46600
rect 33137 46597 33149 46600
rect 33183 46597 33195 46631
rect 33137 46591 33195 46597
rect 34609 46631 34667 46637
rect 34609 46597 34621 46631
rect 34655 46628 34667 46631
rect 35434 46628 35440 46640
rect 34655 46600 35440 46628
rect 34655 46597 34667 46600
rect 34609 46591 34667 46597
rect 35434 46588 35440 46600
rect 35492 46588 35498 46640
rect 29641 46563 29699 46569
rect 29641 46560 29653 46563
rect 28828 46532 29653 46560
rect 27249 46523 27307 46529
rect 29641 46529 29653 46532
rect 29687 46560 29699 46563
rect 29730 46560 29736 46572
rect 29687 46532 29736 46560
rect 29687 46529 29699 46532
rect 29641 46523 29699 46529
rect 29730 46520 29736 46532
rect 29788 46520 29794 46572
rect 29822 46520 29828 46572
rect 29880 46560 29886 46572
rect 30098 46560 30104 46572
rect 29880 46532 30104 46560
rect 29880 46520 29886 46532
rect 30098 46520 30104 46532
rect 30156 46520 30162 46572
rect 30653 46563 30711 46569
rect 30653 46529 30665 46563
rect 30699 46529 30711 46563
rect 30834 46560 30840 46572
rect 30795 46532 30840 46560
rect 30653 46523 30711 46529
rect 20717 46495 20775 46501
rect 20717 46461 20729 46495
rect 20763 46492 20775 46495
rect 21818 46492 21824 46504
rect 20763 46464 21824 46492
rect 20763 46461 20775 46464
rect 20717 46455 20775 46461
rect 21818 46452 21824 46464
rect 21876 46492 21882 46504
rect 22278 46492 22284 46504
rect 21876 46464 22284 46492
rect 21876 46452 21882 46464
rect 22278 46452 22284 46464
rect 22336 46452 22342 46504
rect 24305 46495 24363 46501
rect 24305 46461 24317 46495
rect 24351 46492 24363 46495
rect 24486 46492 24492 46504
rect 24351 46464 24492 46492
rect 24351 46461 24363 46464
rect 24305 46455 24363 46461
rect 24486 46452 24492 46464
rect 24544 46452 24550 46504
rect 25498 46452 25504 46504
rect 25556 46492 25562 46504
rect 25777 46495 25835 46501
rect 25777 46492 25789 46495
rect 25556 46464 25789 46492
rect 25556 46452 25562 46464
rect 25777 46461 25789 46464
rect 25823 46461 25835 46495
rect 25777 46455 25835 46461
rect 25961 46495 26019 46501
rect 25961 46461 25973 46495
rect 26007 46461 26019 46495
rect 25961 46455 26019 46461
rect 30193 46495 30251 46501
rect 30193 46461 30205 46495
rect 30239 46492 30251 46495
rect 30668 46492 30696 46523
rect 30834 46520 30840 46532
rect 30892 46520 30898 46572
rect 32122 46520 32128 46572
rect 32180 46560 32186 46572
rect 32309 46563 32367 46569
rect 32309 46560 32321 46563
rect 32180 46532 32321 46560
rect 32180 46520 32186 46532
rect 32309 46529 32321 46532
rect 32355 46529 32367 46563
rect 32309 46523 32367 46529
rect 32582 46520 32588 46572
rect 32640 46560 32646 46572
rect 33321 46563 33379 46569
rect 33321 46560 33333 46563
rect 32640 46532 33333 46560
rect 32640 46520 32646 46532
rect 33321 46529 33333 46532
rect 33367 46529 33379 46563
rect 33594 46560 33600 46572
rect 33555 46532 33600 46560
rect 33321 46523 33379 46529
rect 33594 46520 33600 46532
rect 33652 46520 33658 46572
rect 34790 46560 34796 46572
rect 34751 46532 34796 46560
rect 34790 46520 34796 46532
rect 34848 46560 34854 46572
rect 35802 46560 35808 46572
rect 34848 46532 35808 46560
rect 34848 46520 34854 46532
rect 35802 46520 35808 46532
rect 35860 46560 35866 46572
rect 35989 46563 36047 46569
rect 35989 46560 36001 46563
rect 35860 46532 36001 46560
rect 35860 46520 35866 46532
rect 35989 46529 36001 46532
rect 36035 46529 36047 46563
rect 53377 46563 53435 46569
rect 53377 46560 53389 46563
rect 35989 46523 36047 46529
rect 52840 46532 53389 46560
rect 32214 46492 32220 46504
rect 30239 46464 32220 46492
rect 30239 46461 30251 46464
rect 30193 46455 30251 46461
rect 22833 46427 22891 46433
rect 22833 46424 22845 46427
rect 22066 46396 22845 46424
rect 18874 46356 18880 46368
rect 18835 46328 18880 46356
rect 18874 46316 18880 46328
rect 18932 46316 18938 46368
rect 19334 46316 19340 46368
rect 19392 46356 19398 46368
rect 19981 46359 20039 46365
rect 19392 46328 19437 46356
rect 19392 46316 19398 46328
rect 19981 46325 19993 46359
rect 20027 46356 20039 46359
rect 20990 46356 20996 46368
rect 20027 46328 20996 46356
rect 20027 46325 20039 46328
rect 19981 46319 20039 46325
rect 20990 46316 20996 46328
rect 21048 46356 21054 46368
rect 22066 46356 22094 46396
rect 22833 46393 22845 46396
rect 22879 46424 22891 46427
rect 23198 46424 23204 46436
rect 22879 46396 23204 46424
rect 22879 46393 22891 46396
rect 22833 46387 22891 46393
rect 23198 46384 23204 46396
rect 23256 46384 23262 46436
rect 25406 46384 25412 46436
rect 25464 46424 25470 46436
rect 25976 46424 26004 46455
rect 32214 46452 32220 46464
rect 32272 46452 32278 46504
rect 33134 46452 33140 46504
rect 33192 46492 33198 46504
rect 33505 46495 33563 46501
rect 33505 46492 33517 46495
rect 33192 46464 33517 46492
rect 33192 46452 33198 46464
rect 33505 46461 33517 46464
rect 33551 46461 33563 46495
rect 33505 46455 33563 46461
rect 33870 46452 33876 46504
rect 33928 46492 33934 46504
rect 35529 46495 35587 46501
rect 35529 46492 35541 46495
rect 33928 46464 35541 46492
rect 33928 46452 33934 46464
rect 35529 46461 35541 46464
rect 35575 46492 35587 46495
rect 36630 46492 36636 46504
rect 35575 46464 36636 46492
rect 35575 46461 35587 46464
rect 35529 46455 35587 46461
rect 36630 46452 36636 46464
rect 36688 46452 36694 46504
rect 52840 46501 52868 46532
rect 53377 46529 53389 46532
rect 53423 46529 53435 46563
rect 53377 46523 53435 46529
rect 52825 46495 52883 46501
rect 52825 46492 52837 46495
rect 41386 46464 52837 46492
rect 25464 46396 26004 46424
rect 25464 46384 25470 46396
rect 30926 46384 30932 46436
rect 30984 46424 30990 46436
rect 31662 46424 31668 46436
rect 30984 46396 31668 46424
rect 30984 46384 30990 46396
rect 31662 46384 31668 46396
rect 31720 46424 31726 46436
rect 41386 46424 41414 46464
rect 52825 46461 52837 46464
rect 52871 46461 52883 46495
rect 52825 46455 52883 46461
rect 31720 46396 41414 46424
rect 31720 46384 31726 46396
rect 22370 46356 22376 46368
rect 21048 46328 22094 46356
rect 22331 46328 22376 46356
rect 21048 46316 21054 46328
rect 22370 46316 22376 46328
rect 22428 46316 22434 46368
rect 26418 46316 26424 46368
rect 26476 46356 26482 46368
rect 26694 46356 26700 46368
rect 26476 46328 26700 46356
rect 26476 46316 26482 46328
rect 26694 46316 26700 46328
rect 26752 46356 26758 46368
rect 27065 46359 27123 46365
rect 27065 46356 27077 46359
rect 26752 46328 27077 46356
rect 26752 46316 26758 46328
rect 27065 46325 27077 46328
rect 27111 46325 27123 46359
rect 27430 46356 27436 46368
rect 27391 46328 27436 46356
rect 27065 46319 27123 46325
rect 27430 46316 27436 46328
rect 27488 46316 27494 46368
rect 28258 46356 28264 46368
rect 28219 46328 28264 46356
rect 28258 46316 28264 46328
rect 28316 46316 28322 46368
rect 28994 46356 29000 46368
rect 28907 46328 29000 46356
rect 28994 46316 29000 46328
rect 29052 46356 29058 46368
rect 29822 46356 29828 46368
rect 29052 46328 29828 46356
rect 29052 46316 29058 46328
rect 29822 46316 29828 46328
rect 29880 46316 29886 46368
rect 32398 46316 32404 46368
rect 32456 46356 32462 46368
rect 34790 46356 34796 46368
rect 32456 46328 34796 46356
rect 32456 46316 32462 46328
rect 34790 46316 34796 46328
rect 34848 46316 34854 46368
rect 34977 46359 35035 46365
rect 34977 46325 34989 46359
rect 35023 46356 35035 46359
rect 35342 46356 35348 46368
rect 35023 46328 35348 46356
rect 35023 46325 35035 46328
rect 34977 46319 35035 46325
rect 35342 46316 35348 46328
rect 35400 46316 35406 46368
rect 36630 46356 36636 46368
rect 36591 46328 36636 46356
rect 36630 46316 36636 46328
rect 36688 46316 36694 46368
rect 37274 46356 37280 46368
rect 37235 46328 37280 46356
rect 37274 46316 37280 46328
rect 37332 46316 37338 46368
rect 37826 46356 37832 46368
rect 37787 46328 37832 46356
rect 37826 46316 37832 46328
rect 37884 46316 37890 46368
rect 53558 46356 53564 46368
rect 53519 46328 53564 46356
rect 53558 46316 53564 46328
rect 53616 46316 53622 46368
rect 1104 46266 54372 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 54372 46266
rect 1104 46192 54372 46214
rect 18693 46155 18751 46161
rect 18693 46121 18705 46155
rect 18739 46152 18751 46155
rect 19334 46152 19340 46164
rect 18739 46124 19340 46152
rect 18739 46121 18751 46124
rect 18693 46115 18751 46121
rect 19334 46112 19340 46124
rect 19392 46112 19398 46164
rect 20990 46152 20996 46164
rect 20951 46124 20996 46152
rect 20990 46112 20996 46124
rect 21048 46112 21054 46164
rect 23198 46152 23204 46164
rect 23159 46124 23204 46152
rect 23198 46112 23204 46124
rect 23256 46112 23262 46164
rect 25038 46112 25044 46164
rect 25096 46152 25102 46164
rect 25593 46155 25651 46161
rect 25593 46152 25605 46155
rect 25096 46124 25605 46152
rect 25096 46112 25102 46124
rect 25593 46121 25605 46124
rect 25639 46121 25651 46155
rect 29546 46152 29552 46164
rect 29507 46124 29552 46152
rect 25593 46115 25651 46121
rect 29546 46112 29552 46124
rect 29604 46112 29610 46164
rect 32309 46155 32367 46161
rect 32309 46121 32321 46155
rect 32355 46152 32367 46155
rect 32398 46152 32404 46164
rect 32355 46124 32404 46152
rect 32355 46121 32367 46124
rect 32309 46115 32367 46121
rect 32398 46112 32404 46124
rect 32456 46112 32462 46164
rect 32490 46112 32496 46164
rect 32548 46152 32554 46164
rect 32953 46155 33011 46161
rect 32953 46152 32965 46155
rect 32548 46124 32965 46152
rect 32548 46112 32554 46124
rect 32953 46121 32965 46124
rect 32999 46121 33011 46155
rect 33134 46152 33140 46164
rect 33095 46124 33140 46152
rect 32953 46115 33011 46121
rect 33134 46112 33140 46124
rect 33192 46112 33198 46164
rect 32122 46044 32128 46096
rect 32180 46084 32186 46096
rect 34238 46084 34244 46096
rect 32180 46056 34244 46084
rect 32180 46044 32186 46056
rect 34238 46044 34244 46056
rect 34296 46044 34302 46096
rect 34514 46044 34520 46096
rect 34572 46084 34578 46096
rect 35161 46087 35219 46093
rect 35161 46084 35173 46087
rect 34572 46056 35173 46084
rect 34572 46044 34578 46056
rect 35161 46053 35173 46056
rect 35207 46053 35219 46087
rect 35161 46047 35219 46053
rect 18874 45976 18880 46028
rect 18932 46016 18938 46028
rect 19242 46016 19248 46028
rect 18932 45988 19248 46016
rect 18932 45976 18938 45988
rect 19242 45976 19248 45988
rect 19300 46016 19306 46028
rect 22189 46019 22247 46025
rect 19300 45988 21680 46016
rect 19300 45976 19306 45988
rect 19978 45908 19984 45960
rect 20036 45948 20042 45960
rect 20165 45951 20223 45957
rect 20165 45948 20177 45951
rect 20036 45920 20177 45948
rect 20036 45908 20042 45920
rect 20165 45917 20177 45920
rect 20211 45917 20223 45951
rect 20165 45911 20223 45917
rect 20349 45951 20407 45957
rect 20349 45917 20361 45951
rect 20395 45948 20407 45951
rect 20990 45948 20996 45960
rect 20395 45920 20996 45948
rect 20395 45917 20407 45920
rect 20349 45911 20407 45917
rect 20990 45908 20996 45920
rect 21048 45908 21054 45960
rect 21652 45957 21680 45988
rect 22189 45985 22201 46019
rect 22235 46016 22247 46019
rect 27982 46016 27988 46028
rect 22235 45988 25728 46016
rect 27943 45988 27988 46016
rect 22235 45985 22247 45988
rect 22189 45979 22247 45985
rect 21637 45951 21695 45957
rect 21637 45917 21649 45951
rect 21683 45948 21695 45951
rect 22830 45948 22836 45960
rect 21683 45920 22836 45948
rect 21683 45917 21695 45920
rect 21637 45911 21695 45917
rect 22830 45908 22836 45920
rect 22888 45908 22894 45960
rect 25130 45908 25136 45960
rect 25188 45948 25194 45960
rect 25700 45957 25728 45988
rect 27982 45976 27988 45988
rect 28040 45976 28046 46028
rect 30834 45976 30840 46028
rect 30892 46016 30898 46028
rect 33226 46016 33232 46028
rect 30892 45988 33232 46016
rect 30892 45976 30898 45988
rect 33226 45976 33232 45988
rect 33284 46016 33290 46028
rect 33870 46016 33876 46028
rect 33284 45988 33876 46016
rect 33284 45976 33290 45988
rect 33870 45976 33876 45988
rect 33928 45976 33934 46028
rect 34072 45988 35020 46016
rect 25501 45951 25559 45957
rect 25501 45948 25513 45951
rect 25188 45920 25513 45948
rect 25188 45908 25194 45920
rect 25501 45917 25513 45920
rect 25547 45917 25559 45951
rect 25501 45911 25559 45917
rect 25685 45951 25743 45957
rect 25685 45917 25697 45951
rect 25731 45948 25743 45951
rect 26326 45948 26332 45960
rect 25731 45920 26332 45948
rect 25731 45917 25743 45920
rect 25685 45911 25743 45917
rect 26326 45908 26332 45920
rect 26384 45908 26390 45960
rect 27430 45908 27436 45960
rect 27488 45948 27494 45960
rect 27718 45951 27776 45957
rect 27718 45948 27730 45951
rect 27488 45920 27730 45948
rect 27488 45908 27494 45920
rect 27718 45917 27730 45920
rect 27764 45917 27776 45951
rect 29730 45948 29736 45960
rect 29691 45920 29736 45948
rect 27718 45911 27776 45917
rect 29730 45908 29736 45920
rect 29788 45908 29794 45960
rect 29822 45908 29828 45960
rect 29880 45948 29886 45960
rect 30190 45948 30196 45960
rect 29880 45920 30196 45948
rect 29880 45908 29886 45920
rect 30190 45908 30196 45920
rect 30248 45908 30254 45960
rect 34072 45957 34100 45988
rect 34992 45960 35020 45988
rect 30377 45951 30435 45957
rect 30377 45917 30389 45951
rect 30423 45948 30435 45951
rect 33321 45951 33379 45957
rect 30423 45920 31524 45948
rect 30423 45917 30435 45920
rect 30377 45911 30435 45917
rect 1578 45840 1584 45892
rect 1636 45880 1642 45892
rect 1857 45883 1915 45889
rect 1857 45880 1869 45883
rect 1636 45852 1869 45880
rect 1636 45840 1642 45852
rect 1857 45849 1869 45852
rect 1903 45849 1915 45883
rect 1857 45843 1915 45849
rect 2041 45883 2099 45889
rect 2041 45849 2053 45883
rect 2087 45880 2099 45883
rect 2130 45880 2136 45892
rect 2087 45852 2136 45880
rect 2087 45849 2099 45852
rect 2041 45843 2099 45849
rect 2130 45840 2136 45852
rect 2188 45840 2194 45892
rect 19705 45883 19763 45889
rect 19705 45849 19717 45883
rect 19751 45880 19763 45883
rect 21818 45880 21824 45892
rect 19751 45852 21824 45880
rect 19751 45849 19763 45852
rect 19705 45843 19763 45849
rect 21818 45840 21824 45852
rect 21876 45840 21882 45892
rect 23845 45883 23903 45889
rect 23845 45849 23857 45883
rect 23891 45880 23903 45883
rect 24394 45880 24400 45892
rect 23891 45852 24400 45880
rect 23891 45849 23903 45852
rect 23845 45843 23903 45849
rect 24394 45840 24400 45852
rect 24452 45840 24458 45892
rect 29454 45840 29460 45892
rect 29512 45880 29518 45892
rect 29549 45883 29607 45889
rect 29549 45880 29561 45883
rect 29512 45852 29561 45880
rect 29512 45840 29518 45852
rect 29549 45849 29561 45852
rect 29595 45849 29607 45883
rect 30926 45880 30932 45892
rect 29549 45843 29607 45849
rect 30300 45852 30932 45880
rect 17494 45812 17500 45824
rect 17455 45784 17500 45812
rect 17494 45772 17500 45784
rect 17552 45772 17558 45824
rect 20070 45772 20076 45824
rect 20128 45812 20134 45824
rect 20257 45815 20315 45821
rect 20257 45812 20269 45815
rect 20128 45784 20269 45812
rect 20128 45772 20134 45784
rect 20257 45781 20269 45784
rect 20303 45781 20315 45815
rect 20257 45775 20315 45781
rect 22741 45815 22799 45821
rect 22741 45781 22753 45815
rect 22787 45812 22799 45815
rect 23014 45812 23020 45824
rect 22787 45784 23020 45812
rect 22787 45781 22799 45784
rect 22741 45775 22799 45781
rect 23014 45772 23020 45784
rect 23072 45772 23078 45824
rect 24486 45812 24492 45824
rect 24447 45784 24492 45812
rect 24486 45772 24492 45784
rect 24544 45772 24550 45824
rect 25041 45815 25099 45821
rect 25041 45781 25053 45815
rect 25087 45812 25099 45815
rect 26605 45815 26663 45821
rect 26605 45812 26617 45815
rect 25087 45784 26617 45812
rect 25087 45781 25099 45784
rect 25041 45775 25099 45781
rect 26605 45781 26617 45784
rect 26651 45812 26663 45815
rect 26694 45812 26700 45824
rect 26651 45784 26700 45812
rect 26651 45781 26663 45784
rect 26605 45775 26663 45781
rect 26694 45772 26700 45784
rect 26752 45772 26758 45824
rect 28350 45772 28356 45824
rect 28408 45812 28414 45824
rect 28445 45815 28503 45821
rect 28445 45812 28457 45815
rect 28408 45784 28457 45812
rect 28408 45772 28414 45784
rect 28445 45781 28457 45784
rect 28491 45812 28503 45815
rect 30300 45812 30328 45852
rect 30926 45840 30932 45852
rect 30984 45840 30990 45892
rect 31496 45824 31524 45920
rect 33321 45917 33333 45951
rect 33367 45917 33379 45951
rect 33321 45911 33379 45917
rect 34057 45951 34115 45957
rect 34057 45917 34069 45951
rect 34103 45917 34115 45951
rect 34057 45911 34115 45917
rect 32122 45880 32128 45892
rect 32083 45852 32128 45880
rect 32122 45840 32128 45852
rect 32180 45840 32186 45892
rect 32214 45840 32220 45892
rect 32272 45880 32278 45892
rect 32325 45883 32383 45889
rect 32325 45880 32337 45883
rect 32272 45852 32337 45880
rect 32272 45840 32278 45852
rect 32325 45849 32337 45852
rect 32371 45849 32383 45883
rect 32325 45843 32383 45849
rect 33336 45824 33364 45911
rect 34146 45908 34152 45960
rect 34204 45948 34210 45960
rect 34204 45920 34560 45948
rect 34204 45908 34210 45920
rect 33410 45840 33416 45892
rect 33468 45880 33474 45892
rect 33870 45880 33876 45892
rect 33468 45852 33876 45880
rect 33468 45840 33474 45852
rect 33870 45840 33876 45852
rect 33928 45840 33934 45892
rect 28491 45784 30328 45812
rect 28491 45781 28503 45784
rect 28445 45775 28503 45781
rect 30374 45772 30380 45824
rect 30432 45812 30438 45824
rect 30837 45815 30895 45821
rect 30837 45812 30849 45815
rect 30432 45784 30849 45812
rect 30432 45772 30438 45784
rect 30837 45781 30849 45784
rect 30883 45781 30895 45815
rect 31478 45812 31484 45824
rect 31439 45784 31484 45812
rect 30837 45775 30895 45781
rect 31478 45772 31484 45784
rect 31536 45772 31542 45824
rect 32493 45815 32551 45821
rect 32493 45781 32505 45815
rect 32539 45812 32551 45815
rect 33318 45812 33324 45824
rect 32539 45784 33324 45812
rect 32539 45781 32551 45784
rect 32493 45775 32551 45781
rect 33318 45772 33324 45784
rect 33376 45772 33382 45824
rect 33594 45772 33600 45824
rect 33652 45812 33658 45824
rect 33965 45815 34023 45821
rect 33965 45812 33977 45815
rect 33652 45784 33977 45812
rect 33652 45772 33658 45784
rect 33965 45781 33977 45784
rect 34011 45812 34023 45815
rect 34422 45812 34428 45824
rect 34011 45784 34428 45812
rect 34011 45781 34023 45784
rect 33965 45775 34023 45781
rect 34422 45772 34428 45784
rect 34480 45772 34486 45824
rect 34532 45812 34560 45920
rect 34606 45908 34612 45960
rect 34664 45948 34670 45960
rect 34701 45951 34759 45957
rect 34701 45948 34713 45951
rect 34664 45920 34713 45948
rect 34664 45908 34670 45920
rect 34701 45917 34713 45920
rect 34747 45917 34759 45951
rect 34974 45948 34980 45960
rect 34935 45920 34980 45948
rect 34701 45911 34759 45917
rect 34974 45908 34980 45920
rect 35032 45908 35038 45960
rect 35434 45908 35440 45960
rect 35492 45948 35498 45960
rect 35621 45951 35679 45957
rect 35621 45948 35633 45951
rect 35492 45920 35633 45948
rect 35492 45908 35498 45920
rect 35621 45917 35633 45920
rect 35667 45917 35679 45951
rect 35802 45948 35808 45960
rect 35763 45920 35808 45948
rect 35621 45911 35679 45917
rect 35802 45908 35808 45920
rect 35860 45948 35866 45960
rect 36265 45951 36323 45957
rect 36265 45948 36277 45951
rect 35860 45920 36277 45948
rect 35860 45908 35866 45920
rect 36265 45917 36277 45920
rect 36311 45948 36323 45951
rect 37369 45951 37427 45957
rect 37369 45948 37381 45951
rect 36311 45920 37381 45948
rect 36311 45917 36323 45920
rect 36265 45911 36323 45917
rect 37369 45917 37381 45920
rect 37415 45948 37427 45951
rect 37826 45948 37832 45960
rect 37415 45920 37832 45948
rect 37415 45917 37427 45920
rect 37369 45911 37427 45917
rect 37826 45908 37832 45920
rect 37884 45908 37890 45960
rect 34606 45812 34612 45824
rect 34532 45784 34612 45812
rect 34606 45772 34612 45784
rect 34664 45812 34670 45824
rect 34793 45815 34851 45821
rect 34793 45812 34805 45815
rect 34664 45784 34805 45812
rect 34664 45772 34670 45784
rect 34793 45781 34805 45784
rect 34839 45781 34851 45815
rect 35802 45812 35808 45824
rect 35763 45784 35808 45812
rect 34793 45775 34851 45781
rect 35802 45772 35808 45784
rect 35860 45772 35866 45824
rect 36538 45772 36544 45824
rect 36596 45812 36602 45824
rect 36909 45815 36967 45821
rect 36909 45812 36921 45815
rect 36596 45784 36921 45812
rect 36596 45772 36602 45784
rect 36909 45781 36921 45784
rect 36955 45812 36967 45815
rect 37734 45812 37740 45824
rect 36955 45784 37740 45812
rect 36955 45781 36967 45784
rect 36909 45775 36967 45781
rect 37734 45772 37740 45784
rect 37792 45772 37798 45824
rect 1104 45722 54372 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 54372 45722
rect 1104 45648 54372 45670
rect 1578 45608 1584 45620
rect 1539 45580 1584 45608
rect 1578 45568 1584 45580
rect 1636 45568 1642 45620
rect 20073 45611 20131 45617
rect 20073 45577 20085 45611
rect 20119 45608 20131 45611
rect 20990 45608 20996 45620
rect 20119 45580 20996 45608
rect 20119 45577 20131 45580
rect 20073 45571 20131 45577
rect 20990 45568 20996 45580
rect 21048 45568 21054 45620
rect 22370 45568 22376 45620
rect 22428 45608 22434 45620
rect 22465 45611 22523 45617
rect 22465 45608 22477 45611
rect 22428 45580 22477 45608
rect 22428 45568 22434 45580
rect 22465 45577 22477 45580
rect 22511 45608 22523 45611
rect 24394 45608 24400 45620
rect 22511 45580 24400 45608
rect 22511 45577 22523 45580
rect 22465 45571 22523 45577
rect 24394 45568 24400 45580
rect 24452 45568 24458 45620
rect 25130 45568 25136 45620
rect 25188 45608 25194 45620
rect 27433 45611 27491 45617
rect 27433 45608 27445 45611
rect 25188 45580 27445 45608
rect 25188 45568 25194 45580
rect 27433 45577 27445 45580
rect 27479 45608 27491 45611
rect 27522 45608 27528 45620
rect 27479 45580 27528 45608
rect 27479 45577 27491 45580
rect 27433 45571 27491 45577
rect 27522 45568 27528 45580
rect 27580 45568 27586 45620
rect 30285 45611 30343 45617
rect 30285 45577 30297 45611
rect 30331 45608 30343 45611
rect 31202 45608 31208 45620
rect 30331 45580 31208 45608
rect 30331 45577 30343 45580
rect 30285 45571 30343 45577
rect 31202 45568 31208 45580
rect 31260 45568 31266 45620
rect 32122 45568 32128 45620
rect 32180 45608 32186 45620
rect 32309 45611 32367 45617
rect 32309 45608 32321 45611
rect 32180 45580 32321 45608
rect 32180 45568 32186 45580
rect 32309 45577 32321 45580
rect 32355 45577 32367 45611
rect 32309 45571 32367 45577
rect 33594 45568 33600 45620
rect 33652 45617 33658 45620
rect 33652 45611 33671 45617
rect 33659 45577 33671 45611
rect 33652 45571 33671 45577
rect 33652 45568 33658 45571
rect 33870 45568 33876 45620
rect 33928 45608 33934 45620
rect 34425 45611 34483 45617
rect 34425 45608 34437 45611
rect 33928 45580 34437 45608
rect 33928 45568 33934 45580
rect 34425 45577 34437 45580
rect 34471 45577 34483 45611
rect 34425 45571 34483 45577
rect 34609 45611 34667 45617
rect 34609 45577 34621 45611
rect 34655 45608 34667 45611
rect 34974 45608 34980 45620
rect 34655 45580 34980 45608
rect 34655 45577 34667 45580
rect 34609 45571 34667 45577
rect 34974 45568 34980 45580
rect 35032 45608 35038 45620
rect 35437 45611 35495 45617
rect 35437 45608 35449 45611
rect 35032 45580 35449 45608
rect 35032 45568 35038 45580
rect 35437 45577 35449 45580
rect 35483 45577 35495 45611
rect 35437 45571 35495 45577
rect 19429 45543 19487 45549
rect 19429 45509 19441 45543
rect 19475 45540 19487 45543
rect 21358 45540 21364 45552
rect 19475 45512 21364 45540
rect 19475 45509 19487 45512
rect 19429 45503 19487 45509
rect 18690 45432 18696 45484
rect 18748 45472 18754 45484
rect 19337 45475 19395 45481
rect 19337 45472 19349 45475
rect 18748 45444 19349 45472
rect 18748 45432 18754 45444
rect 19337 45441 19349 45444
rect 19383 45441 19395 45475
rect 19337 45435 19395 45441
rect 19521 45475 19579 45481
rect 19521 45441 19533 45475
rect 19567 45441 19579 45475
rect 19978 45472 19984 45484
rect 19939 45444 19984 45472
rect 19521 45435 19579 45441
rect 17770 45404 17776 45416
rect 17683 45376 17776 45404
rect 17770 45364 17776 45376
rect 17828 45404 17834 45416
rect 19426 45404 19432 45416
rect 17828 45376 19432 45404
rect 17828 45364 17834 45376
rect 19426 45364 19432 45376
rect 19484 45364 19490 45416
rect 19536 45404 19564 45435
rect 19978 45432 19984 45444
rect 20036 45432 20042 45484
rect 20732 45481 20760 45512
rect 21358 45500 21364 45512
rect 21416 45500 21422 45552
rect 25774 45540 25780 45552
rect 23124 45512 23888 45540
rect 25735 45512 25780 45540
rect 20257 45475 20315 45481
rect 20257 45441 20269 45475
rect 20303 45441 20315 45475
rect 20257 45435 20315 45441
rect 20717 45475 20775 45481
rect 20717 45441 20729 45475
rect 20763 45441 20775 45475
rect 20717 45435 20775 45441
rect 20901 45475 20959 45481
rect 20901 45441 20913 45475
rect 20947 45472 20959 45475
rect 21450 45472 21456 45484
rect 20947 45444 21456 45472
rect 20947 45441 20959 45444
rect 20901 45435 20959 45441
rect 20272 45404 20300 45435
rect 21450 45432 21456 45444
rect 21508 45432 21514 45484
rect 22738 45432 22744 45484
rect 22796 45472 22802 45484
rect 23124 45481 23152 45512
rect 22925 45475 22983 45481
rect 22925 45472 22937 45475
rect 22796 45444 22937 45472
rect 22796 45432 22802 45444
rect 22925 45441 22937 45444
rect 22971 45441 22983 45475
rect 22925 45435 22983 45441
rect 23109 45475 23167 45481
rect 23109 45441 23121 45475
rect 23155 45441 23167 45475
rect 23569 45475 23627 45481
rect 23569 45472 23581 45475
rect 23109 45435 23167 45441
rect 23216 45444 23581 45472
rect 21174 45404 21180 45416
rect 19536 45376 21180 45404
rect 21174 45364 21180 45376
rect 21232 45364 21238 45416
rect 22094 45364 22100 45416
rect 22152 45404 22158 45416
rect 22370 45404 22376 45416
rect 22152 45376 22376 45404
rect 22152 45364 22158 45376
rect 22370 45364 22376 45376
rect 22428 45364 22434 45416
rect 23017 45407 23075 45413
rect 23017 45373 23029 45407
rect 23063 45404 23075 45407
rect 23216 45404 23244 45444
rect 23569 45441 23581 45444
rect 23615 45472 23627 45475
rect 23750 45472 23756 45484
rect 23615 45444 23756 45472
rect 23615 45441 23627 45444
rect 23569 45435 23627 45441
rect 23750 45432 23756 45444
rect 23808 45432 23814 45484
rect 23860 45413 23888 45512
rect 25774 45500 25780 45512
rect 25832 45500 25838 45552
rect 26326 45540 26332 45552
rect 26287 45512 26332 45540
rect 26326 45500 26332 45512
rect 26384 45540 26390 45552
rect 28074 45540 28080 45552
rect 26384 45512 28080 45540
rect 26384 45500 26390 45512
rect 28074 45500 28080 45512
rect 28132 45540 28138 45552
rect 28902 45540 28908 45552
rect 28132 45512 28908 45540
rect 28132 45500 28138 45512
rect 28902 45500 28908 45512
rect 28960 45540 28966 45552
rect 29089 45543 29147 45549
rect 29089 45540 29101 45543
rect 28960 45512 29101 45540
rect 28960 45500 28966 45512
rect 29089 45509 29101 45512
rect 29135 45509 29147 45543
rect 29089 45503 29147 45509
rect 32398 45500 32404 45552
rect 32456 45540 32462 45552
rect 32493 45543 32551 45549
rect 32493 45540 32505 45543
rect 32456 45512 32505 45540
rect 32456 45500 32462 45512
rect 32493 45509 32505 45512
rect 32539 45509 32551 45543
rect 32493 45503 32551 45509
rect 33413 45543 33471 45549
rect 33413 45509 33425 45543
rect 33459 45540 33471 45543
rect 34054 45540 34060 45552
rect 33459 45512 34060 45540
rect 33459 45509 33471 45512
rect 33413 45503 33471 45509
rect 34054 45500 34060 45512
rect 34112 45540 34118 45552
rect 34330 45540 34336 45552
rect 34112 45512 34336 45540
rect 34112 45500 34118 45512
rect 34330 45500 34336 45512
rect 34388 45500 34394 45552
rect 36265 45543 36323 45549
rect 36265 45540 36277 45543
rect 34440 45512 36277 45540
rect 26694 45432 26700 45484
rect 26752 45472 26758 45484
rect 27249 45475 27307 45481
rect 27249 45472 27261 45475
rect 26752 45444 27261 45472
rect 26752 45432 26758 45444
rect 27249 45441 27261 45444
rect 27295 45441 27307 45475
rect 32214 45472 32220 45484
rect 32175 45444 32220 45472
rect 27249 45435 27307 45441
rect 32214 45432 32220 45444
rect 32272 45432 32278 45484
rect 32582 45432 32588 45484
rect 32640 45472 32646 45484
rect 34440 45472 34468 45512
rect 36265 45509 36277 45512
rect 36311 45540 36323 45543
rect 37274 45540 37280 45552
rect 36311 45512 37280 45540
rect 36311 45509 36323 45512
rect 36265 45503 36323 45509
rect 37274 45500 37280 45512
rect 37332 45500 37338 45552
rect 32640 45444 34468 45472
rect 32640 45432 32646 45444
rect 34606 45432 34612 45484
rect 34664 45472 34670 45484
rect 34701 45475 34759 45481
rect 34701 45472 34713 45475
rect 34664 45444 34713 45472
rect 34664 45432 34670 45444
rect 34701 45441 34713 45444
rect 34747 45441 34759 45475
rect 34701 45435 34759 45441
rect 35342 45432 35348 45484
rect 35400 45472 35406 45484
rect 35621 45475 35679 45481
rect 35621 45472 35633 45475
rect 35400 45444 35633 45472
rect 35400 45432 35406 45444
rect 35621 45441 35633 45444
rect 35667 45441 35679 45475
rect 35621 45435 35679 45441
rect 23063 45376 23244 45404
rect 23845 45407 23903 45413
rect 23063 45373 23075 45376
rect 23017 45367 23075 45373
rect 23845 45373 23857 45407
rect 23891 45404 23903 45407
rect 23934 45404 23940 45416
rect 23891 45376 23940 45404
rect 23891 45373 23903 45376
rect 23845 45367 23903 45373
rect 23934 45364 23940 45376
rect 23992 45364 23998 45416
rect 25317 45407 25375 45413
rect 25317 45373 25329 45407
rect 25363 45404 25375 45407
rect 26878 45404 26884 45416
rect 25363 45376 26884 45404
rect 25363 45373 25375 45376
rect 25317 45367 25375 45373
rect 26878 45364 26884 45376
rect 26936 45364 26942 45416
rect 34330 45404 34336 45416
rect 34291 45376 34336 45404
rect 34330 45364 34336 45376
rect 34388 45364 34394 45416
rect 34790 45364 34796 45416
rect 34848 45404 34854 45416
rect 35802 45404 35808 45416
rect 34848 45376 34893 45404
rect 35763 45376 35808 45404
rect 34848 45364 34854 45376
rect 35802 45364 35808 45376
rect 35860 45364 35866 45416
rect 18325 45339 18383 45345
rect 18325 45305 18337 45339
rect 18371 45336 18383 45339
rect 19242 45336 19248 45348
rect 18371 45308 19248 45336
rect 18371 45305 18383 45308
rect 18325 45299 18383 45305
rect 19242 45296 19248 45308
rect 19300 45296 19306 45348
rect 20257 45339 20315 45345
rect 20257 45305 20269 45339
rect 20303 45336 20315 45339
rect 20714 45336 20720 45348
rect 20303 45308 20720 45336
rect 20303 45305 20315 45308
rect 20257 45299 20315 45305
rect 20714 45296 20720 45308
rect 20772 45336 20778 45348
rect 21634 45336 21640 45348
rect 20772 45308 21640 45336
rect 20772 45296 20778 45308
rect 21634 45296 21640 45308
rect 21692 45296 21698 45348
rect 22554 45296 22560 45348
rect 22612 45336 22618 45348
rect 27798 45336 27804 45348
rect 22612 45308 27804 45336
rect 22612 45296 22618 45308
rect 27798 45296 27804 45308
rect 27856 45296 27862 45348
rect 32493 45339 32551 45345
rect 32493 45305 32505 45339
rect 32539 45336 32551 45339
rect 33134 45336 33140 45348
rect 32539 45308 33140 45336
rect 32539 45305 32551 45308
rect 32493 45299 32551 45305
rect 33134 45296 33140 45308
rect 33192 45296 33198 45348
rect 33502 45296 33508 45348
rect 33560 45336 33566 45348
rect 33781 45339 33839 45345
rect 33781 45336 33793 45339
rect 33560 45308 33793 45336
rect 33560 45296 33566 45308
rect 33781 45305 33793 45308
rect 33827 45305 33839 45339
rect 33781 45299 33839 45305
rect 35342 45296 35348 45348
rect 35400 45336 35406 45348
rect 37829 45339 37887 45345
rect 37829 45336 37841 45339
rect 35400 45308 37841 45336
rect 35400 45296 35406 45308
rect 37829 45305 37841 45308
rect 37875 45305 37887 45339
rect 37829 45299 37887 45305
rect 17221 45271 17279 45277
rect 17221 45237 17233 45271
rect 17267 45268 17279 45271
rect 18046 45268 18052 45280
rect 17267 45240 18052 45268
rect 17267 45237 17279 45240
rect 17221 45231 17279 45237
rect 18046 45228 18052 45240
rect 18104 45228 18110 45280
rect 18874 45268 18880 45280
rect 18835 45240 18880 45268
rect 18874 45228 18880 45240
rect 18932 45228 18938 45280
rect 20809 45271 20867 45277
rect 20809 45237 20821 45271
rect 20855 45268 20867 45271
rect 21082 45268 21088 45280
rect 20855 45240 21088 45268
rect 20855 45237 20867 45240
rect 20809 45231 20867 45237
rect 21082 45228 21088 45240
rect 21140 45228 21146 45280
rect 21913 45271 21971 45277
rect 21913 45237 21925 45271
rect 21959 45268 21971 45271
rect 22094 45268 22100 45280
rect 21959 45240 22100 45268
rect 21959 45237 21971 45240
rect 21913 45231 21971 45237
rect 22094 45228 22100 45240
rect 22152 45228 22158 45280
rect 23382 45228 23388 45280
rect 23440 45268 23446 45280
rect 23661 45271 23719 45277
rect 23661 45268 23673 45271
rect 23440 45240 23673 45268
rect 23440 45228 23446 45240
rect 23661 45237 23673 45240
rect 23707 45237 23719 45271
rect 23661 45231 23719 45237
rect 23753 45271 23811 45277
rect 23753 45237 23765 45271
rect 23799 45268 23811 45271
rect 24210 45268 24216 45280
rect 23799 45240 24216 45268
rect 23799 45237 23811 45240
rect 23753 45231 23811 45237
rect 24210 45228 24216 45240
rect 24268 45228 24274 45280
rect 24394 45228 24400 45280
rect 24452 45268 24458 45280
rect 24765 45271 24823 45277
rect 24765 45268 24777 45271
rect 24452 45240 24777 45268
rect 24452 45228 24458 45240
rect 24765 45237 24777 45240
rect 24811 45268 24823 45271
rect 25406 45268 25412 45280
rect 24811 45240 25412 45268
rect 24811 45237 24823 45240
rect 24765 45231 24823 45237
rect 25406 45228 25412 45240
rect 25464 45228 25470 45280
rect 27522 45228 27528 45280
rect 27580 45268 27586 45280
rect 27985 45271 28043 45277
rect 27985 45268 27997 45271
rect 27580 45240 27997 45268
rect 27580 45228 27586 45240
rect 27985 45237 27997 45240
rect 28031 45268 28043 45271
rect 28350 45268 28356 45280
rect 28031 45240 28356 45268
rect 28031 45237 28043 45240
rect 27985 45231 28043 45237
rect 28350 45228 28356 45240
rect 28408 45228 28414 45280
rect 28442 45228 28448 45280
rect 28500 45268 28506 45280
rect 28537 45271 28595 45277
rect 28537 45268 28549 45271
rect 28500 45240 28549 45268
rect 28500 45228 28506 45240
rect 28537 45237 28549 45240
rect 28583 45237 28595 45271
rect 28537 45231 28595 45237
rect 28994 45228 29000 45280
rect 29052 45268 29058 45280
rect 29641 45271 29699 45277
rect 29641 45268 29653 45271
rect 29052 45240 29653 45268
rect 29052 45228 29058 45240
rect 29641 45237 29653 45240
rect 29687 45268 29699 45271
rect 30374 45268 30380 45280
rect 29687 45240 30380 45268
rect 29687 45237 29699 45240
rect 29641 45231 29699 45237
rect 30374 45228 30380 45240
rect 30432 45228 30438 45280
rect 33597 45271 33655 45277
rect 33597 45237 33609 45271
rect 33643 45268 33655 45271
rect 34514 45268 34520 45280
rect 33643 45240 34520 45268
rect 33643 45237 33655 45240
rect 33597 45231 33655 45237
rect 34514 45228 34520 45240
rect 34572 45228 34578 45280
rect 34698 45228 34704 45280
rect 34756 45268 34762 45280
rect 34977 45271 35035 45277
rect 34977 45268 34989 45271
rect 34756 45240 34989 45268
rect 34756 45228 34762 45240
rect 34977 45237 34989 45240
rect 35023 45237 35035 45271
rect 34977 45231 35035 45237
rect 37369 45271 37427 45277
rect 37369 45237 37381 45271
rect 37415 45268 37427 45271
rect 37734 45268 37740 45280
rect 37415 45240 37740 45268
rect 37415 45237 37427 45240
rect 37369 45231 37427 45237
rect 37734 45228 37740 45240
rect 37792 45228 37798 45280
rect 1104 45178 54372 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 54372 45178
rect 1104 45104 54372 45126
rect 16485 45067 16543 45073
rect 16485 45033 16497 45067
rect 16531 45064 16543 45067
rect 16942 45064 16948 45076
rect 16531 45036 16948 45064
rect 16531 45033 16543 45036
rect 16485 45027 16543 45033
rect 16942 45024 16948 45036
rect 17000 45064 17006 45076
rect 17310 45064 17316 45076
rect 17000 45036 17316 45064
rect 17000 45024 17006 45036
rect 17310 45024 17316 45036
rect 17368 45064 17374 45076
rect 17770 45064 17776 45076
rect 17368 45036 17776 45064
rect 17368 45024 17374 45036
rect 17770 45024 17776 45036
rect 17828 45024 17834 45076
rect 19242 45064 19248 45076
rect 19203 45036 19248 45064
rect 19242 45024 19248 45036
rect 19300 45024 19306 45076
rect 19426 45024 19432 45076
rect 19484 45064 19490 45076
rect 22554 45064 22560 45076
rect 19484 45036 22560 45064
rect 19484 45024 19490 45036
rect 22554 45024 22560 45036
rect 22612 45024 22618 45076
rect 22738 45064 22744 45076
rect 22699 45036 22744 45064
rect 22738 45024 22744 45036
rect 22796 45024 22802 45076
rect 23106 45064 23112 45076
rect 23019 45036 23112 45064
rect 23106 45024 23112 45036
rect 23164 45064 23170 45076
rect 27522 45064 27528 45076
rect 23164 45036 27528 45064
rect 23164 45024 23170 45036
rect 27522 45024 27528 45036
rect 27580 45024 27586 45076
rect 28258 45024 28264 45076
rect 28316 45064 28322 45076
rect 30926 45064 30932 45076
rect 28316 45036 30604 45064
rect 30887 45036 30932 45064
rect 28316 45024 28322 45036
rect 17218 44996 17224 45008
rect 17179 44968 17224 44996
rect 17218 44956 17224 44968
rect 17276 44956 17282 45008
rect 18693 44999 18751 45005
rect 18693 44965 18705 44999
rect 18739 44996 18751 44999
rect 19334 44996 19340 45008
rect 18739 44968 19340 44996
rect 18739 44965 18751 44968
rect 18693 44959 18751 44965
rect 19334 44956 19340 44968
rect 19392 44996 19398 45008
rect 21177 44999 21235 45005
rect 19392 44968 21036 44996
rect 19392 44956 19398 44968
rect 19812 44937 19840 44968
rect 21008 44940 21036 44968
rect 21177 44965 21189 44999
rect 21223 44996 21235 44999
rect 22922 44996 22928 45008
rect 21223 44968 22928 44996
rect 21223 44965 21235 44968
rect 21177 44959 21235 44965
rect 22922 44956 22928 44968
rect 22980 44956 22986 45008
rect 19797 44931 19855 44937
rect 15856 44900 17724 44928
rect 15286 44724 15292 44736
rect 15247 44696 15292 44724
rect 15286 44684 15292 44696
rect 15344 44724 15350 44736
rect 15856 44733 15884 44900
rect 16850 44820 16856 44872
rect 16908 44860 16914 44872
rect 16945 44863 17003 44869
rect 16945 44860 16957 44863
rect 16908 44832 16957 44860
rect 16908 44820 16914 44832
rect 16945 44829 16957 44832
rect 16991 44829 17003 44863
rect 17494 44860 17500 44872
rect 16945 44823 17003 44829
rect 17052 44832 17500 44860
rect 16298 44752 16304 44804
rect 16356 44792 16362 44804
rect 17052 44792 17080 44832
rect 17494 44820 17500 44832
rect 17552 44860 17558 44872
rect 17696 44869 17724 44900
rect 19797 44897 19809 44931
rect 19843 44897 19855 44931
rect 20898 44928 20904 44940
rect 20859 44900 20904 44928
rect 19797 44891 19855 44897
rect 20898 44888 20904 44900
rect 20956 44888 20962 44940
rect 20990 44888 20996 44940
rect 21048 44928 21054 44940
rect 23124 44928 23152 45024
rect 30576 45008 30604 45036
rect 30926 45024 30932 45036
rect 30984 45024 30990 45076
rect 31941 45067 31999 45073
rect 31941 45033 31953 45067
rect 31987 45064 31999 45067
rect 33962 45064 33968 45076
rect 31987 45036 33968 45064
rect 31987 45033 31999 45036
rect 31941 45027 31999 45033
rect 23845 44999 23903 45005
rect 23845 44965 23857 44999
rect 23891 44996 23903 44999
rect 24489 44999 24547 45005
rect 24489 44996 24501 44999
rect 23891 44968 24501 44996
rect 23891 44965 23903 44968
rect 23845 44959 23903 44965
rect 24489 44965 24501 44968
rect 24535 44965 24547 44999
rect 24489 44959 24547 44965
rect 24670 44956 24676 45008
rect 24728 44996 24734 45008
rect 24728 44968 24900 44996
rect 24728 44956 24734 44968
rect 23382 44928 23388 44940
rect 21048 44900 22048 44928
rect 21048 44888 21054 44900
rect 22020 44872 22048 44900
rect 22388 44900 23152 44928
rect 23343 44900 23388 44928
rect 17681 44863 17739 44869
rect 17552 44832 17632 44860
rect 17552 44820 17558 44832
rect 16356 44764 17080 44792
rect 16356 44752 16362 44764
rect 17126 44752 17132 44804
rect 17184 44792 17190 44804
rect 17221 44795 17279 44801
rect 17221 44792 17233 44795
rect 17184 44764 17233 44792
rect 17184 44752 17190 44764
rect 17221 44761 17233 44764
rect 17267 44761 17279 44795
rect 17604 44792 17632 44832
rect 17681 44829 17693 44863
rect 17727 44829 17739 44863
rect 17681 44823 17739 44829
rect 17865 44863 17923 44869
rect 17865 44829 17877 44863
rect 17911 44829 17923 44863
rect 19978 44860 19984 44872
rect 19939 44832 19984 44860
rect 17865 44823 17923 44829
rect 17880 44792 17908 44823
rect 19978 44820 19984 44832
rect 20036 44820 20042 44872
rect 20806 44860 20812 44872
rect 20767 44832 20812 44860
rect 20806 44820 20812 44832
rect 20864 44820 20870 44872
rect 21634 44860 21640 44872
rect 21595 44832 21640 44860
rect 21634 44820 21640 44832
rect 21692 44820 21698 44872
rect 21821 44863 21879 44869
rect 21821 44829 21833 44863
rect 21867 44829 21879 44863
rect 21821 44823 21879 44829
rect 18322 44792 18328 44804
rect 17604 44764 18328 44792
rect 17221 44755 17279 44761
rect 18322 44752 18328 44764
rect 18380 44752 18386 44804
rect 20070 44752 20076 44804
rect 20128 44792 20134 44804
rect 21836 44792 21864 44823
rect 22002 44820 22008 44872
rect 22060 44860 22066 44872
rect 22388 44869 22416 44900
rect 23382 44888 23388 44900
rect 23440 44888 23446 44940
rect 22373 44863 22431 44869
rect 22373 44860 22385 44863
rect 22060 44832 22385 44860
rect 22060 44820 22066 44832
rect 22373 44829 22385 44832
rect 22419 44829 22431 44863
rect 22373 44823 22431 44829
rect 22462 44820 22468 44872
rect 22520 44860 22526 44872
rect 22557 44863 22615 44869
rect 22557 44860 22569 44863
rect 22520 44832 22569 44860
rect 22520 44820 22526 44832
rect 22557 44829 22569 44832
rect 22603 44829 22615 44863
rect 22557 44823 22615 44829
rect 23555 44863 23613 44869
rect 23555 44829 23567 44863
rect 23601 44860 23613 44863
rect 23750 44860 23756 44872
rect 23601 44832 23756 44860
rect 23601 44829 23613 44832
rect 23555 44823 23613 44829
rect 23750 44820 23756 44832
rect 23808 44820 23814 44872
rect 24394 44860 24400 44872
rect 24355 44832 24400 44860
rect 24394 44820 24400 44832
rect 24452 44820 24458 44872
rect 24670 44860 24676 44872
rect 24631 44832 24676 44860
rect 24670 44820 24676 44832
rect 24728 44820 24734 44872
rect 24765 44863 24823 44869
rect 24765 44829 24777 44863
rect 24811 44829 24823 44863
rect 24872 44860 24900 44968
rect 25314 44956 25320 45008
rect 25372 44996 25378 45008
rect 25409 44999 25467 45005
rect 25409 44996 25421 44999
rect 25372 44968 25421 44996
rect 25372 44956 25378 44968
rect 25409 44965 25421 44968
rect 25455 44965 25467 44999
rect 25409 44959 25467 44965
rect 26973 44999 27031 45005
rect 26973 44965 26985 44999
rect 27019 44996 27031 44999
rect 28902 44996 28908 45008
rect 27019 44968 28908 44996
rect 27019 44965 27031 44968
rect 26973 44959 27031 44965
rect 28902 44956 28908 44968
rect 28960 44956 28966 45008
rect 28997 44999 29055 45005
rect 28997 44965 29009 44999
rect 29043 44965 29055 44999
rect 28997 44959 29055 44965
rect 24949 44931 25007 44937
rect 24949 44897 24961 44931
rect 24995 44928 25007 44931
rect 24995 44900 28764 44928
rect 24995 44897 25007 44900
rect 24949 44891 25007 44897
rect 25682 44860 25688 44872
rect 24872 44832 25544 44860
rect 25643 44832 25688 44860
rect 24765 44823 24823 44829
rect 20128 44764 21864 44792
rect 20128 44752 20134 44764
rect 22922 44752 22928 44804
rect 22980 44792 22986 44804
rect 24780 44792 24808 44823
rect 25406 44792 25412 44804
rect 22980 44764 24808 44792
rect 25367 44764 25412 44792
rect 22980 44752 22986 44764
rect 25406 44752 25412 44764
rect 25464 44752 25470 44804
rect 25516 44792 25544 44832
rect 25682 44820 25688 44832
rect 25740 44820 25746 44872
rect 27249 44863 27307 44869
rect 27249 44829 27261 44863
rect 27295 44860 27307 44863
rect 27706 44860 27712 44872
rect 27295 44832 27712 44860
rect 27295 44829 27307 44832
rect 27249 44823 27307 44829
rect 27706 44820 27712 44832
rect 27764 44820 27770 44872
rect 28736 44869 28764 44900
rect 28721 44863 28779 44869
rect 28721 44829 28733 44863
rect 28767 44829 28779 44863
rect 29012 44860 29040 44959
rect 30558 44956 30564 45008
rect 30616 44996 30622 45008
rect 31956 44996 31984 45027
rect 33962 45024 33968 45036
rect 34020 45024 34026 45076
rect 34790 45024 34796 45076
rect 34848 45064 34854 45076
rect 35989 45067 36047 45073
rect 35989 45064 36001 45067
rect 34848 45036 36001 45064
rect 34848 45024 34854 45036
rect 35989 45033 36001 45036
rect 36035 45033 36047 45067
rect 35989 45027 36047 45033
rect 37274 45024 37280 45076
rect 37332 45064 37338 45076
rect 37829 45067 37887 45073
rect 37829 45064 37841 45067
rect 37332 45036 37841 45064
rect 37332 45024 37338 45036
rect 37829 45033 37841 45036
rect 37875 45064 37887 45067
rect 38102 45064 38108 45076
rect 37875 45036 38108 45064
rect 37875 45033 37887 45036
rect 37829 45027 37887 45033
rect 38102 45024 38108 45036
rect 38160 45024 38166 45076
rect 30616 44968 31984 44996
rect 30616 44956 30622 44968
rect 34422 44956 34428 45008
rect 34480 44996 34486 45008
rect 34480 44968 35020 44996
rect 34480 44956 34486 44968
rect 29549 44931 29607 44937
rect 29549 44897 29561 44931
rect 29595 44928 29607 44931
rect 30006 44928 30012 44940
rect 29595 44900 30012 44928
rect 29595 44897 29607 44900
rect 29549 44891 29607 44897
rect 30006 44888 30012 44900
rect 30064 44888 30070 44940
rect 34992 44937 35020 44968
rect 33597 44931 33655 44937
rect 33597 44897 33609 44931
rect 33643 44928 33655 44931
rect 34701 44931 34759 44937
rect 34701 44928 34713 44931
rect 33643 44900 34713 44928
rect 33643 44897 33655 44900
rect 33597 44891 33655 44897
rect 34701 44897 34713 44900
rect 34747 44897 34759 44931
rect 34701 44891 34759 44897
rect 34977 44931 35035 44937
rect 34977 44897 34989 44931
rect 35023 44897 35035 44931
rect 34977 44891 35035 44897
rect 35161 44931 35219 44937
rect 35161 44897 35173 44931
rect 35207 44928 35219 44931
rect 35342 44928 35348 44940
rect 35207 44900 35348 44928
rect 35207 44897 35219 44900
rect 35161 44891 35219 44897
rect 35342 44888 35348 44900
rect 35400 44928 35406 44940
rect 35618 44928 35624 44940
rect 35400 44900 35624 44928
rect 35400 44888 35406 44900
rect 35618 44888 35624 44900
rect 35676 44888 35682 44940
rect 36725 44931 36783 44937
rect 36725 44928 36737 44931
rect 35728 44900 36737 44928
rect 35728 44872 35756 44900
rect 36725 44897 36737 44900
rect 36771 44897 36783 44931
rect 36725 44891 36783 44897
rect 29825 44863 29883 44869
rect 29825 44860 29837 44863
rect 29012 44832 29837 44860
rect 28721 44823 28779 44829
rect 29825 44829 29837 44832
rect 29871 44829 29883 44863
rect 29825 44823 29883 44829
rect 31941 44863 31999 44869
rect 31941 44829 31953 44863
rect 31987 44860 31999 44863
rect 32490 44860 32496 44872
rect 31987 44832 32496 44860
rect 31987 44829 31999 44832
rect 31941 44823 31999 44829
rect 32490 44820 32496 44832
rect 32548 44820 32554 44872
rect 32585 44863 32643 44869
rect 32585 44829 32597 44863
rect 32631 44829 32643 44863
rect 32766 44860 32772 44872
rect 32727 44832 32772 44860
rect 32585 44823 32643 44829
rect 26418 44792 26424 44804
rect 25516 44764 26424 44792
rect 26418 44752 26424 44764
rect 26476 44752 26482 44804
rect 26878 44752 26884 44804
rect 26936 44792 26942 44804
rect 26973 44795 27031 44801
rect 26973 44792 26985 44795
rect 26936 44764 26985 44792
rect 26936 44752 26942 44764
rect 26973 44761 26985 44764
rect 27019 44792 27031 44795
rect 28258 44792 28264 44804
rect 27019 44764 28264 44792
rect 27019 44761 27031 44764
rect 26973 44755 27031 44761
rect 28258 44752 28264 44764
rect 28316 44792 28322 44804
rect 28997 44795 29055 44801
rect 28997 44792 29009 44795
rect 28316 44764 29009 44792
rect 28316 44752 28322 44764
rect 28997 44761 29009 44764
rect 29043 44761 29055 44795
rect 32600 44792 32628 44823
rect 32766 44820 32772 44832
rect 32824 44820 32830 44872
rect 33413 44863 33471 44869
rect 33413 44829 33425 44863
rect 33459 44860 33471 44863
rect 33502 44860 33508 44872
rect 33459 44832 33508 44860
rect 33459 44829 33471 44832
rect 33413 44823 33471 44829
rect 33502 44820 33508 44832
rect 33560 44820 33566 44872
rect 33689 44863 33747 44869
rect 33689 44829 33701 44863
rect 33735 44860 33747 44863
rect 34146 44860 34152 44872
rect 33735 44832 34152 44860
rect 33735 44829 33747 44832
rect 33689 44823 33747 44829
rect 34146 44820 34152 44832
rect 34204 44820 34210 44872
rect 34330 44820 34336 44872
rect 34388 44860 34394 44872
rect 34882 44860 34888 44872
rect 34388 44832 34888 44860
rect 34388 44820 34394 44832
rect 34882 44820 34888 44832
rect 34940 44820 34946 44872
rect 35069 44863 35127 44869
rect 35069 44829 35081 44863
rect 35115 44829 35127 44863
rect 35710 44860 35716 44872
rect 35623 44832 35716 44860
rect 35069 44823 35127 44829
rect 33318 44792 33324 44804
rect 32600 44764 33324 44792
rect 28997 44755 29055 44761
rect 33318 44752 33324 44764
rect 33376 44792 33382 44804
rect 33594 44792 33600 44804
rect 33376 44764 33600 44792
rect 33376 44752 33382 44764
rect 33594 44752 33600 44764
rect 33652 44752 33658 44804
rect 34790 44752 34796 44804
rect 34848 44792 34854 44804
rect 35084 44792 35112 44823
rect 35710 44820 35716 44832
rect 35768 44820 35774 44872
rect 36170 44860 36176 44872
rect 36131 44832 36176 44860
rect 36170 44820 36176 44832
rect 36228 44820 36234 44872
rect 36538 44820 36544 44872
rect 36596 44860 36602 44872
rect 36633 44863 36691 44869
rect 36633 44860 36645 44863
rect 36596 44832 36645 44860
rect 36596 44820 36602 44832
rect 36633 44829 36645 44832
rect 36679 44829 36691 44863
rect 36633 44823 36691 44829
rect 36817 44863 36875 44869
rect 36817 44829 36829 44863
rect 36863 44829 36875 44863
rect 36817 44823 36875 44829
rect 35802 44792 35808 44804
rect 34848 44764 35808 44792
rect 34848 44752 34854 44764
rect 35802 44752 35808 44764
rect 35860 44752 35866 44804
rect 36262 44752 36268 44804
rect 36320 44792 36326 44804
rect 36832 44792 36860 44823
rect 37277 44795 37335 44801
rect 37277 44792 37289 44795
rect 36320 44764 37289 44792
rect 36320 44752 36326 44764
rect 37277 44761 37289 44764
rect 37323 44792 37335 44795
rect 38381 44795 38439 44801
rect 38381 44792 38393 44795
rect 37323 44764 38393 44792
rect 37323 44761 37335 44764
rect 37277 44755 37335 44761
rect 38381 44761 38393 44764
rect 38427 44792 38439 44795
rect 38427 44764 38654 44792
rect 38427 44761 38439 44764
rect 38381 44755 38439 44761
rect 15841 44727 15899 44733
rect 15841 44724 15853 44727
rect 15344 44696 15853 44724
rect 15344 44684 15350 44696
rect 15841 44693 15853 44696
rect 15887 44693 15899 44727
rect 15841 44687 15899 44693
rect 17037 44727 17095 44733
rect 17037 44693 17049 44727
rect 17083 44724 17095 44727
rect 17586 44724 17592 44736
rect 17083 44696 17592 44724
rect 17083 44693 17095 44696
rect 17037 44687 17095 44693
rect 17586 44684 17592 44696
rect 17644 44684 17650 44736
rect 17862 44724 17868 44736
rect 17823 44696 17868 44724
rect 17862 44684 17868 44696
rect 17920 44684 17926 44736
rect 20165 44727 20223 44733
rect 20165 44693 20177 44727
rect 20211 44724 20223 44727
rect 20254 44724 20260 44736
rect 20211 44696 20260 44724
rect 20211 44693 20223 44696
rect 20165 44687 20223 44693
rect 20254 44684 20260 44696
rect 20312 44684 20318 44736
rect 20990 44684 20996 44736
rect 21048 44724 21054 44736
rect 21729 44727 21787 44733
rect 21729 44724 21741 44727
rect 21048 44696 21741 44724
rect 21048 44684 21054 44696
rect 21729 44693 21741 44696
rect 21775 44693 21787 44727
rect 21729 44687 21787 44693
rect 23014 44684 23020 44736
rect 23072 44724 23078 44736
rect 24670 44724 24676 44736
rect 23072 44696 24676 44724
rect 23072 44684 23078 44696
rect 24670 44684 24676 44696
rect 24728 44684 24734 44736
rect 25038 44684 25044 44736
rect 25096 44724 25102 44736
rect 25593 44727 25651 44733
rect 25593 44724 25605 44727
rect 25096 44696 25605 44724
rect 25096 44684 25102 44696
rect 25593 44693 25605 44696
rect 25639 44693 25651 44727
rect 27154 44724 27160 44736
rect 27115 44696 27160 44724
rect 25593 44687 25651 44693
rect 27154 44684 27160 44696
rect 27212 44684 27218 44736
rect 28166 44724 28172 44736
rect 28127 44696 28172 44724
rect 28166 44684 28172 44696
rect 28224 44684 28230 44736
rect 28813 44727 28871 44733
rect 28813 44693 28825 44727
rect 28859 44724 28871 44727
rect 30834 44724 30840 44736
rect 28859 44696 30840 44724
rect 28859 44693 28871 44696
rect 28813 44687 28871 44693
rect 30834 44684 30840 44696
rect 30892 44684 30898 44736
rect 32306 44684 32312 44736
rect 32364 44724 32370 44736
rect 32677 44727 32735 44733
rect 32677 44724 32689 44727
rect 32364 44696 32689 44724
rect 32364 44684 32370 44696
rect 32677 44693 32689 44696
rect 32723 44693 32735 44727
rect 33226 44724 33232 44736
rect 33187 44696 33232 44724
rect 32677 44687 32735 44693
rect 33226 44684 33232 44696
rect 33284 44684 33290 44736
rect 38626 44724 38654 44764
rect 38933 44727 38991 44733
rect 38933 44724 38945 44727
rect 38626 44696 38945 44724
rect 38933 44693 38945 44696
rect 38979 44693 38991 44727
rect 38933 44687 38991 44693
rect 1104 44634 54372 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 54372 44634
rect 1104 44560 54372 44582
rect 19353 44523 19411 44529
rect 19353 44520 19365 44523
rect 18432 44492 19365 44520
rect 18432 44396 18460 44492
rect 19353 44489 19365 44492
rect 19399 44489 19411 44523
rect 19353 44483 19411 44489
rect 21082 44480 21088 44532
rect 21140 44520 21146 44532
rect 22021 44523 22079 44529
rect 22021 44520 22033 44523
rect 21140 44492 22033 44520
rect 21140 44480 21146 44492
rect 22021 44489 22033 44492
rect 22067 44489 22079 44523
rect 22021 44483 22079 44489
rect 23382 44480 23388 44532
rect 23440 44520 23446 44532
rect 25133 44523 25191 44529
rect 25133 44520 25145 44523
rect 23440 44492 25145 44520
rect 23440 44480 23446 44492
rect 25133 44489 25145 44492
rect 25179 44489 25191 44523
rect 25133 44483 25191 44489
rect 26421 44523 26479 44529
rect 26421 44489 26433 44523
rect 26467 44520 26479 44523
rect 27154 44520 27160 44532
rect 26467 44492 27160 44520
rect 26467 44489 26479 44492
rect 26421 44483 26479 44489
rect 27154 44480 27160 44492
rect 27212 44480 27218 44532
rect 30834 44520 30840 44532
rect 30795 44492 30840 44520
rect 30834 44480 30840 44492
rect 30892 44480 30898 44532
rect 33502 44520 33508 44532
rect 33463 44492 33508 44520
rect 33502 44480 33508 44492
rect 33560 44480 33566 44532
rect 34333 44523 34391 44529
rect 34333 44489 34345 44523
rect 34379 44520 34391 44523
rect 34790 44520 34796 44532
rect 34379 44492 34796 44520
rect 34379 44489 34391 44492
rect 34333 44483 34391 44489
rect 34790 44480 34796 44492
rect 34848 44480 34854 44532
rect 34882 44480 34888 44532
rect 34940 44520 34946 44532
rect 35345 44523 35403 44529
rect 35345 44520 35357 44523
rect 34940 44492 35357 44520
rect 34940 44480 34946 44492
rect 35345 44489 35357 44492
rect 35391 44489 35403 44523
rect 36170 44520 36176 44532
rect 36131 44492 36176 44520
rect 35345 44483 35403 44489
rect 36170 44480 36176 44492
rect 36228 44480 36234 44532
rect 36630 44480 36636 44532
rect 36688 44520 36694 44532
rect 37277 44523 37335 44529
rect 37277 44520 37289 44523
rect 36688 44492 37289 44520
rect 36688 44480 36694 44492
rect 37277 44489 37289 44492
rect 37323 44489 37335 44523
rect 37277 44483 37335 44489
rect 18693 44455 18751 44461
rect 18693 44421 18705 44455
rect 18739 44452 18751 44455
rect 19153 44455 19211 44461
rect 19153 44452 19165 44455
rect 18739 44424 19165 44452
rect 18739 44421 18751 44424
rect 18693 44415 18751 44421
rect 19153 44421 19165 44424
rect 19199 44452 19211 44455
rect 19242 44452 19248 44464
rect 19199 44424 19248 44452
rect 19199 44421 19211 44424
rect 19153 44415 19211 44421
rect 19242 44412 19248 44424
rect 19300 44412 19306 44464
rect 20070 44452 20076 44464
rect 20031 44424 20076 44452
rect 20070 44412 20076 44424
rect 20128 44412 20134 44464
rect 20254 44452 20260 44464
rect 20215 44424 20260 44452
rect 20254 44412 20260 44424
rect 20312 44412 20318 44464
rect 20901 44455 20959 44461
rect 20901 44421 20913 44455
rect 20947 44452 20959 44455
rect 21450 44452 21456 44464
rect 20947 44424 21456 44452
rect 20947 44421 20959 44424
rect 20901 44415 20959 44421
rect 21450 44412 21456 44424
rect 21508 44412 21514 44464
rect 21818 44452 21824 44464
rect 21779 44424 21824 44452
rect 21818 44412 21824 44424
rect 21876 44412 21882 44464
rect 22741 44455 22799 44461
rect 22741 44421 22753 44455
rect 22787 44452 22799 44455
rect 23293 44455 23351 44461
rect 23293 44452 23305 44455
rect 22787 44424 23305 44452
rect 22787 44421 22799 44424
rect 22741 44415 22799 44421
rect 23293 44421 23305 44424
rect 23339 44452 23351 44455
rect 23566 44452 23572 44464
rect 23339 44424 23572 44452
rect 23339 44421 23351 44424
rect 23293 44415 23351 44421
rect 23566 44412 23572 44424
rect 23624 44452 23630 44464
rect 23624 44424 25360 44452
rect 23624 44412 23630 44424
rect 15102 44344 15108 44396
rect 15160 44384 15166 44396
rect 15565 44387 15623 44393
rect 15565 44384 15577 44387
rect 15160 44356 15577 44384
rect 15160 44344 15166 44356
rect 15565 44353 15577 44356
rect 15611 44353 15623 44387
rect 15746 44384 15752 44396
rect 15707 44356 15752 44384
rect 15565 44347 15623 44353
rect 15746 44344 15752 44356
rect 15804 44344 15810 44396
rect 16669 44387 16727 44393
rect 16669 44353 16681 44387
rect 16715 44353 16727 44387
rect 16669 44347 16727 44353
rect 16853 44387 16911 44393
rect 16853 44353 16865 44387
rect 16899 44384 16911 44387
rect 16942 44384 16948 44396
rect 16899 44356 16948 44384
rect 16899 44353 16911 44356
rect 16853 44347 16911 44353
rect 16684 44316 16712 44347
rect 16942 44344 16948 44356
rect 17000 44344 17006 44396
rect 17126 44344 17132 44396
rect 17184 44384 17190 44396
rect 17313 44387 17371 44393
rect 17313 44384 17325 44387
rect 17184 44356 17325 44384
rect 17184 44344 17190 44356
rect 17313 44353 17325 44356
rect 17359 44353 17371 44387
rect 17494 44384 17500 44396
rect 17455 44356 17500 44384
rect 17313 44347 17371 44353
rect 17494 44344 17500 44356
rect 17552 44344 17558 44396
rect 18414 44384 18420 44396
rect 18327 44356 18420 44384
rect 18414 44344 18420 44356
rect 18472 44344 18478 44396
rect 18506 44344 18512 44396
rect 18564 44384 18570 44396
rect 21085 44387 21143 44393
rect 18564 44356 18609 44384
rect 18564 44344 18570 44356
rect 21085 44353 21097 44387
rect 21131 44384 21143 44387
rect 21358 44384 21364 44396
rect 21131 44356 21364 44384
rect 21131 44353 21143 44356
rect 21085 44347 21143 44353
rect 21358 44344 21364 44356
rect 21416 44344 21422 44396
rect 22278 44344 22284 44396
rect 22336 44384 22342 44396
rect 22649 44387 22707 44393
rect 22649 44384 22661 44387
rect 22336 44356 22661 44384
rect 22336 44344 22342 44356
rect 22649 44353 22661 44356
rect 22695 44353 22707 44387
rect 22830 44384 22836 44396
rect 22791 44356 22836 44384
rect 22649 44347 22707 44353
rect 22830 44344 22836 44356
rect 22888 44344 22894 44396
rect 23474 44384 23480 44396
rect 23435 44356 23480 44384
rect 23474 44344 23480 44356
rect 23532 44344 23538 44396
rect 23842 44344 23848 44396
rect 23900 44384 23906 44396
rect 25332 44393 25360 44424
rect 25406 44412 25412 44464
rect 25464 44452 25470 44464
rect 25464 44424 26280 44452
rect 25464 44412 25470 44424
rect 24305 44387 24363 44393
rect 24305 44384 24317 44387
rect 23900 44356 24317 44384
rect 23900 44344 23906 44356
rect 24305 44353 24317 44356
rect 24351 44353 24363 44387
rect 24305 44347 24363 44353
rect 25317 44387 25375 44393
rect 25317 44353 25329 44387
rect 25363 44353 25375 44387
rect 25498 44384 25504 44396
rect 25459 44356 25504 44384
rect 25317 44347 25375 44353
rect 25498 44344 25504 44356
rect 25556 44344 25562 44396
rect 25590 44344 25596 44396
rect 25648 44384 25654 44396
rect 26252 44393 26280 44424
rect 27982 44412 27988 44464
rect 28040 44452 28046 44464
rect 28626 44452 28632 44464
rect 28040 44424 28632 44452
rect 28040 44412 28046 44424
rect 28626 44412 28632 44424
rect 28684 44412 28690 44464
rect 30926 44412 30932 44464
rect 30984 44452 30990 44464
rect 31205 44455 31263 44461
rect 31205 44452 31217 44455
rect 30984 44424 31217 44452
rect 30984 44412 30990 44424
rect 31205 44421 31217 44424
rect 31251 44421 31263 44455
rect 31205 44415 31263 44421
rect 32398 44412 32404 44464
rect 32456 44452 32462 44464
rect 34149 44455 34207 44461
rect 32456 44424 33364 44452
rect 32456 44412 32462 44424
rect 26053 44387 26111 44393
rect 25648 44356 25693 44384
rect 25648 44344 25654 44356
rect 26053 44353 26065 44387
rect 26099 44353 26111 44387
rect 26053 44347 26111 44353
rect 26237 44387 26295 44393
rect 26237 44353 26249 44387
rect 26283 44384 26295 44387
rect 26786 44384 26792 44396
rect 26283 44356 26792 44384
rect 26283 44353 26295 44356
rect 26237 44347 26295 44353
rect 18046 44316 18052 44328
rect 15028 44288 18052 44316
rect 15028 44192 15056 44288
rect 18046 44276 18052 44288
rect 18104 44316 18110 44328
rect 18598 44316 18604 44328
rect 18104 44288 18604 44316
rect 18104 44276 18110 44288
rect 18598 44276 18604 44288
rect 18656 44276 18662 44328
rect 18874 44276 18880 44328
rect 18932 44316 18938 44328
rect 22094 44316 22100 44328
rect 18932 44288 22100 44316
rect 18932 44276 18938 44288
rect 22094 44276 22100 44288
rect 22152 44316 22158 44328
rect 22462 44316 22468 44328
rect 22152 44288 22468 44316
rect 22152 44276 22158 44288
rect 22462 44276 22468 44288
rect 22520 44276 22526 44328
rect 24210 44316 24216 44328
rect 24171 44288 24216 44316
rect 24210 44276 24216 44288
rect 24268 44276 24274 44328
rect 24673 44319 24731 44325
rect 24673 44285 24685 44319
rect 24719 44316 24731 44319
rect 26068 44316 26096 44347
rect 26786 44344 26792 44356
rect 26844 44344 26850 44396
rect 27522 44344 27528 44396
rect 27580 44384 27586 44396
rect 27709 44387 27767 44393
rect 27709 44384 27721 44387
rect 27580 44356 27721 44384
rect 27580 44344 27586 44356
rect 27709 44353 27721 44356
rect 27755 44353 27767 44387
rect 30374 44384 30380 44396
rect 30335 44356 30380 44384
rect 27709 44347 27767 44353
rect 30374 44344 30380 44356
rect 30432 44344 30438 44396
rect 31021 44387 31079 44393
rect 31021 44353 31033 44387
rect 31067 44353 31079 44387
rect 31021 44347 31079 44353
rect 24719 44288 26096 44316
rect 27985 44319 28043 44325
rect 24719 44285 24731 44288
rect 24673 44279 24731 44285
rect 27985 44285 27997 44319
rect 28031 44316 28043 44319
rect 28074 44316 28080 44328
rect 28031 44288 28080 44316
rect 28031 44285 28043 44288
rect 27985 44279 28043 44285
rect 28074 44276 28080 44288
rect 28132 44276 28138 44328
rect 15657 44251 15715 44257
rect 15657 44217 15669 44251
rect 15703 44248 15715 44251
rect 17034 44248 17040 44260
rect 15703 44220 17040 44248
rect 15703 44217 15715 44220
rect 15657 44211 15715 44217
rect 17034 44208 17040 44220
rect 17092 44208 17098 44260
rect 18690 44248 18696 44260
rect 18651 44220 18696 44248
rect 18690 44208 18696 44220
rect 18748 44208 18754 44260
rect 19521 44251 19579 44257
rect 19521 44217 19533 44251
rect 19567 44248 19579 44251
rect 21174 44248 21180 44260
rect 19567 44220 21180 44248
rect 19567 44217 19579 44220
rect 19521 44211 19579 44217
rect 21174 44208 21180 44220
rect 21232 44208 21238 44260
rect 22189 44251 22247 44257
rect 22189 44217 22201 44251
rect 22235 44248 22247 44251
rect 26142 44248 26148 44260
rect 22235 44220 26148 44248
rect 22235 44217 22247 44220
rect 22189 44211 22247 44217
rect 26142 44208 26148 44220
rect 26200 44208 26206 44260
rect 27893 44251 27951 44257
rect 27893 44217 27905 44251
rect 27939 44248 27951 44251
rect 31036 44248 31064 44347
rect 31294 44344 31300 44396
rect 31352 44384 31358 44396
rect 32125 44387 32183 44393
rect 31352 44356 31397 44384
rect 31352 44344 31358 44356
rect 32125 44353 32137 44387
rect 32171 44353 32183 44387
rect 32306 44384 32312 44396
rect 32267 44356 32312 44384
rect 32125 44347 32183 44353
rect 27939 44220 31064 44248
rect 32140 44248 32168 44347
rect 32306 44344 32312 44356
rect 32364 44344 32370 44396
rect 32582 44344 32588 44396
rect 32640 44384 32646 44396
rect 32769 44387 32827 44393
rect 32769 44384 32781 44387
rect 32640 44356 32781 44384
rect 32640 44344 32646 44356
rect 32769 44353 32781 44356
rect 32815 44353 32827 44387
rect 32769 44347 32827 44353
rect 32953 44387 33011 44393
rect 32953 44353 32965 44387
rect 32999 44353 33011 44387
rect 32953 44347 33011 44353
rect 32217 44319 32275 44325
rect 32217 44285 32229 44319
rect 32263 44316 32275 44319
rect 32968 44316 32996 44347
rect 33042 44344 33048 44396
rect 33100 44384 33106 44396
rect 33336 44393 33364 44424
rect 34149 44421 34161 44455
rect 34195 44452 34207 44455
rect 34900 44452 34928 44480
rect 34195 44424 34928 44452
rect 34195 44421 34207 44424
rect 34149 44415 34207 44421
rect 33321 44387 33379 44393
rect 33100 44356 33145 44384
rect 33100 44344 33106 44356
rect 33321 44353 33333 44387
rect 33367 44353 33379 44387
rect 33321 44347 33379 44353
rect 32263 44288 32996 44316
rect 32263 44285 32275 44288
rect 32217 44279 32275 44285
rect 33134 44276 33140 44328
rect 33192 44316 33198 44328
rect 33336 44316 33364 44347
rect 34422 44344 34428 44396
rect 34480 44384 34486 44396
rect 35529 44387 35587 44393
rect 34480 44356 34525 44384
rect 34480 44344 34486 44356
rect 35529 44353 35541 44387
rect 35575 44384 35587 44387
rect 36188 44384 36216 44480
rect 35575 44356 36216 44384
rect 35575 44353 35587 44356
rect 35529 44347 35587 44353
rect 36262 44344 36268 44396
rect 36320 44384 36326 44396
rect 36357 44387 36415 44393
rect 36357 44384 36369 44387
rect 36320 44356 36369 44384
rect 36320 44344 36326 44356
rect 36357 44353 36369 44356
rect 36403 44353 36415 44387
rect 36538 44384 36544 44396
rect 36499 44356 36544 44384
rect 36357 44347 36415 44353
rect 36538 44344 36544 44356
rect 36596 44344 36602 44396
rect 35710 44316 35716 44328
rect 33192 44288 33237 44316
rect 33336 44288 34284 44316
rect 35671 44288 35716 44316
rect 33192 44276 33198 44288
rect 32950 44248 32956 44260
rect 32140 44220 32956 44248
rect 27939 44217 27951 44220
rect 27893 44211 27951 44217
rect 32950 44208 32956 44220
rect 33008 44248 33014 44260
rect 33410 44248 33416 44260
rect 33008 44220 33416 44248
rect 33008 44208 33014 44220
rect 33410 44208 33416 44220
rect 33468 44208 33474 44260
rect 34146 44248 34152 44260
rect 34107 44220 34152 44248
rect 34146 44208 34152 44220
rect 34204 44208 34210 44260
rect 34256 44248 34284 44288
rect 35710 44276 35716 44288
rect 35768 44276 35774 44328
rect 34256 44220 34928 44248
rect 1670 44140 1676 44192
rect 1728 44180 1734 44192
rect 13725 44183 13783 44189
rect 13725 44180 13737 44183
rect 1728 44152 13737 44180
rect 1728 44140 1734 44152
rect 13725 44149 13737 44152
rect 13771 44180 13783 44183
rect 14090 44180 14096 44192
rect 13771 44152 14096 44180
rect 13771 44149 13783 44152
rect 13725 44143 13783 44149
rect 14090 44140 14096 44152
rect 14148 44140 14154 44192
rect 14458 44180 14464 44192
rect 14419 44152 14464 44180
rect 14458 44140 14464 44152
rect 14516 44140 14522 44192
rect 15010 44180 15016 44192
rect 14971 44152 15016 44180
rect 15010 44140 15016 44152
rect 15068 44140 15074 44192
rect 16853 44183 16911 44189
rect 16853 44149 16865 44183
rect 16899 44180 16911 44183
rect 17126 44180 17132 44192
rect 16899 44152 17132 44180
rect 16899 44149 16911 44152
rect 16853 44143 16911 44149
rect 17126 44140 17132 44152
rect 17184 44140 17190 44192
rect 17678 44180 17684 44192
rect 17639 44152 17684 44180
rect 17678 44140 17684 44152
rect 17736 44140 17742 44192
rect 18506 44140 18512 44192
rect 18564 44180 18570 44192
rect 19337 44183 19395 44189
rect 19337 44180 19349 44183
rect 18564 44152 19349 44180
rect 18564 44140 18570 44152
rect 19337 44149 19349 44152
rect 19383 44149 19395 44183
rect 19337 44143 19395 44149
rect 20441 44183 20499 44189
rect 20441 44149 20453 44183
rect 20487 44180 20499 44183
rect 20806 44180 20812 44192
rect 20487 44152 20812 44180
rect 20487 44149 20499 44152
rect 20441 44143 20499 44149
rect 20806 44140 20812 44152
rect 20864 44140 20870 44192
rect 21269 44183 21327 44189
rect 21269 44149 21281 44183
rect 21315 44180 21327 44183
rect 22005 44183 22063 44189
rect 22005 44180 22017 44183
rect 21315 44152 22017 44180
rect 21315 44149 21327 44152
rect 21269 44143 21327 44149
rect 22005 44149 22017 44152
rect 22051 44149 22063 44183
rect 22005 44143 22063 44149
rect 23661 44183 23719 44189
rect 23661 44149 23673 44183
rect 23707 44180 23719 44183
rect 25038 44180 25044 44192
rect 23707 44152 25044 44180
rect 23707 44149 23719 44152
rect 23661 44143 23719 44149
rect 25038 44140 25044 44152
rect 25096 44140 25102 44192
rect 26234 44140 26240 44192
rect 26292 44180 26298 44192
rect 27157 44183 27215 44189
rect 27157 44180 27169 44183
rect 26292 44152 27169 44180
rect 26292 44140 26298 44152
rect 27157 44149 27169 44152
rect 27203 44149 27215 44183
rect 27157 44143 27215 44149
rect 27801 44183 27859 44189
rect 27801 44149 27813 44183
rect 27847 44180 27859 44183
rect 31294 44180 31300 44192
rect 27847 44152 31300 44180
rect 27847 44149 27859 44152
rect 27801 44143 27859 44149
rect 31294 44140 31300 44152
rect 31352 44140 31358 44192
rect 31570 44140 31576 44192
rect 31628 44180 31634 44192
rect 34790 44180 34796 44192
rect 31628 44152 34796 44180
rect 31628 44140 31634 44152
rect 34790 44140 34796 44152
rect 34848 44140 34854 44192
rect 34900 44180 34928 44220
rect 36722 44208 36728 44260
rect 36780 44248 36786 44260
rect 38378 44248 38384 44260
rect 36780 44220 38384 44248
rect 36780 44208 36786 44220
rect 38378 44208 38384 44220
rect 38436 44208 38442 44260
rect 35710 44180 35716 44192
rect 34900 44152 35716 44180
rect 35710 44140 35716 44152
rect 35768 44180 35774 44192
rect 37829 44183 37887 44189
rect 37829 44180 37841 44183
rect 35768 44152 37841 44180
rect 35768 44140 35774 44152
rect 37829 44149 37841 44152
rect 37875 44149 37887 44183
rect 37829 44143 37887 44149
rect 39025 44183 39083 44189
rect 39025 44149 39037 44183
rect 39071 44180 39083 44183
rect 39114 44180 39120 44192
rect 39071 44152 39120 44180
rect 39071 44149 39083 44152
rect 39025 44143 39083 44149
rect 39114 44140 39120 44152
rect 39172 44140 39178 44192
rect 1104 44090 54372 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 54372 44090
rect 1104 44016 54372 44038
rect 10686 43936 10692 43988
rect 10744 43976 10750 43988
rect 13449 43979 13507 43985
rect 13449 43976 13461 43979
rect 10744 43948 13461 43976
rect 10744 43936 10750 43948
rect 13449 43945 13461 43948
rect 13495 43976 13507 43979
rect 15286 43976 15292 43988
rect 13495 43948 15292 43976
rect 13495 43945 13507 43948
rect 13449 43939 13507 43945
rect 15286 43936 15292 43948
rect 15344 43936 15350 43988
rect 17405 43979 17463 43985
rect 17405 43945 17417 43979
rect 17451 43976 17463 43979
rect 18414 43976 18420 43988
rect 17451 43948 18276 43976
rect 18375 43948 18420 43976
rect 17451 43945 17463 43948
rect 17405 43939 17463 43945
rect 15657 43911 15715 43917
rect 15657 43877 15669 43911
rect 15703 43908 15715 43911
rect 16850 43908 16856 43920
rect 15703 43880 16856 43908
rect 15703 43877 15715 43880
rect 15657 43871 15715 43877
rect 16850 43868 16856 43880
rect 16908 43868 16914 43920
rect 17494 43908 17500 43920
rect 16960 43880 17500 43908
rect 2746 43812 9674 43840
rect 2041 43775 2099 43781
rect 2041 43741 2053 43775
rect 2087 43772 2099 43775
rect 2746 43772 2774 43812
rect 2087 43744 2774 43772
rect 2087 43741 2099 43744
rect 2041 43735 2099 43741
rect 1578 43664 1584 43716
rect 1636 43704 1642 43716
rect 1857 43707 1915 43713
rect 1857 43704 1869 43707
rect 1636 43676 1869 43704
rect 1636 43664 1642 43676
rect 1857 43673 1869 43676
rect 1903 43673 1915 43707
rect 1857 43667 1915 43673
rect 9646 43636 9674 43812
rect 14458 43800 14464 43852
rect 14516 43840 14522 43852
rect 16298 43840 16304 43852
rect 14516 43812 16304 43840
rect 14516 43800 14522 43812
rect 14734 43772 14740 43784
rect 14695 43744 14740 43772
rect 14734 43732 14740 43744
rect 14792 43732 14798 43784
rect 14918 43772 14924 43784
rect 14879 43744 14924 43772
rect 14918 43732 14924 43744
rect 14976 43732 14982 43784
rect 15286 43732 15292 43784
rect 15344 43772 15350 43784
rect 15488 43781 15516 43812
rect 16298 43800 16304 43812
rect 16356 43800 16362 43852
rect 15381 43775 15439 43781
rect 15381 43772 15393 43775
rect 15344 43744 15393 43772
rect 15344 43732 15350 43744
rect 15381 43741 15393 43744
rect 15427 43741 15439 43775
rect 15381 43735 15439 43741
rect 15473 43775 15531 43781
rect 15473 43741 15485 43775
rect 15519 43741 15531 43775
rect 15473 43735 15531 43741
rect 15657 43775 15715 43781
rect 15657 43741 15669 43775
rect 15703 43772 15715 43775
rect 16960 43772 16988 43880
rect 17494 43868 17500 43880
rect 17552 43868 17558 43920
rect 18248 43908 18276 43948
rect 18414 43936 18420 43948
rect 18472 43936 18478 43988
rect 18598 43936 18604 43988
rect 18656 43976 18662 43988
rect 18656 43948 20852 43976
rect 18656 43936 18662 43948
rect 19978 43908 19984 43920
rect 18248 43880 19984 43908
rect 19978 43868 19984 43880
rect 20036 43868 20042 43920
rect 20346 43868 20352 43920
rect 20404 43908 20410 43920
rect 20441 43911 20499 43917
rect 20441 43908 20453 43911
rect 20404 43880 20453 43908
rect 20404 43868 20410 43880
rect 20441 43877 20453 43880
rect 20487 43877 20499 43911
rect 20824 43908 20852 43948
rect 20898 43936 20904 43988
rect 20956 43976 20962 43988
rect 21177 43979 21235 43985
rect 21177 43976 21189 43979
rect 20956 43948 21189 43976
rect 20956 43936 20962 43948
rect 21177 43945 21189 43948
rect 21223 43945 21235 43979
rect 21177 43939 21235 43945
rect 23750 43936 23756 43988
rect 23808 43976 23814 43988
rect 23845 43979 23903 43985
rect 23845 43976 23857 43979
rect 23808 43948 23857 43976
rect 23808 43936 23814 43948
rect 23845 43945 23857 43948
rect 23891 43976 23903 43979
rect 24578 43976 24584 43988
rect 23891 43948 24584 43976
rect 23891 43945 23903 43948
rect 23845 43939 23903 43945
rect 24578 43936 24584 43948
rect 24636 43936 24642 43988
rect 25133 43979 25191 43985
rect 25133 43945 25145 43979
rect 25179 43976 25191 43979
rect 25682 43976 25688 43988
rect 25179 43948 25688 43976
rect 25179 43945 25191 43948
rect 25133 43939 25191 43945
rect 25682 43936 25688 43948
rect 25740 43936 25746 43988
rect 28353 43979 28411 43985
rect 28353 43976 28365 43979
rect 26068 43948 28365 43976
rect 22005 43911 22063 43917
rect 20824 43880 21956 43908
rect 20441 43871 20499 43877
rect 17218 43840 17224 43852
rect 17179 43812 17224 43840
rect 17218 43800 17224 43812
rect 17276 43800 17282 43852
rect 17678 43800 17684 43852
rect 17736 43840 17742 43852
rect 21928 43840 21956 43880
rect 22005 43877 22017 43911
rect 22051 43908 22063 43911
rect 23934 43908 23940 43920
rect 22051 43880 23940 43908
rect 22051 43877 22063 43880
rect 22005 43871 22063 43877
rect 23934 43868 23940 43880
rect 23992 43868 23998 43920
rect 26068 43908 26096 43948
rect 28353 43945 28365 43948
rect 28399 43976 28411 43979
rect 28994 43976 29000 43988
rect 28399 43948 29000 43976
rect 28399 43945 28411 43948
rect 28353 43939 28411 43945
rect 28994 43936 29000 43948
rect 29052 43936 29058 43988
rect 32766 43936 32772 43988
rect 32824 43976 32830 43988
rect 32861 43979 32919 43985
rect 32861 43976 32873 43979
rect 32824 43948 32873 43976
rect 32824 43936 32830 43948
rect 32861 43945 32873 43948
rect 32907 43945 32919 43979
rect 33410 43976 33416 43988
rect 33371 43948 33416 43976
rect 32861 43939 32919 43945
rect 25148 43880 26096 43908
rect 22278 43840 22284 43852
rect 17736 43812 18276 43840
rect 21928 43812 22284 43840
rect 17736 43800 17742 43812
rect 15703 43744 16988 43772
rect 15703 43741 15715 43744
rect 15657 43735 15715 43741
rect 15396 43704 15424 43735
rect 17034 43732 17040 43784
rect 17092 43772 17098 43784
rect 17129 43775 17187 43781
rect 17129 43772 17141 43775
rect 17092 43744 17141 43772
rect 17092 43732 17098 43744
rect 17129 43741 17141 43744
rect 17175 43741 17187 43775
rect 17129 43735 17187 43741
rect 17586 43732 17592 43784
rect 17644 43772 17650 43784
rect 18248 43781 18276 43812
rect 22278 43800 22284 43812
rect 22336 43840 22342 43852
rect 22557 43843 22615 43849
rect 22557 43840 22569 43843
rect 22336 43812 22569 43840
rect 22336 43800 22342 43812
rect 22557 43809 22569 43812
rect 22603 43809 22615 43843
rect 23753 43843 23811 43849
rect 22557 43803 22615 43809
rect 22848 43812 23704 43840
rect 22848 43784 22876 43812
rect 17957 43775 18015 43781
rect 17957 43772 17969 43775
rect 17644 43744 17969 43772
rect 17644 43732 17650 43744
rect 17957 43741 17969 43744
rect 18003 43772 18015 43775
rect 18233 43775 18291 43781
rect 18003 43744 18184 43772
rect 18003 43741 18015 43744
rect 17957 43735 18015 43741
rect 16117 43707 16175 43713
rect 16117 43704 16129 43707
rect 15396 43676 16129 43704
rect 16117 43673 16129 43676
rect 16163 43673 16175 43707
rect 16298 43704 16304 43716
rect 16259 43676 16304 43704
rect 16117 43667 16175 43673
rect 16298 43664 16304 43676
rect 16356 43664 16362 43716
rect 17862 43664 17868 43716
rect 17920 43704 17926 43716
rect 18049 43707 18107 43713
rect 18049 43704 18061 43707
rect 17920 43676 18061 43704
rect 17920 43664 17926 43676
rect 18049 43673 18061 43676
rect 18095 43673 18107 43707
rect 18156 43704 18184 43744
rect 18233 43741 18245 43775
rect 18279 43741 18291 43775
rect 18233 43735 18291 43741
rect 19426 43732 19432 43784
rect 19484 43772 19490 43784
rect 19521 43775 19579 43781
rect 19521 43772 19533 43775
rect 19484 43744 19533 43772
rect 19484 43732 19490 43744
rect 19521 43741 19533 43744
rect 19567 43741 19579 43775
rect 19521 43735 19579 43741
rect 20070 43732 20076 43784
rect 20128 43772 20134 43784
rect 20441 43775 20499 43781
rect 20441 43772 20453 43775
rect 20128 43744 20453 43772
rect 20128 43732 20134 43744
rect 20441 43741 20453 43744
rect 20487 43741 20499 43775
rect 20714 43772 20720 43784
rect 20675 43744 20720 43772
rect 20441 43735 20499 43741
rect 20714 43732 20720 43744
rect 20772 43732 20778 43784
rect 21174 43772 21180 43784
rect 21135 43744 21180 43772
rect 21174 43732 21180 43744
rect 21232 43732 21238 43784
rect 21450 43772 21456 43784
rect 21411 43744 21456 43772
rect 21450 43732 21456 43744
rect 21508 43732 21514 43784
rect 21913 43775 21971 43781
rect 21913 43741 21925 43775
rect 21959 43772 21971 43775
rect 22002 43772 22008 43784
rect 21959 43744 22008 43772
rect 21959 43741 21971 43744
rect 21913 43735 21971 43741
rect 22002 43732 22008 43744
rect 22060 43732 22066 43784
rect 22094 43732 22100 43784
rect 22152 43772 22158 43784
rect 22741 43775 22799 43781
rect 22152 43744 22197 43772
rect 22152 43732 22158 43744
rect 22741 43741 22753 43775
rect 22787 43772 22799 43775
rect 22830 43772 22836 43784
rect 22787 43744 22836 43772
rect 22787 43741 22799 43744
rect 22741 43735 22799 43741
rect 22830 43732 22836 43744
rect 22888 43732 22894 43784
rect 23566 43772 23572 43784
rect 23527 43744 23572 43772
rect 23566 43732 23572 43744
rect 23624 43732 23630 43784
rect 23676 43772 23704 43812
rect 23753 43809 23765 43843
rect 23799 43840 23811 43843
rect 24026 43840 24032 43852
rect 23799 43812 24032 43840
rect 23799 43809 23811 43812
rect 23753 43803 23811 43809
rect 24026 43800 24032 43812
rect 24084 43800 24090 43852
rect 25038 43840 25044 43852
rect 24999 43812 25044 43840
rect 25038 43800 25044 43812
rect 25096 43800 25102 43852
rect 25148 43772 25176 43880
rect 26142 43868 26148 43920
rect 26200 43908 26206 43920
rect 26237 43911 26295 43917
rect 26237 43908 26249 43911
rect 26200 43880 26249 43908
rect 26200 43868 26206 43880
rect 26237 43877 26249 43880
rect 26283 43877 26295 43911
rect 26237 43871 26295 43877
rect 25501 43843 25559 43849
rect 25501 43809 25513 43843
rect 25547 43840 25559 43843
rect 26973 43843 27031 43849
rect 25547 43812 26372 43840
rect 25547 43809 25559 43812
rect 25501 43803 25559 43809
rect 25314 43772 25320 43784
rect 23676 43744 25176 43772
rect 25275 43744 25320 43772
rect 25314 43732 25320 43744
rect 25372 43732 25378 43784
rect 25774 43732 25780 43784
rect 25832 43772 25838 43784
rect 26344 43781 26372 43812
rect 26973 43809 26985 43843
rect 27019 43840 27031 43843
rect 28626 43840 28632 43852
rect 27019 43812 28632 43840
rect 27019 43809 27031 43812
rect 26973 43803 27031 43809
rect 28626 43800 28632 43812
rect 28684 43840 28690 43852
rect 29549 43843 29607 43849
rect 29549 43840 29561 43843
rect 28684 43812 29561 43840
rect 28684 43800 28690 43812
rect 29549 43809 29561 43812
rect 29595 43809 29607 43843
rect 32876 43840 32904 43939
rect 33410 43936 33416 43948
rect 33468 43936 33474 43988
rect 34790 43936 34796 43988
rect 34848 43976 34854 43988
rect 35253 43979 35311 43985
rect 35253 43976 35265 43979
rect 34848 43948 35265 43976
rect 34848 43936 34854 43948
rect 35253 43945 35265 43948
rect 35299 43945 35311 43979
rect 35253 43939 35311 43945
rect 36357 43979 36415 43985
rect 36357 43945 36369 43979
rect 36403 43976 36415 43979
rect 36538 43976 36544 43988
rect 36403 43948 36544 43976
rect 36403 43945 36415 43948
rect 36357 43939 36415 43945
rect 36538 43936 36544 43948
rect 36596 43936 36602 43988
rect 36262 43908 36268 43920
rect 34808 43880 36268 43908
rect 34808 43852 34836 43880
rect 36262 43868 36268 43880
rect 36320 43908 36326 43920
rect 37826 43908 37832 43920
rect 36320 43880 37832 43908
rect 36320 43868 36326 43880
rect 37826 43868 37832 43880
rect 37884 43908 37890 43920
rect 37921 43911 37979 43917
rect 37921 43908 37933 43911
rect 37884 43880 37933 43908
rect 37884 43868 37890 43880
rect 37921 43877 37933 43880
rect 37967 43877 37979 43911
rect 37921 43871 37979 43877
rect 33042 43840 33048 43852
rect 32876 43812 33048 43840
rect 29549 43803 29607 43809
rect 33042 43800 33048 43812
rect 33100 43840 33106 43852
rect 33781 43843 33839 43849
rect 33781 43840 33793 43843
rect 33100 43812 33793 43840
rect 33100 43800 33106 43812
rect 33781 43809 33793 43812
rect 33827 43840 33839 43843
rect 34790 43840 34796 43852
rect 33827 43812 34796 43840
rect 33827 43809 33839 43812
rect 33781 43803 33839 43809
rect 34790 43800 34796 43812
rect 34848 43800 34854 43852
rect 35894 43840 35900 43852
rect 35855 43812 35900 43840
rect 35894 43800 35900 43812
rect 35952 43800 35958 43852
rect 26053 43775 26111 43781
rect 26053 43772 26065 43775
rect 25832 43744 26065 43772
rect 25832 43732 25838 43744
rect 26053 43741 26065 43744
rect 26099 43741 26111 43775
rect 26053 43735 26111 43741
rect 26145 43775 26203 43781
rect 26145 43741 26157 43775
rect 26191 43741 26203 43775
rect 26145 43735 26203 43741
rect 26329 43775 26387 43781
rect 26329 43741 26341 43775
rect 26375 43741 26387 43775
rect 26329 43735 26387 43741
rect 26513 43775 26571 43781
rect 26513 43741 26525 43775
rect 26559 43772 26571 43775
rect 27249 43775 27307 43781
rect 27249 43772 27261 43775
rect 26559 43744 27261 43772
rect 26559 43741 26571 43744
rect 26513 43735 26571 43741
rect 27249 43741 27261 43744
rect 27295 43741 27307 43775
rect 27249 43735 27307 43741
rect 18598 43704 18604 43716
rect 18156 43676 18604 43704
rect 18049 43667 18107 43673
rect 18598 43664 18604 43676
rect 18656 43664 18662 43716
rect 19613 43707 19671 43713
rect 19613 43673 19625 43707
rect 19659 43673 19671 43707
rect 19613 43667 19671 43673
rect 19797 43707 19855 43713
rect 19797 43673 19809 43707
rect 19843 43704 19855 43707
rect 19978 43704 19984 43716
rect 19843 43676 19984 43704
rect 19843 43673 19855 43676
rect 19797 43667 19855 43673
rect 14185 43639 14243 43645
rect 14185 43636 14197 43639
rect 9646 43608 14197 43636
rect 14185 43605 14197 43608
rect 14231 43636 14243 43639
rect 14458 43636 14464 43648
rect 14231 43608 14464 43636
rect 14231 43605 14243 43608
rect 14185 43599 14243 43605
rect 14458 43596 14464 43608
rect 14516 43596 14522 43648
rect 14921 43639 14979 43645
rect 14921 43605 14933 43639
rect 14967 43636 14979 43639
rect 15378 43636 15384 43648
rect 14967 43608 15384 43636
rect 14967 43605 14979 43608
rect 14921 43599 14979 43605
rect 15378 43596 15384 43608
rect 15436 43596 15442 43648
rect 16485 43639 16543 43645
rect 16485 43605 16497 43639
rect 16531 43636 16543 43639
rect 17402 43636 17408 43648
rect 16531 43608 17408 43636
rect 16531 43605 16543 43608
rect 16485 43599 16543 43605
rect 17402 43596 17408 43608
rect 17460 43596 17466 43648
rect 17770 43596 17776 43648
rect 17828 43636 17834 43648
rect 19334 43636 19340 43648
rect 17828 43608 19340 43636
rect 17828 43596 17834 43608
rect 19334 43596 19340 43608
rect 19392 43636 19398 43648
rect 19628 43636 19656 43667
rect 19978 43664 19984 43676
rect 20036 43664 20042 43716
rect 20625 43707 20683 43713
rect 20625 43673 20637 43707
rect 20671 43704 20683 43707
rect 21082 43704 21088 43716
rect 20671 43676 21088 43704
rect 20671 43673 20683 43676
rect 20625 43667 20683 43673
rect 21082 43664 21088 43676
rect 21140 43664 21146 43716
rect 22925 43707 22983 43713
rect 22925 43673 22937 43707
rect 22971 43704 22983 43707
rect 23474 43704 23480 43716
rect 22971 43676 23480 43704
rect 22971 43673 22983 43676
rect 22925 43667 22983 43673
rect 23474 43664 23480 43676
rect 23532 43664 23538 43716
rect 23842 43704 23848 43716
rect 23803 43676 23848 43704
rect 23842 43664 23848 43676
rect 23900 43664 23906 43716
rect 24026 43664 24032 43716
rect 24084 43704 24090 43716
rect 25590 43704 25596 43716
rect 24084 43676 25596 43704
rect 24084 43664 24090 43676
rect 25590 43664 25596 43676
rect 25648 43664 25654 43716
rect 19392 43608 19656 43636
rect 19705 43639 19763 43645
rect 19392 43596 19398 43608
rect 19705 43605 19717 43639
rect 19751 43636 19763 43639
rect 20070 43636 20076 43648
rect 19751 43608 20076 43636
rect 19751 43605 19763 43608
rect 19705 43599 19763 43605
rect 20070 43596 20076 43608
rect 20128 43596 20134 43648
rect 21358 43636 21364 43648
rect 21319 43608 21364 43636
rect 21358 43596 21364 43608
rect 21416 43596 21422 43648
rect 23385 43639 23443 43645
rect 23385 43605 23397 43639
rect 23431 43636 23443 43639
rect 23566 43636 23572 43648
rect 23431 43608 23572 43636
rect 23431 43605 23443 43608
rect 23385 43599 23443 43605
rect 23566 43596 23572 43608
rect 23624 43596 23630 43648
rect 24394 43636 24400 43648
rect 24355 43608 24400 43636
rect 24394 43596 24400 43608
rect 24452 43596 24458 43648
rect 26160 43636 26188 43735
rect 28902 43732 28908 43784
rect 28960 43772 28966 43784
rect 29805 43775 29863 43781
rect 29805 43772 29817 43775
rect 28960 43744 29817 43772
rect 28960 43732 28966 43744
rect 29805 43741 29817 43744
rect 29851 43741 29863 43775
rect 29805 43735 29863 43741
rect 30098 43732 30104 43784
rect 30156 43772 30162 43784
rect 30926 43772 30932 43784
rect 30156 43744 30932 43772
rect 30156 43732 30162 43744
rect 30926 43732 30932 43744
rect 30984 43772 30990 43784
rect 31481 43775 31539 43781
rect 31481 43772 31493 43775
rect 30984 43744 31493 43772
rect 30984 43732 30990 43744
rect 31481 43741 31493 43744
rect 31527 43741 31539 43775
rect 31481 43735 31539 43741
rect 31748 43775 31806 43781
rect 31748 43741 31760 43775
rect 31794 43772 31806 43775
rect 33226 43772 33232 43784
rect 31794 43744 33232 43772
rect 31794 43741 31806 43744
rect 31748 43735 31806 43741
rect 33226 43732 33232 43744
rect 33284 43732 33290 43784
rect 33594 43772 33600 43784
rect 33555 43744 33600 43772
rect 33594 43732 33600 43744
rect 33652 43732 33658 43784
rect 35989 43775 36047 43781
rect 35989 43741 36001 43775
rect 36035 43772 36047 43775
rect 36262 43772 36268 43784
rect 36035 43744 36268 43772
rect 36035 43741 36047 43744
rect 35989 43735 36047 43741
rect 36262 43732 36268 43744
rect 36320 43772 36326 43784
rect 36446 43772 36452 43784
rect 36320 43744 36452 43772
rect 36320 43732 36326 43744
rect 36446 43732 36452 43744
rect 36504 43732 36510 43784
rect 53377 43775 53435 43781
rect 53377 43772 53389 43775
rect 52840 43744 53389 43772
rect 32674 43704 32680 43716
rect 30944 43676 32680 43704
rect 28258 43636 28264 43648
rect 26160 43608 28264 43636
rect 28258 43596 28264 43608
rect 28316 43596 28322 43648
rect 30742 43596 30748 43648
rect 30800 43636 30806 43648
rect 30944 43645 30972 43676
rect 32674 43664 32680 43676
rect 32732 43664 32738 43716
rect 34701 43707 34759 43713
rect 34701 43704 34713 43707
rect 32784 43676 34713 43704
rect 30929 43639 30987 43645
rect 30929 43636 30941 43639
rect 30800 43608 30941 43636
rect 30800 43596 30806 43608
rect 30929 43605 30941 43608
rect 30975 43605 30987 43639
rect 30929 43599 30987 43605
rect 31478 43596 31484 43648
rect 31536 43636 31542 43648
rect 32784 43636 32812 43676
rect 34701 43673 34713 43676
rect 34747 43673 34759 43707
rect 34701 43667 34759 43673
rect 37461 43707 37519 43713
rect 37461 43673 37473 43707
rect 37507 43704 37519 43707
rect 37507 43676 39160 43704
rect 37507 43673 37519 43676
rect 37461 43667 37519 43673
rect 39132 43648 39160 43676
rect 31536 43608 32812 43636
rect 31536 43596 31542 43608
rect 36722 43596 36728 43648
rect 36780 43636 36786 43648
rect 36817 43639 36875 43645
rect 36817 43636 36829 43639
rect 36780 43608 36829 43636
rect 36780 43596 36786 43608
rect 36817 43605 36829 43608
rect 36863 43605 36875 43639
rect 36817 43599 36875 43605
rect 38565 43639 38623 43645
rect 38565 43605 38577 43639
rect 38611 43636 38623 43639
rect 38654 43636 38660 43648
rect 38611 43608 38660 43636
rect 38611 43605 38623 43608
rect 38565 43599 38623 43605
rect 38654 43596 38660 43608
rect 38712 43596 38718 43648
rect 39114 43636 39120 43648
rect 39075 43608 39120 43636
rect 39114 43596 39120 43608
rect 39172 43596 39178 43648
rect 52362 43596 52368 43648
rect 52420 43636 52426 43648
rect 52840 43645 52868 43744
rect 53377 43741 53389 43744
rect 53423 43741 53435 43775
rect 53377 43735 53435 43741
rect 52825 43639 52883 43645
rect 52825 43636 52837 43639
rect 52420 43608 52837 43636
rect 52420 43596 52426 43608
rect 52825 43605 52837 43608
rect 52871 43605 52883 43639
rect 53558 43636 53564 43648
rect 53519 43608 53564 43636
rect 52825 43599 52883 43605
rect 53558 43596 53564 43608
rect 53616 43596 53622 43648
rect 1104 43546 54372 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 54372 43546
rect 1104 43472 54372 43494
rect 1578 43432 1584 43444
rect 1539 43404 1584 43432
rect 1578 43392 1584 43404
rect 1636 43392 1642 43444
rect 14461 43435 14519 43441
rect 14461 43401 14473 43435
rect 14507 43432 14519 43435
rect 14918 43432 14924 43444
rect 14507 43404 14924 43432
rect 14507 43401 14519 43404
rect 14461 43395 14519 43401
rect 14918 43392 14924 43404
rect 14976 43392 14982 43444
rect 16942 43392 16948 43444
rect 17000 43432 17006 43444
rect 17586 43432 17592 43444
rect 17000 43404 17592 43432
rect 17000 43392 17006 43404
rect 17586 43392 17592 43404
rect 17644 43392 17650 43444
rect 18506 43432 18512 43444
rect 18467 43404 18512 43432
rect 18506 43392 18512 43404
rect 18564 43392 18570 43444
rect 19334 43392 19340 43444
rect 19392 43432 19398 43444
rect 19521 43435 19579 43441
rect 19521 43432 19533 43435
rect 19392 43404 19533 43432
rect 19392 43392 19398 43404
rect 19521 43401 19533 43404
rect 19567 43401 19579 43435
rect 23198 43432 23204 43444
rect 19521 43395 19579 43401
rect 21928 43404 23204 43432
rect 14090 43364 14096 43376
rect 14051 43336 14096 43364
rect 14090 43324 14096 43336
rect 14148 43324 14154 43376
rect 13081 43299 13139 43305
rect 13081 43265 13093 43299
rect 13127 43296 13139 43299
rect 13633 43299 13691 43305
rect 13633 43296 13645 43299
rect 13127 43268 13645 43296
rect 13127 43265 13139 43268
rect 13081 43259 13139 43265
rect 13633 43265 13645 43268
rect 13679 43296 13691 43299
rect 14274 43296 14280 43308
rect 13679 43268 14280 43296
rect 13679 43265 13691 43268
rect 13633 43259 13691 43265
rect 14274 43256 14280 43268
rect 14332 43256 14338 43308
rect 14734 43256 14740 43308
rect 14792 43296 14798 43308
rect 15381 43299 15439 43305
rect 15381 43296 15393 43299
rect 14792 43268 15393 43296
rect 14792 43256 14798 43268
rect 15381 43265 15393 43268
rect 15427 43265 15439 43299
rect 16850 43296 16856 43308
rect 16811 43268 16856 43296
rect 15381 43259 15439 43265
rect 16850 43256 16856 43268
rect 16908 43256 16914 43308
rect 16960 43305 16988 43392
rect 17310 43324 17316 43376
rect 17368 43364 17374 43376
rect 17368 43336 17632 43364
rect 17368 43324 17374 43336
rect 16945 43299 17003 43305
rect 16945 43265 16957 43299
rect 16991 43265 17003 43299
rect 16945 43259 17003 43265
rect 17034 43256 17040 43308
rect 17092 43296 17098 43308
rect 17129 43299 17187 43305
rect 17129 43296 17141 43299
rect 17092 43268 17141 43296
rect 17092 43256 17098 43268
rect 17129 43265 17141 43268
rect 17175 43265 17187 43299
rect 17129 43259 17187 43265
rect 17218 43256 17224 43308
rect 17276 43296 17282 43308
rect 17604 43296 17632 43336
rect 17678 43324 17684 43376
rect 17736 43364 17742 43376
rect 18785 43367 18843 43373
rect 18785 43364 18797 43367
rect 17736 43336 18797 43364
rect 17736 43324 17742 43336
rect 18785 43333 18797 43336
rect 18831 43333 18843 43367
rect 19978 43364 19984 43376
rect 18785 43327 18843 43333
rect 19444 43336 19984 43364
rect 17865 43299 17923 43305
rect 17865 43296 17877 43299
rect 17276 43268 17321 43296
rect 17604 43268 17877 43296
rect 17276 43256 17282 43268
rect 17865 43265 17877 43268
rect 17911 43265 17923 43299
rect 17865 43259 17923 43265
rect 17954 43256 17960 43308
rect 18012 43296 18018 43308
rect 18509 43299 18567 43305
rect 18509 43296 18521 43299
rect 18012 43268 18521 43296
rect 18012 43256 18018 43268
rect 18509 43265 18521 43268
rect 18555 43265 18567 43299
rect 18509 43259 18567 43265
rect 18598 43256 18604 43308
rect 18656 43296 18662 43308
rect 19444 43305 19472 43336
rect 19978 43324 19984 43336
rect 20036 43324 20042 43376
rect 20806 43364 20812 43376
rect 20767 43336 20812 43364
rect 20806 43324 20812 43336
rect 20864 43324 20870 43376
rect 21928 43305 21956 43404
rect 22741 43367 22799 43373
rect 22741 43364 22753 43367
rect 22388 43336 22753 43364
rect 22388 43308 22416 43336
rect 22741 43333 22753 43336
rect 22787 43333 22799 43367
rect 22741 43327 22799 43333
rect 19429 43299 19487 43305
rect 18656 43268 18701 43296
rect 18656 43256 18662 43268
rect 19429 43265 19441 43299
rect 19475 43265 19487 43299
rect 19705 43299 19763 43305
rect 19705 43296 19717 43299
rect 19429 43259 19487 43265
rect 19628 43268 19717 43296
rect 15289 43231 15347 43237
rect 15289 43197 15301 43231
rect 15335 43228 15347 43231
rect 15746 43228 15752 43240
rect 15335 43200 15752 43228
rect 15335 43197 15347 43200
rect 15289 43191 15347 43197
rect 15746 43188 15752 43200
rect 15804 43188 15810 43240
rect 16117 43231 16175 43237
rect 16117 43197 16129 43231
rect 16163 43228 16175 43231
rect 16163 43200 17448 43228
rect 16163 43197 16175 43200
rect 16117 43191 16175 43197
rect 15565 43163 15623 43169
rect 15565 43129 15577 43163
rect 15611 43160 15623 43163
rect 16758 43160 16764 43172
rect 15611 43132 16764 43160
rect 15611 43129 15623 43132
rect 15565 43123 15623 43129
rect 16758 43120 16764 43132
rect 16816 43120 16822 43172
rect 16666 43092 16672 43104
rect 16627 43064 16672 43092
rect 16666 43052 16672 43064
rect 16724 43052 16730 43104
rect 17420 43092 17448 43200
rect 17494 43188 17500 43240
rect 17552 43228 17558 43240
rect 17681 43231 17739 43237
rect 17681 43228 17693 43231
rect 17552 43200 17693 43228
rect 17552 43188 17558 43200
rect 17681 43197 17693 43200
rect 17727 43197 17739 43231
rect 18046 43228 18052 43240
rect 18007 43200 18052 43228
rect 17681 43191 17739 43197
rect 18046 43188 18052 43200
rect 18104 43188 18110 43240
rect 17586 43120 17592 43172
rect 17644 43160 17650 43172
rect 19444 43160 19472 43259
rect 17644 43132 19472 43160
rect 17644 43120 17650 43132
rect 19426 43092 19432 43104
rect 17420 43064 19432 43092
rect 19426 43052 19432 43064
rect 19484 43092 19490 43104
rect 19628 43092 19656 43268
rect 19705 43265 19717 43268
rect 19751 43296 19763 43299
rect 21913 43299 21971 43305
rect 21913 43296 21925 43299
rect 19751 43268 21925 43296
rect 19751 43265 19763 43268
rect 19705 43259 19763 43265
rect 21913 43265 21925 43268
rect 21959 43265 21971 43299
rect 21913 43259 21971 43265
rect 22094 43256 22100 43308
rect 22152 43296 22158 43308
rect 22370 43296 22376 43308
rect 22152 43268 22376 43296
rect 22152 43256 22158 43268
rect 22370 43256 22376 43268
rect 22428 43256 22434 43308
rect 22557 43299 22615 43305
rect 22557 43265 22569 43299
rect 22603 43296 22615 43299
rect 22848 43296 22876 43404
rect 23198 43392 23204 43404
rect 23256 43392 23262 43444
rect 25682 43392 25688 43444
rect 25740 43432 25746 43444
rect 25777 43435 25835 43441
rect 25777 43432 25789 43435
rect 25740 43404 25789 43432
rect 25740 43392 25746 43404
rect 25777 43401 25789 43404
rect 25823 43401 25835 43435
rect 27706 43432 27712 43444
rect 27667 43404 27712 43432
rect 25777 43395 25835 43401
rect 27706 43392 27712 43404
rect 27764 43392 27770 43444
rect 30098 43432 30104 43444
rect 30059 43404 30104 43432
rect 30098 43392 30104 43404
rect 30156 43392 30162 43444
rect 31021 43435 31079 43441
rect 31021 43401 31033 43435
rect 31067 43432 31079 43435
rect 31110 43432 31116 43444
rect 31067 43404 31116 43432
rect 31067 43401 31079 43404
rect 31021 43395 31079 43401
rect 31110 43392 31116 43404
rect 31168 43392 31174 43444
rect 31202 43392 31208 43444
rect 31260 43432 31266 43444
rect 31260 43404 31432 43432
rect 31260 43392 31266 43404
rect 31404 43376 31432 43404
rect 32674 43392 32680 43444
rect 32732 43432 32738 43444
rect 51626 43432 51632 43444
rect 32732 43404 51632 43432
rect 32732 43392 32738 43404
rect 51626 43392 51632 43404
rect 51684 43392 51690 43444
rect 23842 43324 23848 43376
rect 23900 43364 23906 43376
rect 24489 43367 24547 43373
rect 24489 43364 24501 43367
rect 23900 43336 24501 43364
rect 23900 43324 23906 43336
rect 24489 43333 24501 43336
rect 24535 43333 24547 43367
rect 24489 43327 24547 43333
rect 28994 43324 29000 43376
rect 29052 43364 29058 43376
rect 30006 43364 30012 43376
rect 29052 43336 30012 43364
rect 29052 43324 29058 43336
rect 30006 43324 30012 43336
rect 30064 43364 30070 43376
rect 30834 43364 30840 43376
rect 30064 43336 30512 43364
rect 30747 43336 30840 43364
rect 30064 43324 30070 43336
rect 23382 43296 23388 43308
rect 22603 43268 22876 43296
rect 22940 43268 23388 43296
rect 22603 43265 22615 43268
rect 22557 43259 22615 43265
rect 22005 43231 22063 43237
rect 22005 43197 22017 43231
rect 22051 43228 22063 43231
rect 22940 43228 22968 43268
rect 23382 43256 23388 43268
rect 23440 43256 23446 43308
rect 23566 43296 23572 43308
rect 23527 43268 23572 43296
rect 23566 43256 23572 43268
rect 23624 43256 23630 43308
rect 23661 43299 23719 43305
rect 23661 43265 23673 43299
rect 23707 43265 23719 43299
rect 23661 43259 23719 43265
rect 23753 43299 23811 43305
rect 23753 43265 23765 43299
rect 23799 43296 23811 43299
rect 23934 43296 23940 43308
rect 23799 43268 23940 43296
rect 23799 43265 23811 43268
rect 23753 43259 23811 43265
rect 22051 43200 22968 43228
rect 22051 43197 22063 43200
rect 22005 43191 22063 43197
rect 23676 43172 23704 43259
rect 23934 43256 23940 43268
rect 23992 43256 23998 43308
rect 24765 43299 24823 43305
rect 24765 43265 24777 43299
rect 24811 43296 24823 43299
rect 25314 43296 25320 43308
rect 24811 43268 25320 43296
rect 24811 43265 24823 43268
rect 24765 43259 24823 43265
rect 25314 43256 25320 43268
rect 25372 43256 25378 43308
rect 25498 43256 25504 43308
rect 25556 43296 25562 43308
rect 25593 43299 25651 43305
rect 25593 43296 25605 43299
rect 25556 43268 25605 43296
rect 25556 43256 25562 43268
rect 25593 43265 25605 43268
rect 25639 43265 25651 43299
rect 27062 43296 27068 43308
rect 27023 43268 27068 43296
rect 25593 43259 25651 43265
rect 27062 43256 27068 43268
rect 27120 43256 27126 43308
rect 27525 43299 27583 43305
rect 27525 43296 27537 43299
rect 27172 43268 27537 43296
rect 24578 43228 24584 43240
rect 24539 43200 24584 43228
rect 24578 43188 24584 43200
rect 24636 43188 24642 43240
rect 25038 43188 25044 43240
rect 25096 43188 25102 43240
rect 25406 43228 25412 43240
rect 25367 43200 25412 43228
rect 25406 43188 25412 43200
rect 25464 43188 25470 43240
rect 26418 43188 26424 43240
rect 26476 43228 26482 43240
rect 27172 43228 27200 43268
rect 27525 43265 27537 43268
rect 27571 43296 27583 43299
rect 28442 43296 28448 43308
rect 27571 43268 28448 43296
rect 27571 43265 27583 43268
rect 27525 43259 27583 43265
rect 28442 43256 28448 43268
rect 28500 43256 28506 43308
rect 28629 43299 28687 43305
rect 28629 43265 28641 43299
rect 28675 43296 28687 43299
rect 30374 43296 30380 43308
rect 28675 43268 30380 43296
rect 28675 43265 28687 43268
rect 28629 43259 28687 43265
rect 30374 43256 30380 43268
rect 30432 43256 30438 43308
rect 30484 43296 30512 43336
rect 30834 43324 30840 43336
rect 30892 43364 30898 43376
rect 31294 43364 31300 43376
rect 30892 43336 31300 43364
rect 30892 43324 30898 43336
rect 31294 43324 31300 43336
rect 31352 43324 31358 43376
rect 31386 43324 31392 43376
rect 31444 43364 31450 43376
rect 31444 43336 31537 43364
rect 31444 43324 31450 43336
rect 32582 43324 32588 43376
rect 32640 43364 32646 43376
rect 34885 43367 34943 43373
rect 34885 43364 34897 43367
rect 32640 43336 34897 43364
rect 32640 43324 32646 43336
rect 34885 43333 34897 43336
rect 34931 43333 34943 43367
rect 35986 43364 35992 43376
rect 34885 43327 34943 43333
rect 35728 43336 35992 43364
rect 31113 43299 31171 43305
rect 31113 43296 31125 43299
rect 30484 43268 31125 43296
rect 31113 43265 31125 43268
rect 31159 43265 31171 43299
rect 31113 43259 31171 43265
rect 26476 43200 27200 43228
rect 27249 43231 27307 43237
rect 26476 43188 26482 43200
rect 27249 43197 27261 43231
rect 27295 43197 27307 43231
rect 27249 43191 27307 43197
rect 27341 43231 27399 43237
rect 27341 43197 27353 43231
rect 27387 43228 27399 43231
rect 28534 43228 28540 43240
rect 27387 43200 28540 43228
rect 27387 43197 27399 43200
rect 27341 43191 27399 43197
rect 21177 43163 21235 43169
rect 21177 43129 21189 43163
rect 21223 43160 21235 43163
rect 22370 43160 22376 43172
rect 21223 43132 22376 43160
rect 21223 43129 21235 43132
rect 21177 43123 21235 43129
rect 22370 43120 22376 43132
rect 22428 43120 22434 43172
rect 23658 43120 23664 43172
rect 23716 43120 23722 43172
rect 25056 43160 25084 43188
rect 24780 43132 25084 43160
rect 19484 43064 19656 43092
rect 19889 43095 19947 43101
rect 19484 43052 19490 43064
rect 19889 43061 19901 43095
rect 19935 43092 19947 43095
rect 19978 43092 19984 43104
rect 19935 43064 19984 43092
rect 19935 43061 19947 43064
rect 19889 43055 19947 43061
rect 19978 43052 19984 43064
rect 20036 43052 20042 43104
rect 21082 43052 21088 43104
rect 21140 43092 21146 43104
rect 21269 43095 21327 43101
rect 21269 43092 21281 43095
rect 21140 43064 21281 43092
rect 21140 43052 21146 43064
rect 21269 43061 21281 43064
rect 21315 43061 21327 43095
rect 21269 43055 21327 43061
rect 22925 43095 22983 43101
rect 22925 43061 22937 43095
rect 22971 43092 22983 43095
rect 23198 43092 23204 43104
rect 22971 43064 23204 43092
rect 22971 43061 22983 43064
rect 22925 43055 22983 43061
rect 23198 43052 23204 43064
rect 23256 43052 23262 43104
rect 24029 43095 24087 43101
rect 24029 43061 24041 43095
rect 24075 43092 24087 43095
rect 24302 43092 24308 43104
rect 24075 43064 24308 43092
rect 24075 43061 24087 43064
rect 24029 43055 24087 43061
rect 24302 43052 24308 43064
rect 24360 43052 24366 43104
rect 24780 43101 24808 43132
rect 26510 43120 26516 43172
rect 26568 43160 26574 43172
rect 27264 43160 27292 43191
rect 28534 43188 28540 43200
rect 28592 43188 28598 43240
rect 31128 43228 31156 43259
rect 31202 43256 31208 43308
rect 31260 43296 31266 43308
rect 31478 43296 31484 43308
rect 31260 43268 31484 43296
rect 31260 43256 31266 43268
rect 31478 43256 31484 43268
rect 31536 43256 31542 43308
rect 32122 43256 32128 43308
rect 32180 43296 32186 43308
rect 32677 43299 32735 43305
rect 32677 43296 32689 43299
rect 32180 43268 32689 43296
rect 32180 43256 32186 43268
rect 32677 43265 32689 43268
rect 32723 43296 32735 43299
rect 33778 43296 33784 43308
rect 32723 43268 33784 43296
rect 32723 43265 32735 43268
rect 32677 43259 32735 43265
rect 33778 43256 33784 43268
rect 33836 43256 33842 43308
rect 34238 43296 34244 43308
rect 34199 43268 34244 43296
rect 34238 43256 34244 43268
rect 34296 43256 34302 43308
rect 34330 43256 34336 43308
rect 34388 43296 34394 43308
rect 34425 43299 34483 43305
rect 34425 43296 34437 43299
rect 34388 43268 34437 43296
rect 34388 43256 34394 43268
rect 34425 43265 34437 43268
rect 34471 43265 34483 43299
rect 35526 43296 35532 43308
rect 35487 43268 35532 43296
rect 34425 43259 34483 43265
rect 35526 43256 35532 43268
rect 35584 43256 35590 43308
rect 35728 43305 35756 43336
rect 35986 43324 35992 43336
rect 36044 43364 36050 43376
rect 36449 43367 36507 43373
rect 36449 43364 36461 43367
rect 36044 43336 36461 43364
rect 36044 43324 36050 43336
rect 36449 43333 36461 43336
rect 36495 43333 36507 43367
rect 36449 43327 36507 43333
rect 37182 43324 37188 43376
rect 37240 43364 37246 43376
rect 37277 43367 37335 43373
rect 37277 43364 37289 43367
rect 37240 43336 37289 43364
rect 37240 43324 37246 43336
rect 37277 43333 37289 43336
rect 37323 43333 37335 43367
rect 37826 43364 37832 43376
rect 37787 43336 37832 43364
rect 37277 43327 37335 43333
rect 37826 43324 37832 43336
rect 37884 43364 37890 43376
rect 38381 43367 38439 43373
rect 38381 43364 38393 43367
rect 37884 43336 38393 43364
rect 37884 43324 37890 43336
rect 38381 43333 38393 43336
rect 38427 43364 38439 43367
rect 38427 43336 38654 43364
rect 38427 43333 38439 43336
rect 38381 43327 38439 43333
rect 35713 43299 35771 43305
rect 35713 43265 35725 43299
rect 35759 43265 35771 43299
rect 35713 43259 35771 43265
rect 36173 43299 36231 43305
rect 36173 43265 36185 43299
rect 36219 43265 36231 43299
rect 36173 43259 36231 43265
rect 31294 43228 31300 43240
rect 31128 43200 31300 43228
rect 31294 43188 31300 43200
rect 31352 43188 31358 43240
rect 32769 43231 32827 43237
rect 32769 43197 32781 43231
rect 32815 43197 32827 43231
rect 32769 43191 32827 43197
rect 33045 43231 33103 43237
rect 33045 43197 33057 43231
rect 33091 43228 33103 43231
rect 33134 43228 33140 43240
rect 33091 43200 33140 43228
rect 33091 43197 33103 43200
rect 33045 43191 33103 43197
rect 26568 43132 27292 43160
rect 27433 43163 27491 43169
rect 26568 43120 26574 43132
rect 27433 43129 27445 43163
rect 27479 43129 27491 43163
rect 32784 43160 32812 43191
rect 33134 43188 33140 43200
rect 33192 43188 33198 43240
rect 33505 43231 33563 43237
rect 33505 43197 33517 43231
rect 33551 43228 33563 43231
rect 33962 43228 33968 43240
rect 33551 43200 33968 43228
rect 33551 43197 33563 43200
rect 33505 43191 33563 43197
rect 33962 43188 33968 43200
rect 34020 43188 34026 43240
rect 35621 43231 35679 43237
rect 35621 43197 35633 43231
rect 35667 43228 35679 43231
rect 35894 43228 35900 43240
rect 35667 43200 35900 43228
rect 35667 43197 35679 43200
rect 35621 43191 35679 43197
rect 35894 43188 35900 43200
rect 35952 43228 35958 43240
rect 36188 43228 36216 43259
rect 36262 43256 36268 43308
rect 36320 43296 36326 43308
rect 37366 43296 37372 43308
rect 36320 43268 37372 43296
rect 36320 43256 36326 43268
rect 37366 43256 37372 43268
rect 37424 43256 37430 43308
rect 37182 43228 37188 43240
rect 35952 43200 37188 43228
rect 35952 43188 35958 43200
rect 37182 43188 37188 43200
rect 37240 43188 37246 43240
rect 33686 43160 33692 43172
rect 32784 43132 33692 43160
rect 27433 43123 27491 43129
rect 24765 43095 24823 43101
rect 24765 43061 24777 43095
rect 24811 43061 24823 43095
rect 24765 43055 24823 43061
rect 24949 43095 25007 43101
rect 24949 43061 24961 43095
rect 24995 43092 25007 43095
rect 25038 43092 25044 43104
rect 24995 43064 25044 43092
rect 24995 43061 25007 43064
rect 24949 43055 25007 43061
rect 25038 43052 25044 43064
rect 25096 43052 25102 43104
rect 26421 43095 26479 43101
rect 26421 43061 26433 43095
rect 26467 43092 26479 43095
rect 27246 43092 27252 43104
rect 26467 43064 27252 43092
rect 26467 43061 26479 43064
rect 26421 43055 26479 43061
rect 27246 43052 27252 43064
rect 27304 43052 27310 43104
rect 27338 43052 27344 43104
rect 27396 43092 27402 43104
rect 27448 43092 27476 43123
rect 33686 43120 33692 43132
rect 33744 43160 33750 43172
rect 33870 43160 33876 43172
rect 33744 43132 33876 43160
rect 33744 43120 33750 43132
rect 33870 43120 33876 43132
rect 33928 43120 33934 43172
rect 38626 43160 38654 43336
rect 39942 43160 39948 43172
rect 38626 43132 39948 43160
rect 39942 43120 39948 43132
rect 40000 43120 40006 43172
rect 27396 43064 27476 43092
rect 27396 43052 27402 43064
rect 29822 43052 29828 43104
rect 29880 43092 29886 43104
rect 32398 43092 32404 43104
rect 29880 43064 32404 43092
rect 29880 43052 29886 43064
rect 32398 43052 32404 43064
rect 32456 43052 32462 43104
rect 33226 43052 33232 43104
rect 33284 43092 33290 43104
rect 33597 43095 33655 43101
rect 33597 43092 33609 43095
rect 33284 43064 33609 43092
rect 33284 43052 33290 43064
rect 33597 43061 33609 43064
rect 33643 43061 33655 43095
rect 33597 43055 33655 43061
rect 34333 43095 34391 43101
rect 34333 43061 34345 43095
rect 34379 43092 34391 43095
rect 36170 43092 36176 43104
rect 34379 43064 36176 43092
rect 34379 43061 34391 43064
rect 34333 43055 34391 43061
rect 36170 43052 36176 43064
rect 36228 43052 36234 43104
rect 36354 43052 36360 43104
rect 36412 43092 36418 43104
rect 36449 43095 36507 43101
rect 36449 43092 36461 43095
rect 36412 43064 36461 43092
rect 36412 43052 36418 43064
rect 36449 43061 36461 43064
rect 36495 43061 36507 43095
rect 36449 43055 36507 43061
rect 38378 43052 38384 43104
rect 38436 43092 38442 43104
rect 38933 43095 38991 43101
rect 38933 43092 38945 43095
rect 38436 43064 38945 43092
rect 38436 43052 38442 43064
rect 38933 43061 38945 43064
rect 38979 43061 38991 43095
rect 39482 43092 39488 43104
rect 39443 43064 39488 43092
rect 38933 43055 38991 43061
rect 39482 43052 39488 43064
rect 39540 43092 39546 43104
rect 40037 43095 40095 43101
rect 40037 43092 40049 43095
rect 39540 43064 40049 43092
rect 39540 43052 39546 43064
rect 40037 43061 40049 43064
rect 40083 43092 40095 43095
rect 40494 43092 40500 43104
rect 40083 43064 40500 43092
rect 40083 43061 40095 43064
rect 40037 43055 40095 43061
rect 40494 43052 40500 43064
rect 40552 43052 40558 43104
rect 1104 43002 54372 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 54372 43002
rect 1104 42928 54372 42950
rect 12989 42891 13047 42897
rect 12989 42857 13001 42891
rect 13035 42888 13047 42891
rect 14090 42888 14096 42900
rect 13035 42860 14096 42888
rect 13035 42857 13047 42860
rect 12989 42851 13047 42857
rect 14090 42848 14096 42860
rect 14148 42848 14154 42900
rect 14185 42891 14243 42897
rect 14185 42857 14197 42891
rect 14231 42888 14243 42891
rect 14734 42888 14740 42900
rect 14231 42860 14740 42888
rect 14231 42857 14243 42860
rect 14185 42851 14243 42857
rect 14734 42848 14740 42860
rect 14792 42848 14798 42900
rect 16850 42848 16856 42900
rect 16908 42888 16914 42900
rect 17678 42888 17684 42900
rect 16908 42860 16988 42888
rect 17639 42860 17684 42888
rect 16908 42848 16914 42860
rect 16960 42829 16988 42860
rect 17678 42848 17684 42860
rect 17736 42848 17742 42900
rect 18322 42848 18328 42900
rect 18380 42888 18386 42900
rect 18601 42891 18659 42897
rect 18601 42888 18613 42891
rect 18380 42860 18613 42888
rect 18380 42848 18386 42860
rect 18601 42857 18613 42860
rect 18647 42857 18659 42891
rect 18601 42851 18659 42857
rect 21269 42891 21327 42897
rect 21269 42857 21281 42891
rect 21315 42888 21327 42891
rect 27062 42888 27068 42900
rect 21315 42860 27068 42888
rect 21315 42857 21327 42860
rect 21269 42851 21327 42857
rect 27062 42848 27068 42860
rect 27120 42848 27126 42900
rect 28258 42848 28264 42900
rect 28316 42888 28322 42900
rect 28445 42891 28503 42897
rect 28445 42888 28457 42891
rect 28316 42860 28457 42888
rect 28316 42848 28322 42860
rect 28445 42857 28457 42860
rect 28491 42857 28503 42891
rect 28637 42891 28695 42897
rect 28637 42888 28649 42891
rect 28445 42851 28503 42857
rect 28552 42860 28649 42888
rect 16945 42823 17003 42829
rect 16945 42789 16957 42823
rect 16991 42789 17003 42823
rect 23569 42823 23627 42829
rect 16945 42783 17003 42789
rect 20824 42792 21036 42820
rect 15102 42752 15108 42764
rect 15063 42724 15108 42752
rect 15102 42712 15108 42724
rect 15160 42712 15166 42764
rect 16666 42752 16672 42764
rect 15764 42724 16672 42752
rect 14090 42684 14096 42696
rect 14051 42656 14096 42684
rect 14090 42644 14096 42656
rect 14148 42644 14154 42696
rect 14274 42644 14280 42696
rect 14332 42684 14338 42696
rect 15764 42693 15792 42724
rect 16666 42712 16672 42724
rect 16724 42712 16730 42764
rect 16853 42755 16911 42761
rect 16853 42721 16865 42755
rect 16899 42752 16911 42755
rect 17126 42752 17132 42764
rect 16899 42724 17132 42752
rect 16899 42721 16911 42724
rect 16853 42715 16911 42721
rect 17126 42712 17132 42724
rect 17184 42752 17190 42764
rect 17184 42724 17724 42752
rect 17184 42712 17190 42724
rect 15749 42687 15807 42693
rect 14332 42656 14377 42684
rect 14332 42644 14338 42656
rect 15749 42653 15761 42687
rect 15795 42653 15807 42687
rect 15749 42647 15807 42653
rect 16025 42687 16083 42693
rect 16025 42653 16037 42687
rect 16071 42653 16083 42687
rect 16758 42684 16764 42696
rect 16719 42656 16764 42684
rect 16025 42647 16083 42653
rect 13630 42576 13636 42628
rect 13688 42616 13694 42628
rect 14737 42619 14795 42625
rect 14737 42616 14749 42619
rect 13688 42588 14749 42616
rect 13688 42576 13694 42588
rect 14737 42585 14749 42588
rect 14783 42585 14795 42619
rect 14918 42616 14924 42628
rect 14879 42588 14924 42616
rect 14737 42579 14795 42585
rect 14918 42576 14924 42588
rect 14976 42576 14982 42628
rect 15378 42576 15384 42628
rect 15436 42616 15442 42628
rect 16040 42616 16068 42647
rect 16758 42644 16764 42656
rect 16816 42644 16822 42696
rect 17037 42687 17095 42693
rect 17037 42653 17049 42687
rect 17083 42684 17095 42687
rect 17218 42684 17224 42696
rect 17083 42656 17224 42684
rect 17083 42653 17095 42656
rect 17037 42647 17095 42653
rect 17218 42644 17224 42656
rect 17276 42644 17282 42696
rect 17696 42693 17724 42724
rect 18966 42712 18972 42764
rect 19024 42752 19030 42764
rect 19337 42755 19395 42761
rect 19337 42752 19349 42755
rect 19024 42724 19349 42752
rect 19024 42712 19030 42724
rect 19337 42721 19349 42724
rect 19383 42752 19395 42755
rect 20824 42752 20852 42792
rect 19383 42724 20852 42752
rect 20901 42755 20959 42761
rect 19383 42721 19395 42724
rect 19337 42715 19395 42721
rect 20901 42721 20913 42755
rect 20947 42721 20959 42755
rect 21008 42752 21036 42792
rect 23569 42789 23581 42823
rect 23615 42820 23627 42823
rect 24026 42820 24032 42832
rect 23615 42792 24032 42820
rect 23615 42789 23627 42792
rect 23569 42783 23627 42789
rect 24026 42780 24032 42792
rect 24084 42780 24090 42832
rect 27246 42820 27252 42832
rect 27159 42792 27252 42820
rect 27246 42780 27252 42792
rect 27304 42820 27310 42832
rect 27522 42820 27528 42832
rect 27304 42792 27528 42820
rect 27304 42780 27310 42792
rect 27522 42780 27528 42792
rect 27580 42780 27586 42832
rect 28074 42780 28080 42832
rect 28132 42820 28138 42832
rect 28552 42820 28580 42860
rect 28637 42857 28649 42860
rect 28683 42857 28695 42891
rect 31110 42888 31116 42900
rect 28637 42851 28695 42857
rect 29748 42860 31116 42888
rect 28132 42792 28580 42820
rect 28132 42780 28138 42792
rect 21821 42755 21879 42761
rect 21821 42752 21833 42755
rect 21008 42724 21833 42752
rect 20901 42715 20959 42721
rect 21821 42721 21833 42724
rect 21867 42721 21879 42755
rect 21821 42715 21879 42721
rect 17681 42687 17739 42693
rect 17681 42653 17693 42687
rect 17727 42653 17739 42687
rect 17681 42647 17739 42653
rect 17770 42644 17776 42696
rect 17828 42684 17834 42696
rect 19889 42687 19947 42693
rect 17828 42656 17873 42684
rect 17828 42644 17834 42656
rect 19889 42653 19901 42687
rect 19935 42684 19947 42687
rect 20070 42684 20076 42696
rect 19935 42656 20076 42684
rect 19935 42653 19947 42656
rect 19889 42647 19947 42653
rect 20070 42644 20076 42656
rect 20128 42644 20134 42696
rect 20346 42684 20352 42696
rect 20307 42656 20352 42684
rect 20346 42644 20352 42656
rect 20404 42684 20410 42696
rect 20916 42684 20944 42715
rect 20404 42656 20944 42684
rect 20993 42687 21051 42693
rect 20404 42644 20410 42656
rect 20993 42653 21005 42687
rect 21039 42653 21051 42687
rect 20993 42647 21051 42653
rect 15436 42588 16068 42616
rect 16209 42619 16267 42625
rect 15436 42576 15442 42588
rect 16209 42585 16221 42619
rect 16255 42616 16267 42619
rect 17586 42616 17592 42628
rect 16255 42588 17592 42616
rect 16255 42585 16267 42588
rect 16209 42579 16267 42585
rect 17586 42576 17592 42588
rect 17644 42576 17650 42628
rect 20254 42616 20260 42628
rect 20167 42588 20260 42616
rect 20254 42576 20260 42588
rect 20312 42616 20318 42628
rect 21008 42616 21036 42647
rect 20312 42588 21036 42616
rect 20312 42576 20318 42588
rect 2866 42508 2872 42560
rect 2924 42548 2930 42560
rect 13541 42551 13599 42557
rect 13541 42548 13553 42551
rect 2924 42520 13553 42548
rect 2924 42508 2930 42520
rect 13541 42517 13553 42520
rect 13587 42548 13599 42551
rect 14936 42548 14964 42576
rect 13587 42520 14964 42548
rect 13587 42517 13599 42520
rect 13541 42511 13599 42517
rect 15746 42508 15752 42560
rect 15804 42548 15810 42560
rect 15841 42551 15899 42557
rect 15841 42548 15853 42551
rect 15804 42520 15853 42548
rect 15804 42508 15810 42520
rect 15841 42517 15853 42520
rect 15887 42517 15899 42551
rect 15841 42511 15899 42517
rect 17221 42551 17279 42557
rect 17221 42517 17233 42551
rect 17267 42548 17279 42551
rect 17310 42548 17316 42560
rect 17267 42520 17316 42548
rect 17267 42517 17279 42520
rect 17221 42511 17279 42517
rect 17310 42508 17316 42520
rect 17368 42508 17374 42560
rect 18046 42548 18052 42560
rect 18007 42520 18052 42548
rect 18046 42508 18052 42520
rect 18104 42508 18110 42560
rect 20162 42548 20168 42560
rect 20123 42520 20168 42548
rect 20162 42508 20168 42520
rect 20220 42508 20226 42560
rect 21836 42548 21864 42715
rect 22002 42712 22008 42764
rect 22060 42752 22066 42764
rect 22094 42752 22100 42764
rect 22060 42724 22100 42752
rect 22060 42712 22066 42724
rect 22094 42712 22100 42724
rect 22152 42752 22158 42764
rect 23017 42755 23075 42761
rect 22152 42724 22968 42752
rect 22152 42712 22158 42724
rect 22940 42693 22968 42724
rect 23017 42721 23029 42755
rect 23063 42752 23075 42755
rect 23658 42752 23664 42764
rect 23063 42724 23664 42752
rect 23063 42721 23075 42724
rect 23017 42715 23075 42721
rect 23658 42712 23664 42724
rect 23716 42712 23722 42764
rect 25314 42752 25320 42764
rect 25275 42724 25320 42752
rect 25314 42712 25320 42724
rect 25372 42712 25378 42764
rect 29546 42752 29552 42764
rect 27356 42724 29552 42752
rect 22925 42687 22983 42693
rect 22925 42653 22937 42687
rect 22971 42653 22983 42687
rect 23106 42684 23112 42696
rect 23067 42656 23112 42684
rect 22925 42647 22983 42653
rect 23106 42644 23112 42656
rect 23164 42644 23170 42696
rect 23474 42644 23480 42696
rect 23532 42684 23538 42696
rect 23569 42687 23627 42693
rect 23569 42684 23581 42687
rect 23532 42656 23581 42684
rect 23532 42644 23538 42656
rect 23569 42653 23581 42656
rect 23615 42653 23627 42687
rect 23845 42687 23903 42693
rect 23845 42684 23857 42687
rect 23569 42647 23627 42653
rect 23676 42656 23857 42684
rect 23676 42616 23704 42656
rect 23845 42653 23857 42656
rect 23891 42653 23903 42687
rect 24486 42684 24492 42696
rect 23845 42647 23903 42653
rect 23952 42656 24492 42684
rect 22388 42588 23704 42616
rect 22388 42557 22416 42588
rect 22373 42551 22431 42557
rect 22373 42548 22385 42551
rect 21836 42520 22385 42548
rect 22373 42517 22385 42520
rect 22419 42517 22431 42551
rect 23676 42548 23704 42588
rect 23753 42619 23811 42625
rect 23753 42585 23765 42619
rect 23799 42616 23811 42619
rect 23952 42616 23980 42656
rect 24486 42644 24492 42656
rect 24544 42684 24550 42696
rect 24581 42687 24639 42693
rect 24581 42684 24593 42687
rect 24544 42656 24593 42684
rect 24544 42644 24550 42656
rect 24581 42653 24593 42656
rect 24627 42653 24639 42687
rect 24581 42647 24639 42653
rect 24765 42687 24823 42693
rect 24765 42653 24777 42687
rect 24811 42684 24823 42687
rect 25225 42687 25283 42693
rect 25225 42684 25237 42687
rect 24811 42656 25237 42684
rect 24811 42653 24823 42656
rect 24765 42647 24823 42653
rect 25225 42653 25237 42656
rect 25271 42653 25283 42687
rect 25406 42684 25412 42696
rect 25367 42656 25412 42684
rect 25225 42647 25283 42653
rect 25406 42644 25412 42656
rect 25464 42644 25470 42696
rect 26786 42684 26792 42696
rect 26699 42656 26792 42684
rect 26786 42644 26792 42656
rect 26844 42684 26850 42696
rect 27246 42684 27252 42696
rect 26844 42656 27252 42684
rect 26844 42644 26850 42656
rect 27246 42644 27252 42656
rect 27304 42644 27310 42696
rect 23799 42588 23980 42616
rect 24397 42619 24455 42625
rect 23799 42585 23811 42588
rect 23753 42579 23811 42585
rect 24397 42585 24409 42619
rect 24443 42616 24455 42619
rect 27356 42616 27384 42724
rect 29546 42712 29552 42724
rect 29604 42712 29610 42764
rect 29748 42761 29776 42860
rect 31110 42848 31116 42860
rect 31168 42848 31174 42900
rect 32122 42888 32128 42900
rect 32083 42860 32128 42888
rect 32122 42848 32128 42860
rect 32180 42848 32186 42900
rect 35526 42888 35532 42900
rect 32876 42860 34744 42888
rect 35487 42860 35532 42888
rect 30466 42780 30472 42832
rect 30524 42820 30530 42832
rect 32876 42820 32904 42860
rect 34054 42820 34060 42832
rect 30524 42792 32904 42820
rect 34015 42792 34060 42820
rect 30524 42780 30530 42792
rect 29733 42755 29791 42761
rect 29733 42721 29745 42755
rect 29779 42721 29791 42755
rect 29733 42715 29791 42721
rect 29917 42755 29975 42761
rect 29917 42721 29929 42755
rect 29963 42752 29975 42755
rect 31386 42752 31392 42764
rect 29963 42724 31392 42752
rect 29963 42721 29975 42724
rect 29917 42715 29975 42721
rect 31386 42712 31392 42724
rect 31444 42712 31450 42764
rect 27430 42644 27436 42696
rect 27488 42684 27494 42696
rect 27801 42687 27859 42693
rect 27801 42684 27813 42687
rect 27488 42656 27813 42684
rect 27488 42644 27494 42656
rect 27801 42653 27813 42656
rect 27847 42653 27859 42687
rect 27801 42647 27859 42653
rect 28997 42687 29055 42693
rect 28997 42653 29009 42687
rect 29043 42653 29055 42687
rect 29564 42684 29592 42712
rect 29825 42687 29883 42693
rect 29825 42684 29837 42687
rect 29564 42656 29837 42684
rect 28997 42647 29055 42653
rect 29825 42653 29837 42656
rect 29871 42653 29883 42687
rect 29825 42647 29883 42653
rect 24443 42588 27384 42616
rect 27617 42619 27675 42625
rect 24443 42585 24455 42588
rect 24397 42579 24455 42585
rect 27617 42585 27629 42619
rect 27663 42616 27675 42619
rect 28902 42616 28908 42628
rect 27663 42588 28908 42616
rect 27663 42585 27675 42588
rect 27617 42579 27675 42585
rect 24210 42548 24216 42560
rect 23676 42520 24216 42548
rect 22373 42511 22431 42517
rect 24210 42508 24216 42520
rect 24268 42548 24274 42560
rect 24412 42548 24440 42579
rect 28902 42576 28908 42588
rect 28960 42616 28966 42628
rect 29012 42616 29040 42647
rect 30006 42644 30012 42696
rect 30064 42684 30070 42696
rect 32876 42693 32904 42792
rect 34054 42780 34060 42792
rect 34112 42780 34118 42832
rect 33594 42712 33600 42764
rect 33652 42752 33658 42764
rect 34330 42752 34336 42764
rect 33652 42724 34336 42752
rect 33652 42712 33658 42724
rect 34330 42712 34336 42724
rect 34388 42712 34394 42764
rect 34716 42752 34744 42860
rect 35526 42848 35532 42860
rect 35584 42848 35590 42900
rect 35986 42888 35992 42900
rect 35947 42860 35992 42888
rect 35986 42848 35992 42860
rect 36044 42848 36050 42900
rect 36446 42848 36452 42900
rect 36504 42888 36510 42900
rect 36504 42860 38654 42888
rect 36504 42848 36510 42860
rect 36262 42780 36268 42832
rect 36320 42820 36326 42832
rect 37458 42820 37464 42832
rect 36320 42792 37464 42820
rect 36320 42780 36326 42792
rect 37458 42780 37464 42792
rect 37516 42820 37522 42832
rect 38289 42823 38347 42829
rect 38289 42820 38301 42823
rect 37516 42792 38301 42820
rect 37516 42780 37522 42792
rect 38289 42789 38301 42792
rect 38335 42789 38347 42823
rect 38626 42820 38654 42860
rect 39482 42820 39488 42832
rect 38626 42792 39488 42820
rect 38289 42783 38347 42789
rect 39482 42780 39488 42792
rect 39540 42780 39546 42832
rect 36357 42755 36415 42761
rect 36357 42752 36369 42755
rect 34716 42724 36369 42752
rect 32033 42687 32091 42693
rect 30064 42656 30109 42684
rect 30064 42644 30070 42656
rect 32033 42653 32045 42687
rect 32079 42653 32091 42687
rect 32033 42647 32091 42653
rect 32217 42687 32275 42693
rect 32217 42653 32229 42687
rect 32263 42684 32275 42687
rect 32861 42687 32919 42693
rect 32263 42656 32812 42684
rect 32263 42653 32275 42656
rect 32217 42647 32275 42653
rect 30834 42616 30840 42628
rect 28960 42588 30840 42616
rect 28960 42576 28966 42588
rect 30834 42576 30840 42588
rect 30892 42576 30898 42628
rect 31018 42576 31024 42628
rect 31076 42616 31082 42628
rect 31113 42619 31171 42625
rect 31113 42616 31125 42619
rect 31076 42588 31125 42616
rect 31076 42576 31082 42588
rect 31113 42585 31125 42588
rect 31159 42585 31171 42619
rect 32048 42616 32076 42647
rect 32677 42619 32735 42625
rect 32677 42616 32689 42619
rect 32048 42588 32689 42616
rect 31113 42579 31171 42585
rect 32677 42585 32689 42588
rect 32723 42585 32735 42619
rect 32784 42616 32812 42656
rect 32861 42653 32873 42687
rect 32907 42653 32919 42687
rect 32861 42647 32919 42653
rect 33042 42644 33048 42696
rect 33100 42684 33106 42696
rect 33100 42656 33145 42684
rect 33100 42644 33106 42656
rect 33686 42644 33692 42696
rect 33744 42684 33750 42696
rect 33781 42687 33839 42693
rect 33781 42684 33793 42687
rect 33744 42656 33793 42684
rect 33744 42644 33750 42656
rect 33781 42653 33793 42656
rect 33827 42684 33839 42687
rect 34238 42684 34244 42696
rect 33827 42656 34244 42684
rect 33827 42653 33839 42656
rect 33781 42647 33839 42653
rect 34238 42644 34244 42656
rect 34296 42644 34302 42696
rect 34716 42693 34744 42724
rect 35360 42696 35388 42724
rect 36357 42721 36369 42724
rect 36403 42752 36415 42755
rect 36722 42752 36728 42764
rect 36403 42724 36728 42752
rect 36403 42721 36415 42724
rect 36357 42715 36415 42721
rect 36722 42712 36728 42724
rect 36780 42712 36786 42764
rect 36814 42712 36820 42764
rect 36872 42752 36878 42764
rect 36872 42724 37780 42752
rect 36872 42712 36878 42724
rect 34701 42687 34759 42693
rect 34701 42653 34713 42687
rect 34747 42653 34759 42687
rect 34701 42647 34759 42653
rect 34790 42644 34796 42696
rect 34848 42684 34854 42696
rect 34885 42687 34943 42693
rect 34885 42684 34897 42687
rect 34848 42656 34897 42684
rect 34848 42644 34854 42656
rect 34885 42653 34897 42656
rect 34931 42653 34943 42687
rect 35342 42684 35348 42696
rect 35255 42656 35348 42684
rect 34885 42647 34943 42653
rect 35342 42644 35348 42656
rect 35400 42644 35406 42696
rect 35526 42684 35532 42696
rect 35487 42656 35532 42684
rect 35526 42644 35532 42656
rect 35584 42684 35590 42696
rect 36173 42687 36231 42693
rect 36173 42684 36185 42687
rect 35584 42656 36185 42684
rect 35584 42644 35590 42656
rect 36173 42653 36185 42656
rect 36219 42684 36231 42687
rect 36446 42684 36452 42696
rect 36219 42656 36452 42684
rect 36219 42653 36231 42656
rect 36173 42647 36231 42653
rect 36446 42644 36452 42656
rect 36504 42644 36510 42696
rect 36924 42693 36952 42724
rect 36909 42687 36967 42693
rect 36909 42653 36921 42687
rect 36955 42653 36967 42687
rect 36909 42647 36967 42653
rect 36998 42644 37004 42696
rect 37056 42686 37062 42696
rect 37185 42687 37243 42693
rect 37056 42658 37099 42686
rect 37056 42644 37062 42658
rect 37185 42653 37197 42687
rect 37231 42684 37243 42687
rect 37645 42687 37703 42693
rect 37645 42684 37657 42687
rect 37231 42656 37657 42684
rect 37231 42653 37243 42656
rect 37185 42647 37243 42653
rect 37645 42653 37657 42656
rect 37691 42653 37703 42687
rect 37645 42647 37703 42653
rect 34057 42619 34115 42625
rect 32784 42588 34008 42616
rect 32677 42579 32735 42585
rect 33980 42560 34008 42588
rect 34057 42585 34069 42619
rect 34103 42616 34115 42619
rect 34974 42616 34980 42628
rect 34103 42588 34980 42616
rect 34103 42585 34115 42588
rect 34057 42579 34115 42585
rect 34974 42576 34980 42588
rect 35032 42576 35038 42628
rect 37752 42616 37780 42724
rect 38654 42712 38660 42764
rect 38712 42752 38718 42764
rect 38841 42755 38899 42761
rect 38841 42752 38853 42755
rect 38712 42724 38853 42752
rect 38712 42712 38718 42724
rect 38841 42721 38853 42724
rect 38887 42752 38899 42755
rect 40034 42752 40040 42764
rect 38887 42724 40040 42752
rect 38887 42721 38899 42724
rect 38841 42715 38899 42721
rect 40034 42712 40040 42724
rect 40092 42712 40098 42764
rect 37829 42687 37887 42693
rect 37829 42653 37841 42687
rect 37875 42684 37887 42687
rect 38930 42684 38936 42696
rect 37875 42656 38936 42684
rect 37875 42653 37887 42656
rect 37829 42647 37887 42653
rect 38930 42644 38936 42656
rect 38988 42644 38994 42696
rect 39114 42616 39120 42628
rect 37752 42588 39120 42616
rect 39114 42576 39120 42588
rect 39172 42576 39178 42628
rect 40405 42619 40463 42625
rect 40405 42616 40417 42619
rect 39224 42588 40417 42616
rect 26234 42548 26240 42560
rect 24268 42520 24440 42548
rect 26195 42520 26240 42548
rect 24268 42508 24274 42520
rect 26234 42508 26240 42520
rect 26292 42548 26298 42560
rect 27433 42551 27491 42557
rect 27433 42548 27445 42551
rect 26292 42520 27445 42548
rect 26292 42508 26298 42520
rect 27433 42517 27445 42520
rect 27479 42517 27491 42551
rect 27433 42511 27491 42517
rect 27525 42551 27583 42557
rect 27525 42517 27537 42551
rect 27571 42548 27583 42551
rect 27706 42548 27712 42560
rect 27571 42520 27712 42548
rect 27571 42517 27583 42520
rect 27525 42511 27583 42517
rect 27706 42508 27712 42520
rect 27764 42548 27770 42560
rect 28166 42548 28172 42560
rect 27764 42520 28172 42548
rect 27764 42508 27770 42520
rect 28166 42508 28172 42520
rect 28224 42508 28230 42560
rect 28629 42551 28687 42557
rect 28629 42517 28641 42551
rect 28675 42548 28687 42551
rect 29549 42551 29607 42557
rect 29549 42548 29561 42551
rect 28675 42520 29561 42548
rect 28675 42517 28687 42520
rect 28629 42511 28687 42517
rect 29549 42517 29561 42520
rect 29595 42517 29607 42551
rect 29549 42511 29607 42517
rect 29638 42508 29644 42560
rect 29696 42548 29702 42560
rect 30558 42548 30564 42560
rect 29696 42520 30564 42548
rect 29696 42508 29702 42520
rect 30558 42508 30564 42520
rect 30616 42508 30622 42560
rect 33594 42508 33600 42560
rect 33652 42548 33658 42560
rect 33873 42551 33931 42557
rect 33873 42548 33885 42551
rect 33652 42520 33885 42548
rect 33652 42508 33658 42520
rect 33873 42517 33885 42520
rect 33919 42517 33931 42551
rect 33873 42511 33931 42517
rect 33962 42508 33968 42560
rect 34020 42548 34026 42560
rect 34701 42551 34759 42557
rect 34701 42548 34713 42551
rect 34020 42520 34713 42548
rect 34020 42508 34026 42520
rect 34701 42517 34713 42520
rect 34747 42517 34759 42551
rect 34701 42511 34759 42517
rect 37458 42508 37464 42560
rect 37516 42548 37522 42560
rect 37737 42551 37795 42557
rect 37737 42548 37749 42551
rect 37516 42520 37749 42548
rect 37516 42508 37522 42520
rect 37737 42517 37749 42520
rect 37783 42517 37795 42551
rect 37737 42511 37795 42517
rect 38378 42508 38384 42560
rect 38436 42548 38442 42560
rect 39224 42548 39252 42588
rect 40405 42585 40417 42588
rect 40451 42585 40463 42619
rect 40405 42579 40463 42585
rect 39942 42548 39948 42560
rect 38436 42520 39252 42548
rect 39903 42520 39948 42548
rect 38436 42508 38442 42520
rect 39942 42508 39948 42520
rect 40000 42508 40006 42560
rect 40954 42548 40960 42560
rect 40915 42520 40960 42548
rect 40954 42508 40960 42520
rect 41012 42508 41018 42560
rect 1104 42458 54372 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 54372 42458
rect 1104 42384 54372 42406
rect 14921 42347 14979 42353
rect 14921 42313 14933 42347
rect 14967 42344 14979 42347
rect 15746 42344 15752 42356
rect 14967 42316 15752 42344
rect 14967 42313 14979 42316
rect 14921 42307 14979 42313
rect 15746 42304 15752 42316
rect 15804 42344 15810 42356
rect 16666 42344 16672 42356
rect 15804 42316 15976 42344
rect 15804 42304 15810 42316
rect 15378 42236 15384 42288
rect 15436 42276 15442 42288
rect 15841 42279 15899 42285
rect 15841 42276 15853 42279
rect 15436 42248 15853 42276
rect 15436 42236 15442 42248
rect 15841 42245 15853 42248
rect 15887 42245 15899 42279
rect 15841 42239 15899 42245
rect 13630 42168 13636 42220
rect 13688 42208 13694 42220
rect 14737 42211 14795 42217
rect 14737 42208 14749 42211
rect 13688 42180 14749 42208
rect 13688 42168 13694 42180
rect 14737 42177 14749 42180
rect 14783 42177 14795 42211
rect 14737 42171 14795 42177
rect 14918 42168 14924 42220
rect 14976 42208 14982 42220
rect 14976 42180 15069 42208
rect 14976 42168 14982 42180
rect 14277 42143 14335 42149
rect 14277 42109 14289 42143
rect 14323 42140 14335 42143
rect 14936 42140 14964 42168
rect 14323 42112 14964 42140
rect 15856 42140 15884 42239
rect 15948 42208 15976 42316
rect 16040 42316 16672 42344
rect 16040 42285 16068 42316
rect 16666 42304 16672 42316
rect 16724 42304 16730 42356
rect 17037 42347 17095 42353
rect 17037 42313 17049 42347
rect 17083 42344 17095 42347
rect 17126 42344 17132 42356
rect 17083 42316 17132 42344
rect 17083 42313 17095 42316
rect 17037 42307 17095 42313
rect 17126 42304 17132 42316
rect 17184 42304 17190 42356
rect 17589 42347 17647 42353
rect 17589 42313 17601 42347
rect 17635 42344 17647 42347
rect 17770 42344 17776 42356
rect 17635 42316 17776 42344
rect 17635 42313 17647 42316
rect 17589 42307 17647 42313
rect 17770 42304 17776 42316
rect 17828 42304 17834 42356
rect 19797 42347 19855 42353
rect 19797 42313 19809 42347
rect 19843 42344 19855 42347
rect 20254 42344 20260 42356
rect 19843 42316 20260 42344
rect 19843 42313 19855 42316
rect 19797 42307 19855 42313
rect 20254 42304 20260 42316
rect 20312 42304 20318 42356
rect 20438 42304 20444 42356
rect 20496 42344 20502 42356
rect 22097 42347 22155 42353
rect 22097 42344 22109 42347
rect 20496 42316 22109 42344
rect 20496 42304 20502 42316
rect 22097 42313 22109 42316
rect 22143 42313 22155 42347
rect 22370 42344 22376 42356
rect 22331 42316 22376 42344
rect 22097 42307 22155 42313
rect 22370 42304 22376 42316
rect 22428 42304 22434 42356
rect 23385 42347 23443 42353
rect 23385 42313 23397 42347
rect 23431 42344 23443 42347
rect 23842 42344 23848 42356
rect 23431 42316 23848 42344
rect 23431 42313 23443 42316
rect 23385 42307 23443 42313
rect 23842 42304 23848 42316
rect 23900 42304 23906 42356
rect 24581 42347 24639 42353
rect 24581 42313 24593 42347
rect 24627 42344 24639 42347
rect 25406 42344 25412 42356
rect 24627 42316 25412 42344
rect 24627 42313 24639 42316
rect 24581 42307 24639 42313
rect 25406 42304 25412 42316
rect 25464 42304 25470 42356
rect 25774 42304 25780 42356
rect 25832 42344 25838 42356
rect 26326 42344 26332 42356
rect 25832 42316 26332 42344
rect 25832 42304 25838 42316
rect 26326 42304 26332 42316
rect 26384 42304 26390 42356
rect 27338 42304 27344 42356
rect 27396 42344 27402 42356
rect 27801 42347 27859 42353
rect 27801 42344 27813 42347
rect 27396 42316 27813 42344
rect 27396 42304 27402 42316
rect 27801 42313 27813 42316
rect 27847 42313 27859 42347
rect 27801 42307 27859 42313
rect 27969 42347 28027 42353
rect 27969 42313 27981 42347
rect 28015 42344 28027 42347
rect 28902 42344 28908 42356
rect 28015 42316 28908 42344
rect 28015 42313 28027 42316
rect 27969 42307 28027 42313
rect 28902 42304 28908 42316
rect 28960 42304 28966 42356
rect 29546 42344 29552 42356
rect 29507 42316 29552 42344
rect 29546 42304 29552 42316
rect 29604 42304 29610 42356
rect 30558 42304 30564 42356
rect 30616 42344 30622 42356
rect 30834 42344 30840 42356
rect 30616 42316 30840 42344
rect 30616 42304 30622 42316
rect 30834 42304 30840 42316
rect 30892 42344 30898 42356
rect 31202 42344 31208 42356
rect 30892 42316 31208 42344
rect 30892 42304 30898 42316
rect 31202 42304 31208 42316
rect 31260 42344 31266 42356
rect 31389 42347 31447 42353
rect 31389 42344 31401 42347
rect 31260 42316 31401 42344
rect 31260 42304 31266 42316
rect 31389 42313 31401 42316
rect 31435 42344 31447 42347
rect 31478 42344 31484 42356
rect 31435 42316 31484 42344
rect 31435 42313 31447 42316
rect 31389 42307 31447 42313
rect 31478 42304 31484 42316
rect 31536 42304 31542 42356
rect 34974 42344 34980 42356
rect 34935 42316 34980 42344
rect 34974 42304 34980 42316
rect 35032 42304 35038 42356
rect 35145 42347 35203 42353
rect 35145 42313 35157 42347
rect 35191 42344 35203 42347
rect 35802 42344 35808 42356
rect 35191 42316 35808 42344
rect 35191 42313 35203 42316
rect 35145 42307 35203 42313
rect 35802 42304 35808 42316
rect 35860 42304 35866 42356
rect 36449 42347 36507 42353
rect 36449 42313 36461 42347
rect 36495 42344 36507 42347
rect 36495 42316 37596 42344
rect 36495 42313 36507 42316
rect 36449 42307 36507 42313
rect 16025 42279 16083 42285
rect 16025 42245 16037 42279
rect 16071 42245 16083 42279
rect 16025 42239 16083 42245
rect 16206 42236 16212 42288
rect 16264 42276 16270 42288
rect 18874 42276 18880 42288
rect 16264 42248 18880 42276
rect 16264 42236 16270 42248
rect 18874 42236 18880 42248
rect 18932 42236 18938 42288
rect 18969 42279 19027 42285
rect 18969 42245 18981 42279
rect 19015 42276 19027 42279
rect 19426 42276 19432 42288
rect 19015 42248 19432 42276
rect 19015 42245 19027 42248
rect 18969 42239 19027 42245
rect 19426 42236 19432 42248
rect 19484 42276 19490 42288
rect 19484 42248 20944 42276
rect 19484 42236 19490 42248
rect 16117 42211 16175 42217
rect 16117 42208 16129 42211
rect 15948 42180 16129 42208
rect 16117 42177 16129 42180
rect 16163 42177 16175 42211
rect 16117 42171 16175 42177
rect 16669 42211 16727 42217
rect 16669 42177 16681 42211
rect 16715 42177 16727 42211
rect 16669 42171 16727 42177
rect 16853 42211 16911 42217
rect 16853 42177 16865 42211
rect 16899 42208 16911 42211
rect 17034 42208 17040 42220
rect 16899 42180 17040 42208
rect 16899 42177 16911 42180
rect 16853 42171 16911 42177
rect 16684 42140 16712 42171
rect 17034 42168 17040 42180
rect 17092 42168 17098 42220
rect 17402 42168 17408 42220
rect 17460 42208 17466 42220
rect 17497 42211 17555 42217
rect 17497 42208 17509 42211
rect 17460 42180 17509 42208
rect 17460 42168 17466 42180
rect 17497 42177 17509 42180
rect 17543 42177 17555 42211
rect 17497 42171 17555 42177
rect 17681 42211 17739 42217
rect 17681 42177 17693 42211
rect 17727 42208 17739 42211
rect 17862 42208 17868 42220
rect 17727 42180 17868 42208
rect 17727 42177 17739 42180
rect 17681 42171 17739 42177
rect 17862 42168 17868 42180
rect 17920 42168 17926 42220
rect 19613 42211 19671 42217
rect 19613 42177 19625 42211
rect 19659 42208 19671 42211
rect 20070 42208 20076 42220
rect 19659 42180 20076 42208
rect 19659 42177 19671 42180
rect 19613 42171 19671 42177
rect 20070 42168 20076 42180
rect 20128 42208 20134 42220
rect 20438 42208 20444 42220
rect 20128 42180 20444 42208
rect 20128 42168 20134 42180
rect 20438 42168 20444 42180
rect 20496 42168 20502 42220
rect 20714 42208 20720 42220
rect 20675 42180 20720 42208
rect 20714 42168 20720 42180
rect 20772 42168 20778 42220
rect 20916 42217 20944 42248
rect 21818 42236 21824 42288
rect 21876 42276 21882 42288
rect 22189 42279 22247 42285
rect 22189 42276 22201 42279
rect 21876 42248 22201 42276
rect 21876 42236 21882 42248
rect 22189 42245 22201 42248
rect 22235 42245 22247 42279
rect 22189 42239 22247 42245
rect 23290 42236 23296 42288
rect 23348 42276 23354 42288
rect 23937 42279 23995 42285
rect 23937 42276 23949 42279
rect 23348 42248 23949 42276
rect 23348 42236 23354 42248
rect 23937 42245 23949 42248
rect 23983 42276 23995 42279
rect 27706 42276 27712 42288
rect 23983 42248 27712 42276
rect 23983 42245 23995 42248
rect 23937 42239 23995 42245
rect 20901 42211 20959 42217
rect 20901 42177 20913 42211
rect 20947 42177 20959 42211
rect 20901 42171 20959 42177
rect 22005 42211 22063 42217
rect 22005 42177 22017 42211
rect 22051 42177 22063 42211
rect 23198 42208 23204 42220
rect 23159 42180 23204 42208
rect 22005 42171 22063 42177
rect 15856 42112 16712 42140
rect 19429 42143 19487 42149
rect 14323 42109 14335 42112
rect 14277 42103 14335 42109
rect 14936 42072 14964 42112
rect 19429 42109 19441 42143
rect 19475 42140 19487 42143
rect 19978 42140 19984 42152
rect 19475 42112 19984 42140
rect 19475 42109 19487 42112
rect 19429 42103 19487 42109
rect 19978 42100 19984 42112
rect 20036 42140 20042 42152
rect 22020 42140 22048 42171
rect 23198 42168 23204 42180
rect 23256 42168 23262 42220
rect 23382 42208 23388 42220
rect 23343 42180 23388 42208
rect 23382 42168 23388 42180
rect 23440 42168 23446 42220
rect 24210 42168 24216 42220
rect 24268 42208 24274 42220
rect 24397 42211 24455 42217
rect 24397 42208 24409 42211
rect 24268 42180 24409 42208
rect 24268 42168 24274 42180
rect 24397 42177 24409 42180
rect 24443 42177 24455 42211
rect 24397 42171 24455 42177
rect 24486 42168 24492 42220
rect 24544 42208 24550 42220
rect 27172 42217 27200 42248
rect 27706 42236 27712 42248
rect 27764 42236 27770 42288
rect 28169 42279 28227 42285
rect 28169 42245 28181 42279
rect 28215 42276 28227 42279
rect 28813 42279 28871 42285
rect 28813 42276 28825 42279
rect 28215 42248 28825 42276
rect 28215 42245 28227 42248
rect 28169 42239 28227 42245
rect 28813 42245 28825 42248
rect 28859 42245 28871 42279
rect 30742 42276 30748 42288
rect 28813 42239 28871 42245
rect 29932 42248 30748 42276
rect 24581 42211 24639 42217
rect 24581 42208 24593 42211
rect 24544 42180 24593 42208
rect 24544 42168 24550 42180
rect 24581 42177 24593 42180
rect 24627 42177 24639 42211
rect 24581 42171 24639 42177
rect 27157 42211 27215 42217
rect 27157 42177 27169 42211
rect 27203 42177 27215 42211
rect 27338 42208 27344 42220
rect 27299 42180 27344 42208
rect 27157 42171 27215 42177
rect 27338 42168 27344 42180
rect 27396 42168 27402 42220
rect 27522 42168 27528 42220
rect 27580 42208 27586 42220
rect 28184 42208 28212 42239
rect 27580 42180 28212 42208
rect 28629 42211 28687 42217
rect 28629 42206 28641 42211
rect 27580 42168 27586 42180
rect 28552 42178 28641 42206
rect 20036 42112 22048 42140
rect 20036 42100 20042 42112
rect 23106 42100 23112 42152
rect 23164 42140 23170 42152
rect 25225 42143 25283 42149
rect 25225 42140 25237 42143
rect 23164 42112 25237 42140
rect 23164 42100 23170 42112
rect 25225 42109 25237 42112
rect 25271 42140 25283 42143
rect 26234 42140 26240 42152
rect 25271 42112 26240 42140
rect 25271 42109 25283 42112
rect 25225 42103 25283 42109
rect 26234 42100 26240 42112
rect 26292 42140 26298 42152
rect 28552 42140 28580 42178
rect 28629 42177 28641 42178
rect 28675 42177 28687 42211
rect 28629 42171 28687 42177
rect 28902 42168 28908 42220
rect 28960 42208 28966 42220
rect 28960 42180 29005 42208
rect 28960 42168 28966 42180
rect 29932 42140 29960 42248
rect 30742 42236 30748 42248
rect 30800 42236 30806 42288
rect 33778 42236 33784 42288
rect 33836 42276 33842 42288
rect 35342 42276 35348 42288
rect 33836 42248 34376 42276
rect 35303 42248 35348 42276
rect 33836 42236 33842 42248
rect 30650 42208 30656 42220
rect 30708 42217 30714 42220
rect 30620 42180 30656 42208
rect 30650 42168 30656 42180
rect 30708 42171 30720 42217
rect 30926 42208 30932 42220
rect 30887 42180 30932 42208
rect 30708 42168 30714 42171
rect 30926 42168 30932 42180
rect 30984 42168 30990 42220
rect 32122 42208 32128 42220
rect 32083 42180 32128 42208
rect 32122 42168 32128 42180
rect 32180 42168 32186 42220
rect 33137 42211 33195 42217
rect 33137 42177 33149 42211
rect 33183 42208 33195 42211
rect 34054 42208 34060 42220
rect 33183 42180 33916 42208
rect 34015 42180 34060 42208
rect 33183 42177 33195 42180
rect 33137 42171 33195 42177
rect 33226 42140 33232 42152
rect 26292 42112 29960 42140
rect 33187 42112 33232 42140
rect 26292 42100 26298 42112
rect 16022 42072 16028 42084
rect 14936 42044 16028 42072
rect 16022 42032 16028 42044
rect 16080 42032 16086 42084
rect 16117 42075 16175 42081
rect 16117 42041 16129 42075
rect 16163 42072 16175 42075
rect 17678 42072 17684 42084
rect 16163 42044 17684 42072
rect 16163 42041 16175 42044
rect 16117 42035 16175 42041
rect 17678 42032 17684 42044
rect 17736 42032 17742 42084
rect 17788 42044 20576 42072
rect 13630 42004 13636 42016
rect 13591 41976 13636 42004
rect 13630 41964 13636 41976
rect 13688 41964 13694 42016
rect 14274 41964 14280 42016
rect 14332 42004 14338 42016
rect 17788 42004 17816 42044
rect 14332 41976 17816 42004
rect 18417 42007 18475 42013
rect 14332 41964 14338 41976
rect 18417 41973 18429 42007
rect 18463 42004 18475 42007
rect 18506 42004 18512 42016
rect 18463 41976 18512 42004
rect 18463 41973 18475 41976
rect 18417 41967 18475 41973
rect 18506 41964 18512 41976
rect 18564 41964 18570 42016
rect 20257 42007 20315 42013
rect 20257 41973 20269 42007
rect 20303 42004 20315 42007
rect 20438 42004 20444 42016
rect 20303 41976 20444 42004
rect 20303 41973 20315 41976
rect 20257 41967 20315 41973
rect 20438 41964 20444 41976
rect 20496 41964 20502 42016
rect 20548 42004 20576 42044
rect 21358 42032 21364 42084
rect 21416 42072 21422 42084
rect 21821 42075 21879 42081
rect 21821 42072 21833 42075
rect 21416 42044 21833 42072
rect 21416 42032 21422 42044
rect 21821 42041 21833 42044
rect 21867 42041 21879 42075
rect 21821 42035 21879 42041
rect 25869 42075 25927 42081
rect 25869 42041 25881 42075
rect 25915 42072 25927 42075
rect 26786 42072 26792 42084
rect 25915 42044 26792 42072
rect 25915 42041 25927 42044
rect 25869 42035 25927 42041
rect 26786 42032 26792 42044
rect 26844 42032 26850 42084
rect 22002 42004 22008 42016
rect 20548 41976 22008 42004
rect 22002 41964 22008 41976
rect 22060 41964 22066 42016
rect 27341 42007 27399 42013
rect 27341 41973 27353 42007
rect 27387 42004 27399 42007
rect 27890 42004 27896 42016
rect 27387 41976 27896 42004
rect 27387 41973 27399 41976
rect 27341 41967 27399 41973
rect 27890 41964 27896 41976
rect 27948 41964 27954 42016
rect 28000 42013 28028 42112
rect 33226 42100 33232 42112
rect 33284 42100 33290 42152
rect 33888 42140 33916 42180
rect 34054 42168 34060 42180
rect 34112 42168 34118 42220
rect 34348 42217 34376 42248
rect 35342 42236 35348 42248
rect 35400 42236 35406 42288
rect 36814 42276 36820 42288
rect 36096 42248 36820 42276
rect 34333 42211 34391 42217
rect 34333 42177 34345 42211
rect 34379 42177 34391 42211
rect 34333 42171 34391 42177
rect 34149 42143 34207 42149
rect 34149 42140 34161 42143
rect 33888 42112 34161 42140
rect 34149 42109 34161 42112
rect 34195 42140 34207 42143
rect 34606 42140 34612 42152
rect 34195 42112 34612 42140
rect 34195 42109 34207 42112
rect 34149 42103 34207 42109
rect 34606 42100 34612 42112
rect 34664 42100 34670 42152
rect 35360 42140 35388 42236
rect 35894 42208 35900 42220
rect 35855 42180 35900 42208
rect 35894 42168 35900 42180
rect 35952 42168 35958 42220
rect 35986 42168 35992 42220
rect 36044 42208 36050 42220
rect 36096 42217 36124 42248
rect 36814 42236 36820 42248
rect 36872 42236 36878 42288
rect 37366 42276 37372 42288
rect 37327 42248 37372 42276
rect 37366 42236 37372 42248
rect 37424 42236 37430 42288
rect 37568 42276 37596 42316
rect 38378 42304 38384 42356
rect 38436 42344 38442 42356
rect 39393 42347 39451 42353
rect 39393 42344 39405 42347
rect 38436 42316 39405 42344
rect 38436 42304 38442 42316
rect 39393 42313 39405 42316
rect 39439 42313 39451 42347
rect 40494 42344 40500 42356
rect 40455 42316 40500 42344
rect 39393 42307 39451 42313
rect 38010 42276 38016 42288
rect 37568 42248 38016 42276
rect 36081 42211 36139 42217
rect 36081 42208 36093 42211
rect 36044 42180 36093 42208
rect 36044 42168 36050 42180
rect 36081 42177 36093 42180
rect 36127 42177 36139 42211
rect 36081 42171 36139 42177
rect 36173 42211 36231 42217
rect 36173 42177 36185 42211
rect 36219 42177 36231 42211
rect 36173 42171 36231 42177
rect 36265 42211 36323 42217
rect 36265 42177 36277 42211
rect 36311 42177 36323 42211
rect 36265 42171 36323 42177
rect 36188 42140 36216 42171
rect 35360 42112 36216 42140
rect 28534 42032 28540 42084
rect 28592 42072 28598 42084
rect 28629 42075 28687 42081
rect 28629 42072 28641 42075
rect 28592 42044 28641 42072
rect 28592 42032 28598 42044
rect 28629 42041 28641 42044
rect 28675 42041 28687 42075
rect 28629 42035 28687 42041
rect 33505 42075 33563 42081
rect 33505 42041 33517 42075
rect 33551 42072 33563 42075
rect 33594 42072 33600 42084
rect 33551 42044 33600 42072
rect 33551 42041 33563 42044
rect 33505 42035 33563 42041
rect 33594 42032 33600 42044
rect 33652 42032 33658 42084
rect 33870 42032 33876 42084
rect 33928 42072 33934 42084
rect 34241 42075 34299 42081
rect 34241 42072 34253 42075
rect 33928 42044 34253 42072
rect 33928 42032 33934 42044
rect 34241 42041 34253 42044
rect 34287 42041 34299 42075
rect 34241 42035 34299 42041
rect 35526 42032 35532 42084
rect 35584 42072 35590 42084
rect 36280 42072 36308 42171
rect 37182 42168 37188 42220
rect 37240 42208 37246 42220
rect 37568 42217 37596 42248
rect 38010 42236 38016 42248
rect 38068 42236 38074 42288
rect 39408 42276 39436 42307
rect 40494 42304 40500 42316
rect 40552 42304 40558 42356
rect 41049 42279 41107 42285
rect 41049 42276 41061 42279
rect 39408 42248 41061 42276
rect 41049 42245 41061 42248
rect 41095 42245 41107 42279
rect 41049 42239 41107 42245
rect 37277 42211 37335 42217
rect 37277 42208 37289 42211
rect 37240 42180 37289 42208
rect 37240 42168 37246 42180
rect 37277 42177 37289 42180
rect 37323 42177 37335 42211
rect 37277 42171 37335 42177
rect 37553 42211 37611 42217
rect 37553 42177 37565 42211
rect 37599 42177 37611 42211
rect 37553 42171 37611 42177
rect 37826 42168 37832 42220
rect 37884 42208 37890 42220
rect 38381 42211 38439 42217
rect 38381 42208 38393 42211
rect 37884 42180 38393 42208
rect 37884 42168 37890 42180
rect 38381 42177 38393 42180
rect 38427 42177 38439 42211
rect 38381 42171 38439 42177
rect 38102 42100 38108 42152
rect 38160 42140 38166 42152
rect 38841 42143 38899 42149
rect 38841 42140 38853 42143
rect 38160 42112 38853 42140
rect 38160 42100 38166 42112
rect 38841 42109 38853 42112
rect 38887 42109 38899 42143
rect 38841 42103 38899 42109
rect 35584 42044 36308 42072
rect 35584 42032 35590 42044
rect 37366 42032 37372 42084
rect 37424 42072 37430 42084
rect 38289 42075 38347 42081
rect 38289 42072 38301 42075
rect 37424 42044 38301 42072
rect 37424 42032 37430 42044
rect 38289 42041 38301 42044
rect 38335 42041 38347 42075
rect 38289 42035 38347 42041
rect 41601 42075 41659 42081
rect 41601 42041 41613 42075
rect 41647 42041 41659 42075
rect 41601 42035 41659 42041
rect 27985 42007 28043 42013
rect 27985 41973 27997 42007
rect 28031 41973 28043 42007
rect 27985 41967 28043 41973
rect 32309 42007 32367 42013
rect 32309 41973 32321 42007
rect 32355 42004 32367 42007
rect 32398 42004 32404 42016
rect 32355 41976 32404 42004
rect 32355 41973 32367 41976
rect 32309 41967 32367 41973
rect 32398 41964 32404 41976
rect 32456 41964 32462 42016
rect 34330 41964 34336 42016
rect 34388 42004 34394 42016
rect 34517 42007 34575 42013
rect 34517 42004 34529 42007
rect 34388 41976 34529 42004
rect 34388 41964 34394 41976
rect 34517 41973 34529 41976
rect 34563 41973 34575 42007
rect 34517 41967 34575 41973
rect 34790 41964 34796 42016
rect 34848 42004 34854 42016
rect 35161 42007 35219 42013
rect 35161 42004 35173 42007
rect 34848 41976 35173 42004
rect 34848 41964 34854 41976
rect 35161 41973 35173 41976
rect 35207 41973 35219 42007
rect 35161 41967 35219 41973
rect 37550 41964 37556 42016
rect 37608 42004 37614 42016
rect 37737 42007 37795 42013
rect 37737 42004 37749 42007
rect 37608 41976 37749 42004
rect 37608 41964 37614 41976
rect 37737 41973 37749 41976
rect 37783 41973 37795 42007
rect 37737 41967 37795 41973
rect 39022 41964 39028 42016
rect 39080 42004 39086 42016
rect 40037 42007 40095 42013
rect 40037 42004 40049 42007
rect 39080 41976 40049 42004
rect 39080 41964 39086 41976
rect 40037 41973 40049 41976
rect 40083 42004 40095 42007
rect 40954 42004 40960 42016
rect 40083 41976 40960 42004
rect 40083 41973 40095 41976
rect 40037 41967 40095 41973
rect 40954 41964 40960 41976
rect 41012 42004 41018 42016
rect 41616 42004 41644 42035
rect 41012 41976 41644 42004
rect 41012 41964 41018 41976
rect 1104 41914 54372 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 54372 41914
rect 1104 41840 54372 41862
rect 13630 41760 13636 41812
rect 13688 41800 13694 41812
rect 14369 41803 14427 41809
rect 14369 41800 14381 41803
rect 13688 41772 14381 41800
rect 13688 41760 13694 41772
rect 14369 41769 14381 41772
rect 14415 41769 14427 41803
rect 14369 41763 14427 41769
rect 16942 41760 16948 41812
rect 17000 41800 17006 41812
rect 17586 41800 17592 41812
rect 17000 41772 17592 41800
rect 17000 41760 17006 41772
rect 17586 41760 17592 41772
rect 17644 41760 17650 41812
rect 18322 41760 18328 41812
rect 18380 41800 18386 41812
rect 19705 41803 19763 41809
rect 19705 41800 19717 41803
rect 18380 41772 19717 41800
rect 18380 41760 18386 41772
rect 19705 41769 19717 41772
rect 19751 41800 19763 41803
rect 24486 41800 24492 41812
rect 19751 41772 24492 41800
rect 19751 41769 19763 41772
rect 19705 41763 19763 41769
rect 24486 41760 24492 41772
rect 24544 41760 24550 41812
rect 28442 41800 28448 41812
rect 27356 41772 28448 41800
rect 21634 41732 21640 41744
rect 18064 41704 21640 41732
rect 15473 41667 15531 41673
rect 15473 41633 15485 41667
rect 15519 41664 15531 41667
rect 16577 41667 16635 41673
rect 16577 41664 16589 41667
rect 15519 41636 16589 41664
rect 15519 41633 15531 41636
rect 15473 41627 15531 41633
rect 16577 41633 16589 41636
rect 16623 41664 16635 41667
rect 18064 41664 18092 41704
rect 21634 41692 21640 41704
rect 21692 41692 21698 41744
rect 22189 41735 22247 41741
rect 22189 41701 22201 41735
rect 22235 41732 22247 41735
rect 27249 41735 27307 41741
rect 27249 41732 27261 41735
rect 22235 41704 27261 41732
rect 22235 41701 22247 41704
rect 22189 41695 22247 41701
rect 27249 41701 27261 41704
rect 27295 41701 27307 41735
rect 27249 41695 27307 41701
rect 16623 41636 18092 41664
rect 16623 41633 16635 41636
rect 16577 41627 16635 41633
rect 17972 41608 18000 41636
rect 20162 41624 20168 41676
rect 20220 41664 20226 41676
rect 21729 41667 21787 41673
rect 21729 41664 21741 41667
rect 20220 41636 21741 41664
rect 20220 41624 20226 41636
rect 21729 41633 21741 41636
rect 21775 41633 21787 41667
rect 21729 41627 21787 41633
rect 25041 41667 25099 41673
rect 25041 41633 25053 41667
rect 25087 41664 25099 41667
rect 27356 41664 27384 41772
rect 28442 41760 28448 41772
rect 28500 41760 28506 41812
rect 30374 41800 30380 41812
rect 30335 41772 30380 41800
rect 30374 41760 30380 41772
rect 30432 41760 30438 41812
rect 33505 41803 33563 41809
rect 33505 41769 33517 41803
rect 33551 41800 33563 41803
rect 33686 41800 33692 41812
rect 33551 41772 33692 41800
rect 33551 41769 33563 41772
rect 33505 41763 33563 41769
rect 33686 41760 33692 41772
rect 33744 41800 33750 41812
rect 34146 41800 34152 41812
rect 33744 41772 34152 41800
rect 33744 41760 33750 41772
rect 34146 41760 34152 41772
rect 34204 41760 34210 41812
rect 35621 41803 35679 41809
rect 35621 41769 35633 41803
rect 35667 41800 35679 41803
rect 35710 41800 35716 41812
rect 35667 41772 35716 41800
rect 35667 41769 35679 41772
rect 35621 41763 35679 41769
rect 35710 41760 35716 41772
rect 35768 41760 35774 41812
rect 38930 41800 38936 41812
rect 38891 41772 38936 41800
rect 38930 41760 38936 41772
rect 38988 41760 38994 41812
rect 39945 41803 40003 41809
rect 39945 41769 39957 41803
rect 39991 41800 40003 41803
rect 40034 41800 40040 41812
rect 39991 41772 40040 41800
rect 39991 41769 40003 41772
rect 39945 41763 40003 41769
rect 40034 41760 40040 41772
rect 40092 41800 40098 41812
rect 40402 41800 40408 41812
rect 40092 41772 40408 41800
rect 40092 41760 40098 41772
rect 40402 41760 40408 41772
rect 40460 41760 40466 41812
rect 40954 41760 40960 41812
rect 41012 41800 41018 41812
rect 41509 41803 41567 41809
rect 41509 41800 41521 41803
rect 41012 41772 41521 41800
rect 41012 41760 41018 41772
rect 41509 41769 41521 41772
rect 41555 41769 41567 41803
rect 41509 41763 41567 41769
rect 27430 41692 27436 41744
rect 27488 41732 27494 41744
rect 27488 41704 27844 41732
rect 27488 41692 27494 41704
rect 25087 41636 25636 41664
rect 25087 41633 25099 41636
rect 25041 41627 25099 41633
rect 25608 41608 25636 41636
rect 27080 41636 27384 41664
rect 17770 41596 17776 41608
rect 17731 41568 17776 41596
rect 17770 41556 17776 41568
rect 17828 41556 17834 41608
rect 17954 41596 17960 41608
rect 17867 41568 17960 41596
rect 17954 41556 17960 41568
rect 18012 41556 18018 41608
rect 18049 41599 18107 41605
rect 18049 41565 18061 41599
rect 18095 41596 18107 41599
rect 18230 41596 18236 41608
rect 18095 41568 18236 41596
rect 18095 41565 18107 41568
rect 18049 41559 18107 41565
rect 18230 41556 18236 41568
rect 18288 41556 18294 41608
rect 20254 41596 20260 41608
rect 20215 41568 20260 41596
rect 20254 41556 20260 41568
rect 20312 41556 20318 41608
rect 20438 41596 20444 41608
rect 20399 41568 20444 41596
rect 20438 41556 20444 41568
rect 20496 41556 20502 41608
rect 20625 41599 20683 41605
rect 20625 41565 20637 41599
rect 20671 41565 20683 41599
rect 20990 41596 20996 41608
rect 20951 41568 20996 41596
rect 20625 41559 20683 41565
rect 17126 41528 17132 41540
rect 17039 41500 17132 41528
rect 17126 41488 17132 41500
rect 17184 41528 17190 41540
rect 19426 41528 19432 41540
rect 17184 41500 19432 41528
rect 17184 41488 17190 41500
rect 19426 41488 19432 41500
rect 19484 41488 19490 41540
rect 20346 41488 20352 41540
rect 20404 41528 20410 41540
rect 20640 41528 20668 41559
rect 20990 41556 20996 41568
rect 21048 41556 21054 41608
rect 21174 41596 21180 41608
rect 21087 41568 21180 41596
rect 21174 41556 21180 41568
rect 21232 41596 21238 41608
rect 21818 41596 21824 41608
rect 21232 41568 21824 41596
rect 21232 41556 21238 41568
rect 21818 41556 21824 41568
rect 21876 41556 21882 41608
rect 22738 41556 22744 41608
rect 22796 41596 22802 41608
rect 23290 41596 23296 41608
rect 22796 41568 23296 41596
rect 22796 41556 22802 41568
rect 23290 41556 23296 41568
rect 23348 41596 23354 41608
rect 23477 41599 23535 41605
rect 23477 41596 23489 41599
rect 23348 41568 23489 41596
rect 23348 41556 23354 41568
rect 23477 41565 23489 41568
rect 23523 41565 23535 41599
rect 23477 41559 23535 41565
rect 24857 41599 24915 41605
rect 24857 41565 24869 41599
rect 24903 41596 24915 41599
rect 25314 41596 25320 41608
rect 24903 41568 25320 41596
rect 24903 41565 24915 41568
rect 24857 41559 24915 41565
rect 25314 41556 25320 41568
rect 25372 41556 25378 41608
rect 25498 41596 25504 41608
rect 25459 41568 25504 41596
rect 25498 41556 25504 41568
rect 25556 41556 25562 41608
rect 25590 41556 25596 41608
rect 25648 41596 25654 41608
rect 27080 41605 27108 41636
rect 25685 41599 25743 41605
rect 25685 41596 25697 41599
rect 25648 41568 25697 41596
rect 25648 41556 25654 41568
rect 25685 41565 25697 41568
rect 25731 41565 25743 41599
rect 25685 41559 25743 41565
rect 26973 41599 27031 41605
rect 26973 41565 26985 41599
rect 27019 41565 27031 41599
rect 26973 41559 27031 41565
rect 27065 41599 27123 41605
rect 27065 41565 27077 41599
rect 27111 41565 27123 41599
rect 27065 41559 27123 41565
rect 27341 41599 27399 41605
rect 27341 41565 27353 41599
rect 27387 41596 27399 41599
rect 27706 41596 27712 41608
rect 27387 41568 27712 41596
rect 27387 41565 27399 41568
rect 27341 41559 27399 41565
rect 20404 41500 20668 41528
rect 22925 41531 22983 41537
rect 20404 41488 20410 41500
rect 22925 41497 22937 41531
rect 22971 41528 22983 41531
rect 23842 41528 23848 41540
rect 22971 41500 23848 41528
rect 22971 41497 22983 41500
rect 22925 41491 22983 41497
rect 23842 41488 23848 41500
rect 23900 41488 23906 41540
rect 24670 41528 24676 41540
rect 24631 41500 24676 41528
rect 24670 41488 24676 41500
rect 24728 41488 24734 41540
rect 25869 41531 25927 41537
rect 25869 41497 25881 41531
rect 25915 41528 25927 41531
rect 26988 41528 27016 41559
rect 27706 41556 27712 41568
rect 27764 41556 27770 41608
rect 27816 41605 27844 41704
rect 37182 41692 37188 41744
rect 37240 41732 37246 41744
rect 37645 41735 37703 41741
rect 37645 41732 37657 41735
rect 37240 41704 37657 41732
rect 37240 41692 37246 41704
rect 37645 41701 37657 41704
rect 37691 41701 37703 41735
rect 37645 41695 37703 41701
rect 27890 41624 27896 41676
rect 27948 41624 27954 41676
rect 30926 41624 30932 41676
rect 30984 41664 30990 41676
rect 32125 41667 32183 41673
rect 32125 41664 32137 41667
rect 30984 41636 32137 41664
rect 30984 41624 30990 41636
rect 32125 41633 32137 41636
rect 32171 41633 32183 41667
rect 32125 41627 32183 41633
rect 34422 41624 34428 41676
rect 34480 41664 34486 41676
rect 36354 41664 36360 41676
rect 34480 41636 34928 41664
rect 36315 41636 36360 41664
rect 34480 41624 34486 41636
rect 27801 41599 27859 41605
rect 27801 41565 27813 41599
rect 27847 41565 27859 41599
rect 27908 41596 27936 41624
rect 27985 41599 28043 41605
rect 27985 41596 27997 41599
rect 27908 41568 27997 41596
rect 27801 41559 27859 41565
rect 27985 41565 27997 41568
rect 28031 41565 28043 41599
rect 27985 41559 28043 41565
rect 31570 41556 31576 41608
rect 31628 41596 31634 41608
rect 32398 41605 32404 41608
rect 31665 41599 31723 41605
rect 31665 41596 31677 41599
rect 31628 41568 31677 41596
rect 31628 41556 31634 41568
rect 31665 41565 31677 41568
rect 31711 41565 31723 41599
rect 32392 41596 32404 41605
rect 32359 41568 32404 41596
rect 31665 41559 31723 41565
rect 32392 41559 32404 41568
rect 32398 41556 32404 41559
rect 32456 41556 32462 41608
rect 34146 41556 34152 41608
rect 34204 41596 34210 41608
rect 34900 41605 34928 41636
rect 36354 41624 36360 41636
rect 36412 41624 36418 41676
rect 36998 41624 37004 41676
rect 37056 41664 37062 41676
rect 38948 41664 38976 41760
rect 40034 41664 40040 41676
rect 37056 41636 38516 41664
rect 38948 41636 40040 41664
rect 37056 41624 37062 41636
rect 34701 41599 34759 41605
rect 34701 41596 34713 41599
rect 34204 41568 34713 41596
rect 34204 41556 34210 41568
rect 34701 41565 34713 41568
rect 34747 41565 34759 41599
rect 34701 41559 34759 41565
rect 34885 41599 34943 41605
rect 34885 41565 34897 41599
rect 34931 41596 34943 41599
rect 35986 41596 35992 41608
rect 34931 41568 35992 41596
rect 34931 41565 34943 41568
rect 34885 41559 34943 41565
rect 35986 41556 35992 41568
rect 36044 41556 36050 41608
rect 36449 41599 36507 41605
rect 36449 41565 36461 41599
rect 36495 41565 36507 41599
rect 36449 41559 36507 41565
rect 37277 41599 37335 41605
rect 37277 41565 37289 41599
rect 37323 41596 37335 41599
rect 38102 41596 38108 41608
rect 37323 41568 38108 41596
rect 37323 41565 37335 41568
rect 37277 41559 37335 41565
rect 27893 41531 27951 41537
rect 27893 41528 27905 41531
rect 25915 41500 26924 41528
rect 26988 41500 27905 41528
rect 25915 41497 25927 41500
rect 25869 41491 25927 41497
rect 26896 41472 26924 41500
rect 27893 41497 27905 41500
rect 27939 41497 27951 41531
rect 27893 41491 27951 41497
rect 28994 41488 29000 41540
rect 29052 41528 29058 41540
rect 30282 41528 30288 41540
rect 29052 41500 30288 41528
rect 29052 41488 29058 41500
rect 30282 41488 30288 41500
rect 30340 41528 30346 41540
rect 32214 41528 32220 41540
rect 30340 41500 32220 41528
rect 30340 41488 30346 41500
rect 32214 41488 32220 41500
rect 32272 41528 32278 41540
rect 34057 41531 34115 41537
rect 34057 41528 34069 41531
rect 32272 41500 34069 41528
rect 32272 41488 32278 41500
rect 34057 41497 34069 41500
rect 34103 41497 34115 41531
rect 34057 41491 34115 41497
rect 34238 41488 34244 41540
rect 34296 41528 34302 41540
rect 36262 41528 36268 41540
rect 34296 41500 36268 41528
rect 34296 41488 34302 41500
rect 36262 41488 36268 41500
rect 36320 41488 36326 41540
rect 36464 41528 36492 41559
rect 38102 41556 38108 41568
rect 38160 41556 38166 41608
rect 38488 41605 38516 41636
rect 40034 41624 40040 41636
rect 40092 41624 40098 41676
rect 38473 41599 38531 41605
rect 38473 41565 38485 41599
rect 38519 41596 38531 41599
rect 38933 41599 38991 41605
rect 38933 41596 38945 41599
rect 38519 41568 38945 41596
rect 38519 41565 38531 41568
rect 38473 41559 38531 41565
rect 38933 41565 38945 41568
rect 38979 41596 38991 41599
rect 39022 41596 39028 41608
rect 38979 41568 39028 41596
rect 38979 41565 38991 41568
rect 38933 41559 38991 41565
rect 39022 41556 39028 41568
rect 39080 41556 39086 41608
rect 39114 41556 39120 41608
rect 39172 41596 39178 41608
rect 39172 41568 40540 41596
rect 39172 41556 39178 41568
rect 37458 41528 37464 41540
rect 36464 41500 37464 41528
rect 37458 41488 37464 41500
rect 37516 41488 37522 41540
rect 38289 41531 38347 41537
rect 38289 41497 38301 41531
rect 38335 41528 38347 41531
rect 39132 41528 39160 41556
rect 38335 41500 39160 41528
rect 38335 41497 38347 41500
rect 38289 41491 38347 41497
rect 16022 41460 16028 41472
rect 15983 41432 16028 41460
rect 16022 41420 16028 41432
rect 16080 41420 16086 41472
rect 18693 41463 18751 41469
rect 18693 41429 18705 41463
rect 18739 41460 18751 41463
rect 19334 41460 19340 41472
rect 18739 41432 19340 41460
rect 18739 41429 18751 41432
rect 18693 41423 18751 41429
rect 19334 41420 19340 41432
rect 19392 41420 19398 41472
rect 20165 41463 20223 41469
rect 20165 41429 20177 41463
rect 20211 41460 20223 41463
rect 20622 41460 20628 41472
rect 20211 41432 20628 41460
rect 20211 41429 20223 41432
rect 20165 41423 20223 41429
rect 20622 41420 20628 41432
rect 20680 41420 20686 41472
rect 26602 41420 26608 41472
rect 26660 41460 26666 41472
rect 26789 41463 26847 41469
rect 26789 41460 26801 41463
rect 26660 41432 26801 41460
rect 26660 41420 26666 41432
rect 26789 41429 26801 41432
rect 26835 41429 26847 41463
rect 26789 41423 26847 41429
rect 26878 41420 26884 41472
rect 26936 41420 26942 41472
rect 27062 41420 27068 41472
rect 27120 41460 27126 41472
rect 33870 41460 33876 41472
rect 27120 41432 33876 41460
rect 27120 41420 27126 41432
rect 33870 41420 33876 41432
rect 33928 41420 33934 41472
rect 33962 41420 33968 41472
rect 34020 41460 34026 41472
rect 34422 41460 34428 41472
rect 34020 41432 34428 41460
rect 34020 41420 34026 41432
rect 34422 41420 34428 41432
rect 34480 41420 34486 41472
rect 35069 41463 35127 41469
rect 35069 41429 35081 41463
rect 35115 41460 35127 41463
rect 35342 41460 35348 41472
rect 35115 41432 35348 41460
rect 35115 41429 35127 41432
rect 35069 41423 35127 41429
rect 35342 41420 35348 41432
rect 35400 41460 35406 41472
rect 35802 41460 35808 41472
rect 35400 41432 35808 41460
rect 35400 41420 35406 41432
rect 35802 41420 35808 41432
rect 35860 41420 35866 41472
rect 36081 41463 36139 41469
rect 36081 41429 36093 41463
rect 36127 41460 36139 41463
rect 36354 41460 36360 41472
rect 36127 41432 36360 41460
rect 36127 41429 36139 41432
rect 36081 41423 36139 41429
rect 36354 41420 36360 41432
rect 36412 41420 36418 41472
rect 36722 41420 36728 41472
rect 36780 41460 36786 41472
rect 37093 41463 37151 41469
rect 37093 41460 37105 41463
rect 36780 41432 37105 41460
rect 36780 41420 36786 41432
rect 37093 41429 37105 41432
rect 37139 41429 37151 41463
rect 37366 41460 37372 41472
rect 37327 41432 37372 41460
rect 37093 41423 37151 41429
rect 37366 41420 37372 41432
rect 37424 41420 37430 41472
rect 38105 41463 38163 41469
rect 38105 41429 38117 41463
rect 38151 41460 38163 41463
rect 38194 41460 38200 41472
rect 38151 41432 38200 41460
rect 38151 41429 38163 41432
rect 38105 41423 38163 41429
rect 38194 41420 38200 41432
rect 38252 41420 38258 41472
rect 40512 41469 40540 41568
rect 53374 41528 53380 41540
rect 53335 41500 53380 41528
rect 53374 41488 53380 41500
rect 53432 41488 53438 41540
rect 53558 41528 53564 41540
rect 53519 41500 53564 41528
rect 53558 41488 53564 41500
rect 53616 41488 53622 41540
rect 40497 41463 40555 41469
rect 40497 41429 40509 41463
rect 40543 41460 40555 41463
rect 41049 41463 41107 41469
rect 41049 41460 41061 41463
rect 40543 41432 41061 41460
rect 40543 41429 40555 41432
rect 40497 41423 40555 41429
rect 41049 41429 41061 41432
rect 41095 41460 41107 41463
rect 42058 41460 42064 41472
rect 41095 41432 42064 41460
rect 41095 41429 41107 41432
rect 41049 41423 41107 41429
rect 42058 41420 42064 41432
rect 42116 41460 42122 41472
rect 42613 41463 42671 41469
rect 42613 41460 42625 41463
rect 42116 41432 42625 41460
rect 42116 41420 42122 41432
rect 42613 41429 42625 41432
rect 42659 41429 42671 41463
rect 42613 41423 42671 41429
rect 52917 41463 52975 41469
rect 52917 41429 52929 41463
rect 52963 41460 52975 41463
rect 53576 41460 53604 41488
rect 52963 41432 53604 41460
rect 52963 41429 52975 41432
rect 52917 41423 52975 41429
rect 1104 41370 54372 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 54372 41370
rect 1104 41296 54372 41318
rect 16022 41256 16028 41268
rect 15983 41228 16028 41256
rect 16022 41216 16028 41228
rect 16080 41216 16086 41268
rect 17865 41259 17923 41265
rect 17865 41225 17877 41259
rect 17911 41256 17923 41259
rect 17954 41256 17960 41268
rect 17911 41228 17960 41256
rect 17911 41225 17923 41228
rect 17865 41219 17923 41225
rect 17954 41216 17960 41228
rect 18012 41256 18018 41268
rect 18138 41256 18144 41268
rect 18012 41228 18144 41256
rect 18012 41216 18018 41228
rect 18138 41216 18144 41228
rect 18196 41216 18202 41268
rect 25225 41259 25283 41265
rect 25225 41225 25237 41259
rect 25271 41256 25283 41259
rect 25498 41256 25504 41268
rect 25271 41228 25504 41256
rect 25271 41225 25283 41228
rect 25225 41219 25283 41225
rect 25498 41216 25504 41228
rect 25556 41216 25562 41268
rect 26878 41216 26884 41268
rect 26936 41256 26942 41268
rect 26936 41228 27936 41256
rect 26936 41216 26942 41228
rect 18046 41188 18052 41200
rect 17696 41160 18052 41188
rect 17696 41129 17724 41160
rect 18046 41148 18052 41160
rect 18104 41148 18110 41200
rect 26050 41148 26056 41200
rect 26108 41188 26114 41200
rect 26326 41188 26332 41200
rect 26108 41160 26332 41188
rect 26108 41148 26114 41160
rect 26326 41148 26332 41160
rect 26384 41188 26390 41200
rect 26510 41188 26516 41200
rect 26384 41160 26516 41188
rect 26384 41148 26390 41160
rect 26510 41148 26516 41160
rect 26568 41148 26574 41200
rect 27908 41188 27936 41228
rect 28166 41216 28172 41268
rect 28224 41256 28230 41268
rect 28353 41259 28411 41265
rect 28353 41256 28365 41259
rect 28224 41228 28365 41256
rect 28224 41216 28230 41228
rect 28353 41225 28365 41228
rect 28399 41225 28411 41259
rect 30285 41259 30343 41265
rect 28353 41219 28411 41225
rect 28966 41228 29684 41256
rect 28966 41188 28994 41228
rect 27908 41160 28994 41188
rect 29656 41142 29684 41228
rect 30285 41225 30297 41259
rect 30331 41256 30343 41259
rect 30650 41256 30656 41268
rect 30331 41228 30656 41256
rect 30331 41225 30343 41228
rect 30285 41219 30343 41225
rect 30650 41216 30656 41228
rect 30708 41216 30714 41268
rect 32122 41216 32128 41268
rect 32180 41256 32186 41268
rect 32217 41259 32275 41265
rect 32217 41256 32229 41259
rect 32180 41228 32229 41256
rect 32180 41216 32186 41228
rect 32217 41225 32229 41228
rect 32263 41225 32275 41259
rect 32217 41219 32275 41225
rect 34422 41216 34428 41268
rect 34480 41216 34486 41268
rect 36630 41256 36636 41268
rect 36543 41228 36636 41256
rect 36630 41216 36636 41228
rect 36688 41256 36694 41268
rect 37182 41256 37188 41268
rect 36688 41228 37188 41256
rect 36688 41216 36694 41228
rect 37182 41216 37188 41228
rect 37240 41216 37246 41268
rect 38010 41256 38016 41268
rect 37971 41228 38016 41256
rect 38010 41216 38016 41228
rect 38068 41216 38074 41268
rect 38381 41259 38439 41265
rect 38381 41225 38393 41259
rect 38427 41225 38439 41259
rect 38381 41219 38439 41225
rect 29914 41148 29920 41200
rect 29972 41188 29978 41200
rect 30745 41191 30803 41197
rect 30745 41188 30757 41191
rect 29972 41160 30757 41188
rect 29972 41148 29978 41160
rect 30745 41157 30757 41160
rect 30791 41157 30803 41191
rect 30745 41151 30803 41157
rect 32674 41148 32680 41200
rect 32732 41188 32738 41200
rect 33505 41191 33563 41197
rect 33505 41188 33517 41191
rect 32732 41160 33517 41188
rect 32732 41148 32738 41160
rect 33505 41157 33517 41160
rect 33551 41157 33563 41191
rect 33505 41151 33563 41157
rect 33594 41148 33600 41200
rect 33652 41197 33658 41200
rect 33652 41191 33681 41197
rect 33669 41157 33681 41191
rect 33652 41151 33681 41157
rect 33652 41148 33658 41151
rect 33778 41148 33784 41200
rect 33836 41188 33842 41200
rect 34440 41188 34468 41216
rect 38396 41188 38424 41219
rect 38654 41216 38660 41268
rect 38712 41256 38718 41268
rect 40957 41259 41015 41265
rect 40957 41256 40969 41259
rect 38712 41228 40969 41256
rect 38712 41216 38718 41228
rect 40957 41225 40969 41228
rect 41003 41256 41015 41259
rect 41046 41256 41052 41268
rect 41003 41228 41052 41256
rect 41003 41225 41015 41228
rect 40957 41219 41015 41225
rect 41046 41216 41052 41228
rect 41104 41256 41110 41268
rect 41104 41228 41414 41256
rect 41104 41216 41110 41228
rect 41386 41188 41414 41228
rect 41509 41191 41567 41197
rect 41509 41188 41521 41191
rect 33836 41160 38240 41188
rect 38396 41160 39344 41188
rect 41386 41160 41521 41188
rect 33836 41148 33842 41160
rect 29656 41135 29776 41142
rect 1673 41123 1731 41129
rect 1673 41089 1685 41123
rect 1719 41120 1731 41123
rect 17681 41123 17739 41129
rect 1719 41092 2268 41120
rect 1719 41089 1731 41092
rect 1673 41083 1731 41089
rect 2240 40993 2268 41092
rect 17681 41089 17693 41123
rect 17727 41089 17739 41123
rect 17681 41083 17739 41089
rect 17957 41123 18015 41129
rect 17957 41089 17969 41123
rect 18003 41120 18015 41123
rect 18230 41120 18236 41132
rect 18003 41092 18236 41120
rect 18003 41089 18015 41092
rect 17957 41083 18015 41089
rect 18230 41080 18236 41092
rect 18288 41080 18294 41132
rect 18598 41120 18604 41132
rect 18559 41092 18604 41120
rect 18598 41080 18604 41092
rect 18656 41080 18662 41132
rect 19426 41080 19432 41132
rect 19484 41120 19490 41132
rect 19705 41123 19763 41129
rect 19705 41120 19717 41123
rect 19484 41092 19717 41120
rect 19484 41080 19490 41092
rect 19705 41089 19717 41092
rect 19751 41089 19763 41123
rect 20714 41120 20720 41132
rect 20378 41092 20720 41120
rect 19705 41083 19763 41089
rect 17586 41012 17592 41064
rect 17644 41052 17650 41064
rect 18417 41055 18475 41061
rect 18417 41052 18429 41055
rect 17644 41024 18429 41052
rect 17644 41012 17650 41024
rect 18417 41021 18429 41024
rect 18463 41021 18475 41055
rect 18417 41015 18475 41021
rect 2225 40987 2283 40993
rect 2225 40953 2237 40987
rect 2271 40984 2283 40987
rect 16942 40984 16948 40996
rect 2271 40956 16948 40984
rect 2271 40953 2283 40956
rect 2225 40947 2283 40953
rect 16942 40944 16948 40956
rect 17000 40944 17006 40996
rect 17037 40987 17095 40993
rect 17037 40953 17049 40987
rect 17083 40984 17095 40987
rect 17954 40984 17960 40996
rect 17083 40956 17960 40984
rect 17083 40953 17095 40956
rect 17037 40947 17095 40953
rect 1486 40916 1492 40928
rect 1447 40888 1492 40916
rect 1486 40876 1492 40888
rect 1544 40876 1550 40928
rect 16666 40876 16672 40928
rect 16724 40916 16730 40928
rect 17052 40916 17080 40947
rect 17954 40944 17960 40956
rect 18012 40944 18018 40996
rect 18782 40984 18788 40996
rect 18743 40956 18788 40984
rect 18782 40944 18788 40956
rect 18840 40944 18846 40996
rect 19720 40984 19748 41083
rect 20714 41080 20720 41092
rect 20772 41080 20778 41132
rect 21266 41120 21272 41132
rect 21179 41092 21272 41120
rect 21266 41080 21272 41092
rect 21324 41120 21330 41132
rect 22649 41123 22707 41129
rect 22649 41120 22661 41123
rect 21324 41092 22661 41120
rect 21324 41080 21330 41092
rect 22649 41089 22661 41092
rect 22695 41120 22707 41123
rect 23658 41120 23664 41132
rect 22695 41092 23664 41120
rect 22695 41089 22707 41092
rect 22649 41083 22707 41089
rect 23658 41080 23664 41092
rect 23716 41080 23722 41132
rect 23842 41120 23848 41132
rect 23803 41092 23848 41120
rect 23842 41080 23848 41092
rect 23900 41080 23906 41132
rect 24026 41080 24032 41132
rect 24084 41120 24090 41132
rect 24581 41123 24639 41129
rect 24581 41120 24593 41123
rect 24084 41092 24593 41120
rect 24084 41080 24090 41092
rect 24581 41089 24593 41092
rect 24627 41120 24639 41123
rect 24670 41120 24676 41132
rect 24627 41092 24676 41120
rect 24627 41089 24639 41092
rect 24581 41083 24639 41089
rect 24670 41080 24676 41092
rect 24728 41120 24734 41132
rect 25041 41123 25099 41129
rect 25041 41120 25053 41123
rect 24728 41092 25053 41120
rect 24728 41080 24734 41092
rect 25041 41089 25053 41092
rect 25087 41089 25099 41123
rect 25041 41083 25099 41089
rect 25225 41123 25283 41129
rect 25225 41089 25237 41123
rect 25271 41120 25283 41123
rect 25314 41120 25320 41132
rect 25271 41092 25320 41120
rect 25271 41089 25283 41092
rect 25225 41083 25283 41089
rect 25314 41080 25320 41092
rect 25372 41080 25378 41132
rect 26786 41080 26792 41132
rect 26844 41120 26850 41132
rect 28994 41120 29000 41132
rect 26844 41092 29000 41120
rect 26844 41080 26850 41092
rect 28994 41080 29000 41092
rect 29052 41080 29058 41132
rect 29546 41120 29552 41132
rect 29459 41092 29552 41120
rect 29546 41080 29552 41092
rect 29604 41080 29610 41132
rect 29656 41129 29791 41135
rect 29656 41114 29745 41129
rect 29733 41095 29745 41114
rect 29779 41095 29791 41129
rect 29733 41089 29791 41095
rect 30112 41123 30170 41129
rect 30112 41089 30124 41123
rect 30158 41120 30170 41123
rect 30282 41120 30288 41132
rect 30158 41092 30288 41120
rect 30158 41089 30170 41092
rect 30112 41083 30170 41089
rect 30282 41080 30288 41092
rect 30340 41080 30346 41132
rect 30926 41120 30932 41132
rect 30887 41092 30932 41120
rect 30926 41080 30932 41092
rect 30984 41080 30990 41132
rect 31021 41123 31079 41129
rect 31021 41089 31033 41123
rect 31067 41089 31079 41123
rect 31021 41083 31079 41089
rect 31297 41123 31355 41129
rect 31297 41089 31309 41123
rect 31343 41089 31355 41123
rect 32398 41120 32404 41132
rect 32359 41092 32404 41120
rect 31297 41083 31355 41089
rect 20625 41055 20683 41061
rect 20625 41021 20637 41055
rect 20671 41052 20683 41055
rect 21174 41052 21180 41064
rect 20671 41024 21180 41052
rect 20671 41021 20683 41024
rect 20625 41015 20683 41021
rect 21174 41012 21180 41024
rect 21232 41012 21238 41064
rect 23382 41012 23388 41064
rect 23440 41052 23446 41064
rect 23860 41052 23888 41080
rect 24302 41052 24308 41064
rect 23440 41024 23888 41052
rect 24263 41024 24308 41052
rect 23440 41012 23446 41024
rect 24302 41012 24308 41024
rect 24360 41012 24366 41064
rect 26970 41052 26976 41064
rect 26931 41024 26976 41052
rect 26970 41012 26976 41024
rect 27028 41012 27034 41064
rect 27246 41052 27252 41064
rect 27207 41024 27252 41052
rect 27246 41012 27252 41024
rect 27304 41012 27310 41064
rect 29564 41052 29592 41080
rect 29822 41052 29828 41064
rect 27908 41024 29592 41052
rect 29783 41024 29828 41052
rect 20898 40984 20904 40996
rect 19720 40956 20904 40984
rect 20898 40944 20904 40956
rect 20956 40984 20962 40996
rect 22005 40987 22063 40993
rect 22005 40984 22017 40987
rect 20956 40956 22017 40984
rect 20956 40944 20962 40956
rect 22005 40953 22017 40956
rect 22051 40984 22063 40987
rect 22738 40984 22744 40996
rect 22051 40956 22744 40984
rect 22051 40953 22063 40956
rect 22005 40947 22063 40953
rect 22738 40944 22744 40956
rect 22796 40944 22802 40996
rect 25869 40987 25927 40993
rect 25869 40953 25881 40987
rect 25915 40984 25927 40987
rect 26234 40984 26240 40996
rect 25915 40956 26240 40984
rect 25915 40953 25927 40956
rect 25869 40947 25927 40953
rect 26234 40944 26240 40956
rect 26292 40984 26298 40996
rect 26878 40984 26884 40996
rect 26292 40956 26884 40984
rect 26292 40944 26298 40956
rect 26878 40944 26884 40956
rect 26936 40944 26942 40996
rect 17494 40916 17500 40928
rect 16724 40888 17080 40916
rect 17455 40888 17500 40916
rect 16724 40876 16730 40888
rect 17494 40876 17500 40888
rect 17552 40876 17558 40928
rect 23106 40916 23112 40928
rect 23067 40888 23112 40916
rect 23106 40876 23112 40888
rect 23164 40876 23170 40928
rect 23750 40916 23756 40928
rect 23711 40888 23756 40916
rect 23750 40876 23756 40888
rect 23808 40876 23814 40928
rect 24394 40916 24400 40928
rect 24355 40888 24400 40916
rect 24394 40876 24400 40888
rect 24452 40876 24458 40928
rect 24489 40919 24547 40925
rect 24489 40885 24501 40919
rect 24535 40916 24547 40919
rect 25038 40916 25044 40928
rect 24535 40888 25044 40916
rect 24535 40885 24547 40888
rect 24489 40879 24547 40885
rect 25038 40876 25044 40888
rect 25096 40876 25102 40928
rect 26326 40916 26332 40928
rect 26287 40888 26332 40916
rect 26326 40876 26332 40888
rect 26384 40876 26390 40928
rect 26510 40876 26516 40928
rect 26568 40916 26574 40928
rect 27154 40916 27160 40928
rect 26568 40888 27160 40916
rect 26568 40876 26574 40888
rect 27154 40876 27160 40888
rect 27212 40916 27218 40928
rect 27908 40916 27936 41024
rect 29822 41012 29828 41024
rect 29880 41012 29886 41064
rect 29914 41012 29920 41064
rect 29972 41052 29978 41064
rect 31036 41052 31064 41083
rect 29972 41024 30017 41052
rect 30944 41024 31064 41052
rect 29972 41012 29978 41024
rect 28442 40944 28448 40996
rect 28500 40984 28506 40996
rect 29730 40984 29736 40996
rect 28500 40956 29736 40984
rect 28500 40944 28506 40956
rect 29730 40944 29736 40956
rect 29788 40984 29794 40996
rect 30944 40984 30972 41024
rect 31312 40984 31340 41083
rect 32398 41080 32404 41092
rect 32456 41080 32462 41132
rect 32582 41120 32588 41132
rect 32543 41092 32588 41120
rect 32582 41080 32588 41092
rect 32640 41080 32646 41132
rect 33321 41123 33379 41129
rect 33321 41089 33333 41123
rect 33367 41089 33379 41123
rect 33321 41083 33379 41089
rect 33336 41052 33364 41083
rect 33410 41080 33416 41132
rect 33468 41120 33474 41132
rect 33468 41092 33513 41120
rect 33468 41080 33474 41092
rect 34146 41080 34152 41132
rect 34204 41120 34210 41132
rect 34425 41123 34483 41129
rect 34425 41120 34437 41123
rect 34204 41092 34437 41120
rect 34204 41080 34210 41092
rect 34425 41089 34437 41092
rect 34471 41089 34483 41123
rect 34425 41083 34483 41089
rect 34609 41123 34667 41129
rect 34609 41089 34621 41123
rect 34655 41120 34667 41123
rect 34698 41120 34704 41132
rect 34655 41092 34704 41120
rect 34655 41089 34667 41092
rect 34609 41083 34667 41089
rect 34698 41080 34704 41092
rect 34756 41080 34762 41132
rect 35621 41123 35679 41129
rect 35621 41089 35633 41123
rect 35667 41120 35679 41123
rect 35894 41120 35900 41132
rect 35667 41092 35900 41120
rect 35667 41089 35679 41092
rect 35621 41083 35679 41089
rect 35894 41080 35900 41092
rect 35952 41080 35958 41132
rect 36449 41123 36507 41129
rect 36449 41089 36461 41123
rect 36495 41089 36507 41123
rect 36449 41083 36507 41089
rect 33781 41055 33839 41061
rect 33336 41024 33456 41052
rect 29788 40956 30972 40984
rect 31036 40956 31340 40984
rect 29788 40944 29794 40956
rect 27212 40888 27936 40916
rect 27212 40876 27218 40888
rect 28534 40876 28540 40928
rect 28592 40916 28598 40928
rect 29638 40916 29644 40928
rect 28592 40888 29644 40916
rect 28592 40876 28598 40888
rect 29638 40876 29644 40888
rect 29696 40916 29702 40928
rect 31036 40916 31064 40956
rect 31202 40916 31208 40928
rect 29696 40888 31064 40916
rect 31163 40888 31208 40916
rect 29696 40876 29702 40888
rect 31202 40876 31208 40888
rect 31260 40876 31266 40928
rect 33137 40919 33195 40925
rect 33137 40885 33149 40919
rect 33183 40916 33195 40919
rect 33226 40916 33232 40928
rect 33183 40888 33232 40916
rect 33183 40885 33195 40888
rect 33137 40879 33195 40885
rect 33226 40876 33232 40888
rect 33284 40876 33290 40928
rect 33428 40916 33456 41024
rect 33781 41021 33793 41055
rect 33827 41052 33839 41055
rect 34238 41052 34244 41064
rect 33827 41024 34244 41052
rect 33827 41021 33839 41024
rect 33781 41015 33839 41021
rect 34238 41012 34244 41024
rect 34296 41012 34302 41064
rect 35437 41055 35495 41061
rect 35437 41021 35449 41055
rect 35483 41052 35495 41055
rect 36464 41052 36492 41083
rect 36722 41080 36728 41132
rect 36780 41120 36786 41132
rect 37737 41123 37795 41129
rect 36780 41092 36825 41120
rect 36780 41080 36786 41092
rect 37737 41089 37749 41123
rect 37783 41120 37795 41123
rect 37826 41120 37832 41132
rect 37783 41092 37832 41120
rect 37783 41089 37795 41092
rect 37737 41083 37795 41089
rect 37826 41080 37832 41092
rect 37884 41080 37890 41132
rect 38102 41120 38108 41132
rect 38063 41092 38108 41120
rect 38102 41080 38108 41092
rect 38160 41080 38166 41132
rect 38212 41120 38240 41160
rect 38212 41092 38424 41120
rect 35483 41024 36492 41052
rect 35483 41021 35495 41024
rect 35437 41015 35495 41021
rect 36464 40984 36492 41024
rect 38194 41012 38200 41064
rect 38252 41061 38258 41064
rect 38252 41055 38280 41061
rect 38268 41021 38280 41055
rect 38396 41052 38424 41092
rect 38654 41080 38660 41132
rect 38712 41120 38718 41132
rect 39025 41123 39083 41129
rect 39025 41120 39037 41123
rect 38712 41092 39037 41120
rect 38712 41080 38718 41092
rect 39025 41089 39037 41092
rect 39071 41089 39083 41123
rect 39025 41083 39083 41089
rect 39117 41123 39175 41129
rect 39117 41089 39129 41123
rect 39163 41120 39175 41123
rect 39206 41120 39212 41132
rect 39163 41092 39212 41120
rect 39163 41089 39175 41092
rect 39117 41083 39175 41089
rect 39206 41080 39212 41092
rect 39264 41080 39270 41132
rect 39316 41129 39344 41160
rect 41509 41157 41521 41160
rect 41555 41157 41567 41191
rect 41509 41151 41567 41157
rect 39301 41123 39359 41129
rect 39301 41089 39313 41123
rect 39347 41089 39359 41123
rect 39301 41083 39359 41089
rect 39390 41080 39396 41132
rect 39448 41120 39454 41132
rect 39448 41092 39493 41120
rect 39448 41080 39454 41092
rect 39853 41055 39911 41061
rect 39853 41052 39865 41055
rect 38396 41024 39865 41052
rect 38252 41015 38280 41021
rect 39853 41021 39865 41024
rect 39899 41021 39911 41055
rect 39853 41015 39911 41021
rect 38252 41012 38258 41015
rect 38841 40987 38899 40993
rect 38841 40984 38853 40987
rect 36464 40956 38853 40984
rect 38841 40953 38853 40956
rect 38887 40953 38899 40987
rect 38841 40947 38899 40953
rect 34241 40919 34299 40925
rect 34241 40916 34253 40919
rect 33428 40888 34253 40916
rect 34241 40885 34253 40888
rect 34287 40885 34299 40919
rect 35802 40916 35808 40928
rect 35763 40888 35808 40916
rect 34241 40879 34299 40885
rect 35802 40876 35808 40888
rect 35860 40876 35866 40928
rect 36265 40919 36323 40925
rect 36265 40885 36277 40919
rect 36311 40916 36323 40919
rect 37642 40916 37648 40928
rect 36311 40888 37648 40916
rect 36311 40885 36323 40888
rect 36265 40879 36323 40885
rect 37642 40876 37648 40888
rect 37700 40876 37706 40928
rect 40402 40916 40408 40928
rect 40363 40888 40408 40916
rect 40402 40876 40408 40888
rect 40460 40876 40466 40928
rect 41506 40876 41512 40928
rect 41564 40916 41570 40928
rect 42429 40919 42487 40925
rect 42429 40916 42441 40919
rect 41564 40888 42441 40916
rect 41564 40876 41570 40888
rect 42429 40885 42441 40888
rect 42475 40885 42487 40919
rect 42429 40879 42487 40885
rect 1104 40826 54372 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 54372 40826
rect 1104 40752 54372 40774
rect 16022 40712 16028 40724
rect 15983 40684 16028 40712
rect 16022 40672 16028 40684
rect 16080 40672 16086 40724
rect 16574 40672 16580 40724
rect 16632 40712 16638 40724
rect 17126 40712 17132 40724
rect 16632 40684 17132 40712
rect 16632 40672 16638 40684
rect 17126 40672 17132 40684
rect 17184 40672 17190 40724
rect 17957 40715 18015 40721
rect 17957 40681 17969 40715
rect 18003 40712 18015 40715
rect 18598 40712 18604 40724
rect 18003 40684 18604 40712
rect 18003 40681 18015 40684
rect 17957 40675 18015 40681
rect 18598 40672 18604 40684
rect 18656 40672 18662 40724
rect 20254 40672 20260 40724
rect 20312 40712 20318 40724
rect 20533 40715 20591 40721
rect 20533 40712 20545 40715
rect 20312 40684 20545 40712
rect 20312 40672 20318 40684
rect 20533 40681 20545 40684
rect 20579 40681 20591 40715
rect 20533 40675 20591 40681
rect 26973 40715 27031 40721
rect 26973 40681 26985 40715
rect 27019 40712 27031 40715
rect 27246 40712 27252 40724
rect 27019 40684 27252 40712
rect 27019 40681 27031 40684
rect 26973 40675 27031 40681
rect 27246 40672 27252 40684
rect 27304 40672 27310 40724
rect 30101 40715 30159 40721
rect 30101 40681 30113 40715
rect 30147 40712 30159 40715
rect 30926 40712 30932 40724
rect 30147 40684 30932 40712
rect 30147 40681 30159 40684
rect 30101 40675 30159 40681
rect 30926 40672 30932 40684
rect 30984 40672 30990 40724
rect 32398 40672 32404 40724
rect 32456 40712 32462 40724
rect 33689 40715 33747 40721
rect 33689 40712 33701 40715
rect 32456 40684 33701 40712
rect 32456 40672 32462 40684
rect 33689 40681 33701 40684
rect 33735 40681 33747 40715
rect 33689 40675 33747 40681
rect 34606 40672 34612 40724
rect 34664 40712 34670 40724
rect 35437 40715 35495 40721
rect 35437 40712 35449 40715
rect 34664 40684 35449 40712
rect 34664 40672 34670 40684
rect 35437 40681 35449 40684
rect 35483 40681 35495 40715
rect 36170 40712 36176 40724
rect 35437 40675 35495 40681
rect 35636 40684 36176 40712
rect 16666 40644 16672 40656
rect 16627 40616 16672 40644
rect 16666 40604 16672 40616
rect 16724 40604 16730 40656
rect 16942 40604 16948 40656
rect 17000 40644 17006 40656
rect 18966 40644 18972 40656
rect 17000 40616 18972 40644
rect 17000 40604 17006 40616
rect 18966 40604 18972 40616
rect 19024 40604 19030 40656
rect 23658 40644 23664 40656
rect 23216 40616 23664 40644
rect 15565 40579 15623 40585
rect 15565 40545 15577 40579
rect 15611 40576 15623 40579
rect 18138 40576 18144 40588
rect 15611 40548 18144 40576
rect 15611 40545 15623 40548
rect 15565 40539 15623 40545
rect 17972 40517 18000 40548
rect 18138 40536 18144 40548
rect 18196 40536 18202 40588
rect 18506 40536 18512 40588
rect 18564 40576 18570 40588
rect 19426 40576 19432 40588
rect 18564 40548 19432 40576
rect 18564 40536 18570 40548
rect 19426 40536 19432 40548
rect 19484 40576 19490 40588
rect 20073 40579 20131 40585
rect 20073 40576 20085 40579
rect 19484 40548 20085 40576
rect 19484 40536 19490 40548
rect 20073 40545 20085 40548
rect 20119 40576 20131 40579
rect 20119 40548 22094 40576
rect 20119 40545 20131 40548
rect 20073 40539 20131 40545
rect 17957 40511 18015 40517
rect 17052 40480 17908 40508
rect 16022 40332 16028 40384
rect 16080 40372 16086 40384
rect 17052 40372 17080 40480
rect 17678 40440 17684 40452
rect 17639 40412 17684 40440
rect 17678 40400 17684 40412
rect 17736 40400 17742 40452
rect 17880 40449 17908 40480
rect 17957 40477 17969 40511
rect 18003 40477 18015 40511
rect 17957 40471 18015 40477
rect 18046 40468 18052 40520
rect 18104 40508 18110 40520
rect 18417 40511 18475 40517
rect 18417 40508 18429 40511
rect 18104 40480 18429 40508
rect 18104 40468 18110 40480
rect 18417 40477 18429 40480
rect 18463 40477 18475 40511
rect 18417 40471 18475 40477
rect 18601 40511 18659 40517
rect 18601 40477 18613 40511
rect 18647 40508 18659 40511
rect 18782 40508 18788 40520
rect 18647 40480 18788 40508
rect 18647 40477 18659 40480
rect 18601 40471 18659 40477
rect 18782 40468 18788 40480
rect 18840 40468 18846 40520
rect 20714 40508 20720 40520
rect 20675 40480 20720 40508
rect 20714 40468 20720 40480
rect 20772 40468 20778 40520
rect 20898 40508 20904 40520
rect 20859 40480 20904 40508
rect 20898 40468 20904 40480
rect 20956 40468 20962 40520
rect 22066 40508 22094 40548
rect 22833 40511 22891 40517
rect 22833 40508 22845 40511
rect 22066 40480 22845 40508
rect 22833 40477 22845 40480
rect 22879 40477 22891 40511
rect 22833 40471 22891 40477
rect 23017 40511 23075 40517
rect 23017 40477 23029 40511
rect 23063 40508 23075 40511
rect 23216 40508 23244 40616
rect 23658 40604 23664 40616
rect 23716 40604 23722 40656
rect 27706 40604 27712 40656
rect 27764 40644 27770 40656
rect 28534 40644 28540 40656
rect 27764 40616 28540 40644
rect 27764 40604 27770 40616
rect 23290 40536 23296 40588
rect 23348 40576 23354 40588
rect 24394 40576 24400 40588
rect 23348 40548 24400 40576
rect 23348 40536 23354 40548
rect 24394 40536 24400 40548
rect 24452 40576 24458 40588
rect 24489 40579 24547 40585
rect 24489 40576 24501 40579
rect 24452 40548 24501 40576
rect 24452 40536 24458 40548
rect 24489 40545 24501 40548
rect 24535 40545 24547 40579
rect 26326 40576 26332 40588
rect 24489 40539 24547 40545
rect 25700 40548 26332 40576
rect 23063 40480 23244 40508
rect 23063 40477 23075 40480
rect 23017 40471 23075 40477
rect 17865 40443 17923 40449
rect 17865 40409 17877 40443
rect 17911 40440 17923 40443
rect 18230 40440 18236 40452
rect 17911 40412 18236 40440
rect 17911 40409 17923 40412
rect 17865 40403 17923 40409
rect 18230 40400 18236 40412
rect 18288 40440 18294 40452
rect 18874 40440 18880 40452
rect 18288 40412 18880 40440
rect 18288 40400 18294 40412
rect 18874 40400 18880 40412
rect 18932 40400 18938 40452
rect 19334 40400 19340 40452
rect 19392 40440 19398 40452
rect 19521 40443 19579 40449
rect 19521 40440 19533 40443
rect 19392 40412 19533 40440
rect 19392 40400 19398 40412
rect 19521 40409 19533 40412
rect 19567 40440 19579 40443
rect 20806 40440 20812 40452
rect 19567 40412 20812 40440
rect 19567 40409 19579 40412
rect 19521 40403 19579 40409
rect 20806 40400 20812 40412
rect 20864 40400 20870 40452
rect 22848 40440 22876 40471
rect 23382 40468 23388 40520
rect 23440 40508 23446 40520
rect 23477 40511 23535 40517
rect 23477 40508 23489 40511
rect 23440 40480 23489 40508
rect 23440 40468 23446 40480
rect 23477 40477 23489 40480
rect 23523 40477 23535 40511
rect 23477 40471 23535 40477
rect 23658 40468 23664 40520
rect 23716 40508 23722 40520
rect 24578 40508 24584 40520
rect 23716 40480 24440 40508
rect 24539 40480 24584 40508
rect 23716 40468 23722 40480
rect 23400 40440 23428 40468
rect 24118 40440 24124 40452
rect 22848 40412 23428 40440
rect 23768 40412 24124 40440
rect 16080 40344 17080 40372
rect 18509 40375 18567 40381
rect 16080 40332 16086 40344
rect 18509 40341 18521 40375
rect 18555 40372 18567 40375
rect 18690 40372 18696 40384
rect 18555 40344 18696 40372
rect 18555 40341 18567 40344
rect 18509 40335 18567 40341
rect 18690 40332 18696 40344
rect 18748 40332 18754 40384
rect 21821 40375 21879 40381
rect 21821 40341 21833 40375
rect 21867 40372 21879 40375
rect 21910 40372 21916 40384
rect 21867 40344 21916 40372
rect 21867 40341 21879 40344
rect 21821 40335 21879 40341
rect 21910 40332 21916 40344
rect 21968 40332 21974 40384
rect 22373 40375 22431 40381
rect 22373 40341 22385 40375
rect 22419 40372 22431 40375
rect 22462 40372 22468 40384
rect 22419 40344 22468 40372
rect 22419 40341 22431 40344
rect 22373 40335 22431 40341
rect 22462 40332 22468 40344
rect 22520 40332 22526 40384
rect 22925 40375 22983 40381
rect 22925 40341 22937 40375
rect 22971 40372 22983 40375
rect 23768 40372 23796 40412
rect 24118 40400 24124 40412
rect 24176 40400 24182 40452
rect 24412 40440 24440 40480
rect 24578 40468 24584 40480
rect 24636 40468 24642 40520
rect 25700 40508 25728 40548
rect 26326 40536 26332 40548
rect 26384 40536 26390 40588
rect 26602 40576 26608 40588
rect 26563 40548 26608 40576
rect 26602 40536 26608 40548
rect 26660 40536 26666 40588
rect 24688 40480 25728 40508
rect 24688 40440 24716 40480
rect 26050 40468 26056 40520
rect 26108 40508 26114 40520
rect 26237 40511 26295 40517
rect 26237 40508 26249 40511
rect 26108 40480 26249 40508
rect 26108 40468 26114 40480
rect 26237 40477 26249 40480
rect 26283 40477 26295 40511
rect 26237 40471 26295 40477
rect 26421 40511 26479 40517
rect 26421 40477 26433 40511
rect 26467 40477 26479 40511
rect 26421 40471 26479 40477
rect 26513 40511 26571 40517
rect 26513 40477 26525 40511
rect 26559 40477 26571 40511
rect 26786 40508 26792 40520
rect 26747 40480 26792 40508
rect 26513 40471 26571 40477
rect 26436 40440 26464 40471
rect 24412 40412 24716 40440
rect 24964 40412 26464 40440
rect 26528 40440 26556 40471
rect 26786 40468 26792 40480
rect 26844 40508 26850 40520
rect 27522 40508 27528 40520
rect 26844 40480 27528 40508
rect 26844 40468 26850 40480
rect 27522 40468 27528 40480
rect 27580 40508 27586 40520
rect 28460 40517 28488 40616
rect 28534 40604 28540 40616
rect 28592 40604 28598 40656
rect 31389 40647 31447 40653
rect 31389 40644 31401 40647
rect 29840 40616 31401 40644
rect 29840 40588 29868 40616
rect 31389 40613 31401 40616
rect 31435 40613 31447 40647
rect 31389 40607 31447 40613
rect 31478 40604 31484 40656
rect 31536 40644 31542 40656
rect 31536 40616 32444 40644
rect 31536 40604 31542 40616
rect 28902 40576 28908 40588
rect 28863 40548 28908 40576
rect 28902 40536 28908 40548
rect 28960 40536 28966 40588
rect 29822 40576 29828 40588
rect 29783 40548 29828 40576
rect 29822 40536 29828 40548
rect 29880 40536 29886 40588
rect 30760 40548 32260 40576
rect 30760 40520 30788 40548
rect 27709 40511 27767 40517
rect 27709 40508 27721 40511
rect 27580 40480 27721 40508
rect 27580 40468 27586 40480
rect 27709 40477 27721 40480
rect 27755 40477 27767 40511
rect 27709 40471 27767 40477
rect 28445 40511 28503 40517
rect 28445 40477 28457 40511
rect 28491 40477 28503 40511
rect 28445 40471 28503 40477
rect 29733 40511 29791 40517
rect 29733 40477 29745 40511
rect 29779 40477 29791 40511
rect 30742 40508 30748 40520
rect 30703 40480 30748 40508
rect 29733 40471 29791 40477
rect 26878 40440 26884 40452
rect 26528 40412 26884 40440
rect 22971 40344 23796 40372
rect 23845 40375 23903 40381
rect 22971 40341 22983 40344
rect 22925 40335 22983 40341
rect 23845 40341 23857 40375
rect 23891 40372 23903 40375
rect 24210 40372 24216 40384
rect 23891 40344 24216 40372
rect 23891 40341 23903 40344
rect 23845 40335 23903 40341
rect 24210 40332 24216 40344
rect 24268 40332 24274 40384
rect 24964 40381 24992 40412
rect 26878 40400 26884 40412
rect 26936 40440 26942 40452
rect 27338 40440 27344 40452
rect 26936 40412 27344 40440
rect 26936 40400 26942 40412
rect 27338 40400 27344 40412
rect 27396 40400 27402 40452
rect 29748 40440 29776 40471
rect 30742 40468 30748 40480
rect 30800 40468 30806 40520
rect 30834 40468 30840 40520
rect 30892 40508 30898 40520
rect 30892 40480 30937 40508
rect 30892 40468 30898 40480
rect 31018 40468 31024 40520
rect 31076 40508 31082 40520
rect 32232 40517 32260 40548
rect 32416 40517 32444 40616
rect 33410 40604 33416 40656
rect 33468 40644 33474 40656
rect 34793 40647 34851 40653
rect 34793 40644 34805 40647
rect 33468 40616 34805 40644
rect 33468 40604 33474 40616
rect 34793 40613 34805 40616
rect 34839 40613 34851 40647
rect 34793 40607 34851 40613
rect 33226 40576 33232 40588
rect 33187 40548 33232 40576
rect 33226 40536 33232 40548
rect 33284 40536 33290 40588
rect 33321 40579 33379 40585
rect 33321 40545 33333 40579
rect 33367 40576 33379 40579
rect 33778 40576 33784 40588
rect 33367 40548 33784 40576
rect 33367 40545 33379 40548
rect 33321 40539 33379 40545
rect 33778 40536 33784 40548
rect 33836 40536 33842 40588
rect 34146 40536 34152 40588
rect 34204 40576 34210 40588
rect 34204 40548 34928 40576
rect 34204 40536 34210 40548
rect 31573 40511 31631 40517
rect 31573 40508 31585 40511
rect 31076 40480 31585 40508
rect 31076 40468 31082 40480
rect 31573 40477 31585 40480
rect 31619 40477 31631 40511
rect 31573 40471 31631 40477
rect 31665 40511 31723 40517
rect 31665 40477 31677 40511
rect 31711 40477 31723 40511
rect 31665 40471 31723 40477
rect 32217 40511 32275 40517
rect 32217 40477 32229 40511
rect 32263 40477 32275 40511
rect 32217 40471 32275 40477
rect 32401 40511 32459 40517
rect 32401 40477 32413 40511
rect 32447 40477 32459 40511
rect 33410 40508 33416 40520
rect 33371 40480 33416 40508
rect 32401 40471 32459 40477
rect 30852 40440 30880 40468
rect 29748 40412 30880 40440
rect 31386 40400 31392 40452
rect 31444 40440 31450 40452
rect 31680 40440 31708 40471
rect 33410 40468 33416 40480
rect 33468 40468 33474 40520
rect 33502 40468 33508 40520
rect 33560 40508 33566 40520
rect 34698 40508 34704 40520
rect 33560 40480 33605 40508
rect 33796 40480 34704 40508
rect 33560 40468 33566 40480
rect 31444 40412 31708 40440
rect 31444 40400 31450 40412
rect 31588 40384 31616 40412
rect 32950 40400 32956 40452
rect 33008 40440 33014 40452
rect 33796 40440 33824 40480
rect 34698 40468 34704 40480
rect 34756 40468 34762 40520
rect 34900 40517 34928 40548
rect 34885 40511 34943 40517
rect 34885 40477 34897 40511
rect 34931 40477 34943 40511
rect 35342 40508 35348 40520
rect 35303 40480 35348 40508
rect 34885 40471 34943 40477
rect 35342 40468 35348 40480
rect 35400 40468 35406 40520
rect 35529 40511 35587 40517
rect 35529 40477 35541 40511
rect 35575 40508 35587 40511
rect 35636 40508 35664 40684
rect 36170 40672 36176 40684
rect 36228 40672 36234 40724
rect 41046 40712 41052 40724
rect 41007 40684 41052 40712
rect 41046 40672 41052 40684
rect 41104 40672 41110 40724
rect 35894 40604 35900 40656
rect 35952 40644 35958 40656
rect 35952 40616 37136 40644
rect 35952 40604 35958 40616
rect 35802 40536 35808 40588
rect 35860 40576 35866 40588
rect 36265 40579 36323 40585
rect 36265 40576 36277 40579
rect 35860 40548 36277 40576
rect 35860 40536 35866 40548
rect 36265 40545 36277 40548
rect 36311 40545 36323 40579
rect 36265 40539 36323 40545
rect 37108 40520 37136 40616
rect 37826 40604 37832 40656
rect 37884 40644 37890 40656
rect 38378 40644 38384 40656
rect 37884 40616 38384 40644
rect 37884 40604 37890 40616
rect 38378 40604 38384 40616
rect 38436 40644 38442 40656
rect 38436 40616 39896 40644
rect 38436 40604 38442 40616
rect 36630 40508 36636 40520
rect 35575 40480 35664 40508
rect 36591 40480 36636 40508
rect 35575 40477 35587 40480
rect 35529 40471 35587 40477
rect 36630 40468 36636 40480
rect 36688 40468 36694 40520
rect 36722 40468 36728 40520
rect 36780 40508 36786 40520
rect 36909 40511 36967 40517
rect 36909 40508 36921 40511
rect 36780 40480 36921 40508
rect 36780 40468 36786 40480
rect 36909 40477 36921 40480
rect 36955 40477 36967 40511
rect 36909 40471 36967 40477
rect 37090 40468 37096 40520
rect 37148 40508 37154 40520
rect 37277 40511 37335 40517
rect 37277 40508 37289 40511
rect 37148 40480 37289 40508
rect 37148 40468 37154 40480
rect 37277 40477 37289 40480
rect 37323 40477 37335 40511
rect 37277 40471 37335 40477
rect 38102 40468 38108 40520
rect 38160 40468 38166 40520
rect 38654 40468 38660 40520
rect 38712 40468 38718 40520
rect 39206 40468 39212 40520
rect 39264 40508 39270 40520
rect 39868 40517 39896 40616
rect 39853 40511 39911 40517
rect 39264 40480 39357 40508
rect 39264 40468 39270 40480
rect 39853 40477 39865 40511
rect 39899 40477 39911 40511
rect 40034 40508 40040 40520
rect 39995 40480 40040 40508
rect 39853 40471 39911 40477
rect 40034 40468 40040 40480
rect 40092 40468 40098 40520
rect 33008 40412 33824 40440
rect 33008 40400 33014 40412
rect 33870 40400 33876 40452
rect 33928 40440 33934 40452
rect 36173 40443 36231 40449
rect 36173 40440 36185 40443
rect 33928 40412 36185 40440
rect 33928 40400 33934 40412
rect 36173 40409 36185 40412
rect 36219 40409 36231 40443
rect 38120 40440 38148 40468
rect 38470 40440 38476 40452
rect 38120 40412 38476 40440
rect 36173 40403 36231 40409
rect 38470 40400 38476 40412
rect 38528 40400 38534 40452
rect 39224 40440 39252 40468
rect 39666 40440 39672 40452
rect 39224 40412 39672 40440
rect 39666 40400 39672 40412
rect 39724 40440 39730 40452
rect 41506 40440 41512 40452
rect 39724 40412 41512 40440
rect 39724 40400 39730 40412
rect 41506 40400 41512 40412
rect 41564 40440 41570 40452
rect 41601 40443 41659 40449
rect 41601 40440 41613 40443
rect 41564 40412 41613 40440
rect 41564 40400 41570 40412
rect 41601 40409 41613 40412
rect 41647 40409 41659 40443
rect 41601 40403 41659 40409
rect 24949 40375 25007 40381
rect 24949 40341 24961 40375
rect 24995 40341 25007 40375
rect 25774 40372 25780 40384
rect 25735 40344 25780 40372
rect 24949 40335 25007 40341
rect 25774 40332 25780 40344
rect 25832 40332 25838 40384
rect 26234 40332 26240 40384
rect 26292 40372 26298 40384
rect 26510 40372 26516 40384
rect 26292 40344 26516 40372
rect 26292 40332 26298 40344
rect 26510 40332 26516 40344
rect 26568 40332 26574 40384
rect 30558 40372 30564 40384
rect 30519 40344 30564 40372
rect 30558 40332 30564 40344
rect 30616 40332 30622 40384
rect 31570 40332 31576 40384
rect 31628 40332 31634 40384
rect 31754 40332 31760 40384
rect 31812 40372 31818 40384
rect 32309 40375 32367 40381
rect 32309 40372 32321 40375
rect 31812 40344 32321 40372
rect 31812 40332 31818 40344
rect 32309 40341 32321 40344
rect 32355 40341 32367 40375
rect 32309 40335 32367 40341
rect 35342 40332 35348 40384
rect 35400 40372 35406 40384
rect 35618 40372 35624 40384
rect 35400 40344 35624 40372
rect 35400 40332 35406 40344
rect 35618 40332 35624 40344
rect 35676 40332 35682 40384
rect 38102 40332 38108 40384
rect 38160 40372 38166 40384
rect 39945 40375 40003 40381
rect 39945 40372 39957 40375
rect 38160 40344 39957 40372
rect 38160 40332 38166 40344
rect 39945 40341 39957 40344
rect 39991 40341 40003 40375
rect 39945 40335 40003 40341
rect 40402 40332 40408 40384
rect 40460 40372 40466 40384
rect 40497 40375 40555 40381
rect 40497 40372 40509 40375
rect 40460 40344 40509 40372
rect 40460 40332 40466 40344
rect 40497 40341 40509 40344
rect 40543 40341 40555 40375
rect 40497 40335 40555 40341
rect 1104 40282 54372 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 54372 40282
rect 1104 40208 54372 40230
rect 16758 40128 16764 40180
rect 16816 40168 16822 40180
rect 17237 40171 17295 40177
rect 17237 40168 17249 40171
rect 16816 40140 17249 40168
rect 16816 40128 16822 40140
rect 17237 40137 17249 40140
rect 17283 40137 17295 40171
rect 17237 40131 17295 40137
rect 18325 40171 18383 40177
rect 18325 40137 18337 40171
rect 18371 40168 18383 40171
rect 20714 40168 20720 40180
rect 18371 40140 20720 40168
rect 18371 40137 18383 40140
rect 18325 40131 18383 40137
rect 20714 40128 20720 40140
rect 20772 40128 20778 40180
rect 23109 40171 23167 40177
rect 23109 40137 23121 40171
rect 23155 40168 23167 40171
rect 23934 40168 23940 40180
rect 23155 40140 23940 40168
rect 23155 40137 23167 40140
rect 23109 40131 23167 40137
rect 23934 40128 23940 40140
rect 23992 40168 23998 40180
rect 23992 40140 25544 40168
rect 23992 40128 23998 40140
rect 16942 40060 16948 40112
rect 17000 40100 17006 40112
rect 17037 40103 17095 40109
rect 17037 40100 17049 40103
rect 17000 40072 17049 40100
rect 17000 40060 17006 40072
rect 17037 40069 17049 40072
rect 17083 40100 17095 40103
rect 17494 40100 17500 40112
rect 17083 40072 17500 40100
rect 17083 40069 17095 40072
rect 17037 40063 17095 40069
rect 17494 40060 17500 40072
rect 17552 40060 17558 40112
rect 17954 40060 17960 40112
rect 18012 40100 18018 40112
rect 19153 40103 19211 40109
rect 19153 40100 19165 40103
rect 18012 40072 19165 40100
rect 18012 40060 18018 40072
rect 19153 40069 19165 40072
rect 19199 40100 19211 40103
rect 19199 40072 19840 40100
rect 19199 40069 19211 40072
rect 19153 40063 19211 40069
rect 16117 40035 16175 40041
rect 16117 40001 16129 40035
rect 16163 40032 16175 40035
rect 18969 40035 19027 40041
rect 18969 40032 18981 40035
rect 16163 40004 18981 40032
rect 16163 40001 16175 40004
rect 16117 39995 16175 40001
rect 18969 40001 18981 40004
rect 19015 40032 19027 40035
rect 19426 40032 19432 40044
rect 19015 40004 19432 40032
rect 19015 40001 19027 40004
rect 18969 39995 19027 40001
rect 19426 39992 19432 40004
rect 19484 40032 19490 40044
rect 19812 40041 19840 40072
rect 23860 40072 24348 40100
rect 19613 40035 19671 40041
rect 19613 40032 19625 40035
rect 19484 40004 19625 40032
rect 19484 39992 19490 40004
rect 19613 40001 19625 40004
rect 19659 40001 19671 40035
rect 19613 39995 19671 40001
rect 19797 40035 19855 40041
rect 19797 40001 19809 40035
rect 19843 40032 19855 40035
rect 19978 40032 19984 40044
rect 19843 40004 19984 40032
rect 19843 40001 19855 40004
rect 19797 39995 19855 40001
rect 19978 39992 19984 40004
rect 20036 39992 20042 40044
rect 20717 40035 20775 40041
rect 20717 40001 20729 40035
rect 20763 40032 20775 40035
rect 20806 40032 20812 40044
rect 20763 40004 20812 40032
rect 20763 40001 20775 40004
rect 20717 39995 20775 40001
rect 20806 39992 20812 40004
rect 20864 40032 20870 40044
rect 21266 40032 21272 40044
rect 20864 40004 21272 40032
rect 20864 39992 20870 40004
rect 21266 39992 21272 40004
rect 21324 39992 21330 40044
rect 22189 40035 22247 40041
rect 22189 40001 22201 40035
rect 22235 40001 22247 40035
rect 22189 39995 22247 40001
rect 17865 39967 17923 39973
rect 17865 39933 17877 39967
rect 17911 39933 17923 39967
rect 17865 39927 17923 39933
rect 17405 39899 17463 39905
rect 17405 39865 17417 39899
rect 17451 39896 17463 39899
rect 17880 39896 17908 39927
rect 18046 39924 18052 39976
rect 18104 39964 18110 39976
rect 19705 39967 19763 39973
rect 19705 39964 19717 39967
rect 18104 39936 19717 39964
rect 18104 39924 18110 39936
rect 19705 39933 19717 39936
rect 19751 39933 19763 39967
rect 22204 39964 22232 39995
rect 22370 39992 22376 40044
rect 22428 40032 22434 40044
rect 23201 40035 23259 40041
rect 23201 40032 23213 40035
rect 22428 40004 23213 40032
rect 22428 39992 22434 40004
rect 23201 40001 23213 40004
rect 23247 40001 23259 40035
rect 23201 39995 23259 40001
rect 23290 39992 23296 40044
rect 23348 40032 23354 40044
rect 23348 40004 23393 40032
rect 23348 39992 23354 40004
rect 22830 39964 22836 39976
rect 22204 39936 22836 39964
rect 19705 39927 19763 39933
rect 22830 39924 22836 39936
rect 22888 39924 22894 39976
rect 17451 39868 17908 39896
rect 18141 39899 18199 39905
rect 17451 39865 17463 39868
rect 17405 39859 17463 39865
rect 18141 39865 18153 39899
rect 18187 39865 18199 39899
rect 18141 39859 18199 39865
rect 22281 39899 22339 39905
rect 22281 39865 22293 39899
rect 22327 39896 22339 39899
rect 23860 39896 23888 40072
rect 23934 39992 23940 40044
rect 23992 40032 23998 40044
rect 24210 40032 24216 40044
rect 23992 40004 24037 40032
rect 24171 40004 24216 40032
rect 23992 39992 23998 40004
rect 24210 39992 24216 40004
rect 24268 39992 24274 40044
rect 24320 40032 24348 40072
rect 24578 40032 24584 40044
rect 24320 40004 24584 40032
rect 24578 39992 24584 40004
rect 24636 40032 24642 40044
rect 25516 40041 25544 40140
rect 25774 40128 25780 40180
rect 25832 40168 25838 40180
rect 27062 40168 27068 40180
rect 25832 40140 27068 40168
rect 25832 40128 25838 40140
rect 27062 40128 27068 40140
rect 27120 40168 27126 40180
rect 28074 40168 28080 40180
rect 27120 40140 28080 40168
rect 27120 40128 27126 40140
rect 28074 40128 28080 40140
rect 28132 40128 28138 40180
rect 30469 40171 30527 40177
rect 30469 40137 30481 40171
rect 30515 40168 30527 40171
rect 31202 40168 31208 40180
rect 30515 40140 31208 40168
rect 30515 40137 30527 40140
rect 30469 40131 30527 40137
rect 31202 40128 31208 40140
rect 31260 40128 31266 40180
rect 32214 40168 32220 40180
rect 32175 40140 32220 40168
rect 32214 40128 32220 40140
rect 32272 40128 32278 40180
rect 33502 40128 33508 40180
rect 33560 40168 33566 40180
rect 34241 40171 34299 40177
rect 34241 40168 34253 40171
rect 33560 40140 34253 40168
rect 33560 40128 33566 40140
rect 34241 40137 34253 40140
rect 34287 40137 34299 40171
rect 39390 40168 39396 40180
rect 34241 40131 34299 40137
rect 34348 40140 35848 40168
rect 39351 40140 39396 40168
rect 26602 40060 26608 40112
rect 26660 40100 26666 40112
rect 27154 40100 27160 40112
rect 26660 40072 27160 40100
rect 26660 40060 26666 40072
rect 27154 40060 27160 40072
rect 27212 40060 27218 40112
rect 27522 40060 27528 40112
rect 27580 40100 27586 40112
rect 29730 40100 29736 40112
rect 27580 40072 27936 40100
rect 27580 40060 27586 40072
rect 24857 40035 24915 40041
rect 24857 40032 24869 40035
rect 24636 40004 24869 40032
rect 24636 39992 24642 40004
rect 24857 40001 24869 40004
rect 24903 40001 24915 40035
rect 25041 40035 25099 40041
rect 25041 40032 25053 40035
rect 24857 39995 24915 40001
rect 24964 40004 25053 40032
rect 24964 39976 24992 40004
rect 25041 40001 25053 40004
rect 25087 40001 25099 40035
rect 25041 39995 25099 40001
rect 25501 40035 25559 40041
rect 25501 40001 25513 40035
rect 25547 40001 25559 40035
rect 25501 39995 25559 40001
rect 26326 39992 26332 40044
rect 26384 40032 26390 40044
rect 26421 40035 26479 40041
rect 26421 40032 26433 40035
rect 26384 40004 26433 40032
rect 26384 39992 26390 40004
rect 26421 40001 26433 40004
rect 26467 40032 26479 40035
rect 27338 40032 27344 40044
rect 26467 40004 27344 40032
rect 26467 40001 26479 40004
rect 26421 39995 26479 40001
rect 27338 39992 27344 40004
rect 27396 39992 27402 40044
rect 27908 40041 27936 40072
rect 29012 40072 29736 40100
rect 29012 40041 29040 40072
rect 29730 40060 29736 40072
rect 29788 40060 29794 40112
rect 34146 40060 34152 40112
rect 34204 40100 34210 40112
rect 34348 40100 34376 40140
rect 34204 40072 34376 40100
rect 34425 40103 34483 40109
rect 34204 40060 34210 40072
rect 34425 40069 34437 40103
rect 34471 40100 34483 40103
rect 34471 40072 35388 40100
rect 34471 40069 34483 40072
rect 34425 40063 34483 40069
rect 27893 40035 27951 40041
rect 27893 40001 27905 40035
rect 27939 40001 27951 40035
rect 27893 39995 27951 40001
rect 28997 40035 29055 40041
rect 28997 40001 29009 40035
rect 29043 40001 29055 40035
rect 28997 39995 29055 40001
rect 30101 40035 30159 40041
rect 30101 40001 30113 40035
rect 30147 40032 30159 40035
rect 30147 40004 30512 40032
rect 30147 40001 30159 40004
rect 30101 39995 30159 40001
rect 24118 39964 24124 39976
rect 24079 39936 24124 39964
rect 24118 39924 24124 39936
rect 24176 39964 24182 39976
rect 24946 39964 24952 39976
rect 24176 39936 24952 39964
rect 24176 39924 24182 39936
rect 24946 39924 24952 39936
rect 25004 39924 25010 39976
rect 25777 39967 25835 39973
rect 25777 39964 25789 39967
rect 25056 39936 25789 39964
rect 22327 39868 23888 39896
rect 22327 39865 22339 39868
rect 22281 39859 22339 39865
rect 17221 39831 17279 39837
rect 17221 39797 17233 39831
rect 17267 39828 17279 39831
rect 17310 39828 17316 39840
rect 17267 39800 17316 39828
rect 17267 39797 17279 39800
rect 17221 39791 17279 39797
rect 17310 39788 17316 39800
rect 17368 39788 17374 39840
rect 17494 39788 17500 39840
rect 17552 39828 17558 39840
rect 18156 39828 18184 39859
rect 24210 39856 24216 39908
rect 24268 39896 24274 39908
rect 25056 39896 25084 39936
rect 25777 39933 25789 39936
rect 25823 39933 25835 39967
rect 27062 39964 27068 39976
rect 27023 39936 27068 39964
rect 25777 39927 25835 39933
rect 27062 39924 27068 39936
rect 27120 39924 27126 39976
rect 27249 39967 27307 39973
rect 27249 39933 27261 39967
rect 27295 39964 27307 39967
rect 27430 39964 27436 39976
rect 27295 39936 27436 39964
rect 27295 39933 27307 39936
rect 27249 39927 27307 39933
rect 27430 39924 27436 39936
rect 27488 39924 27494 39976
rect 30006 39964 30012 39976
rect 29967 39936 30012 39964
rect 30006 39924 30012 39936
rect 30064 39924 30070 39976
rect 30484 39964 30512 40004
rect 30558 39992 30564 40044
rect 30616 40032 30622 40044
rect 30929 40035 30987 40041
rect 30929 40032 30941 40035
rect 30616 40004 30941 40032
rect 30616 39992 30622 40004
rect 30929 40001 30941 40004
rect 30975 40001 30987 40035
rect 30929 39995 30987 40001
rect 31110 39992 31116 40044
rect 31168 40032 31174 40044
rect 31754 40032 31760 40044
rect 31168 40004 31760 40032
rect 31168 39992 31174 40004
rect 31754 39992 31760 40004
rect 31812 39992 31818 40044
rect 32950 39992 32956 40044
rect 33008 40032 33014 40044
rect 33045 40035 33103 40041
rect 33045 40032 33057 40035
rect 33008 40004 33057 40032
rect 33008 39992 33014 40004
rect 33045 40001 33057 40004
rect 33091 40001 33103 40035
rect 33045 39995 33103 40001
rect 33137 40035 33195 40041
rect 33137 40001 33149 40035
rect 33183 40001 33195 40035
rect 33318 40032 33324 40044
rect 33279 40004 33324 40032
rect 33137 39995 33195 40001
rect 30742 39964 30748 39976
rect 30484 39936 30748 39964
rect 30742 39924 30748 39936
rect 30800 39964 30806 39976
rect 31021 39967 31079 39973
rect 31021 39964 31033 39967
rect 30800 39936 31033 39964
rect 30800 39924 30806 39936
rect 31021 39933 31033 39936
rect 31067 39933 31079 39967
rect 33152 39964 33180 39995
rect 33318 39992 33324 40004
rect 33376 39992 33382 40044
rect 34609 40035 34667 40041
rect 34609 40001 34621 40035
rect 34655 40032 34667 40035
rect 34790 40032 34796 40044
rect 34655 40004 34796 40032
rect 34655 40001 34667 40004
rect 34609 39995 34667 40001
rect 34790 39992 34796 40004
rect 34848 39992 34854 40044
rect 33502 39964 33508 39976
rect 33152 39936 33508 39964
rect 31021 39927 31079 39933
rect 33502 39924 33508 39936
rect 33560 39964 33566 39976
rect 34146 39964 34152 39976
rect 33560 39936 34152 39964
rect 33560 39924 33566 39936
rect 34146 39924 34152 39936
rect 34204 39924 34210 39976
rect 25593 39899 25651 39905
rect 25593 39896 25605 39899
rect 24268 39868 25084 39896
rect 25148 39868 25605 39896
rect 24268 39856 24274 39868
rect 18782 39828 18788 39840
rect 17552 39800 18184 39828
rect 18743 39800 18788 39828
rect 17552 39788 17558 39800
rect 18782 39788 18788 39800
rect 18840 39788 18846 39840
rect 21174 39828 21180 39840
rect 21135 39800 21180 39828
rect 21174 39788 21180 39800
rect 21232 39788 21238 39840
rect 23474 39788 23480 39840
rect 23532 39828 23538 39840
rect 23753 39831 23811 39837
rect 23753 39828 23765 39831
rect 23532 39800 23765 39828
rect 23532 39788 23538 39800
rect 23753 39797 23765 39800
rect 23799 39797 23811 39831
rect 23753 39791 23811 39797
rect 24486 39788 24492 39840
rect 24544 39828 24550 39840
rect 24872 39837 24900 39868
rect 24673 39831 24731 39837
rect 24673 39828 24685 39831
rect 24544 39800 24685 39828
rect 24544 39788 24550 39800
rect 24673 39797 24685 39800
rect 24719 39797 24731 39831
rect 24673 39791 24731 39797
rect 24857 39831 24915 39837
rect 24857 39797 24869 39831
rect 24903 39797 24915 39831
rect 24857 39791 24915 39797
rect 24946 39788 24952 39840
rect 25004 39828 25010 39840
rect 25148 39828 25176 39868
rect 25593 39865 25605 39868
rect 25639 39865 25651 39899
rect 27080 39896 27108 39924
rect 27338 39896 27344 39908
rect 27080 39868 27344 39896
rect 25593 39859 25651 39865
rect 27338 39856 27344 39868
rect 27396 39856 27402 39908
rect 28074 39856 28080 39908
rect 28132 39896 28138 39908
rect 31662 39896 31668 39908
rect 28132 39868 31668 39896
rect 28132 39856 28138 39868
rect 31662 39856 31668 39868
rect 31720 39856 31726 39908
rect 25498 39828 25504 39840
rect 25004 39800 25176 39828
rect 25459 39800 25504 39828
rect 25004 39788 25010 39800
rect 25498 39788 25504 39800
rect 25556 39788 25562 39840
rect 27154 39828 27160 39840
rect 27115 39800 27160 39828
rect 27154 39788 27160 39800
rect 27212 39788 27218 39840
rect 33226 39788 33232 39840
rect 33284 39828 33290 39840
rect 33321 39831 33379 39837
rect 33321 39828 33333 39831
rect 33284 39800 33333 39828
rect 33284 39788 33290 39800
rect 33321 39797 33333 39800
rect 33367 39797 33379 39831
rect 35360 39828 35388 40072
rect 35529 40035 35587 40041
rect 35529 40001 35541 40035
rect 35575 40001 35587 40035
rect 35529 39995 35587 40001
rect 35713 40035 35771 40041
rect 35713 40001 35725 40035
rect 35759 40001 35771 40035
rect 35820 40032 35848 40140
rect 39390 40128 39396 40140
rect 39448 40128 39454 40180
rect 40034 40128 40040 40180
rect 40092 40168 40098 40180
rect 40402 40168 40408 40180
rect 40092 40140 40408 40168
rect 40092 40128 40098 40140
rect 40402 40128 40408 40140
rect 40460 40168 40466 40180
rect 40497 40171 40555 40177
rect 40497 40168 40509 40171
rect 40460 40140 40509 40168
rect 40460 40128 40466 40140
rect 40497 40137 40509 40140
rect 40543 40168 40555 40171
rect 41046 40168 41052 40180
rect 40543 40140 41052 40168
rect 40543 40137 40555 40140
rect 40497 40131 40555 40137
rect 41046 40128 41052 40140
rect 41104 40128 41110 40180
rect 37568 40072 38332 40100
rect 37568 40044 37596 40072
rect 36170 40032 36176 40044
rect 35820 40004 36176 40032
rect 35713 39995 35771 40001
rect 35544 39896 35572 39995
rect 35728 39964 35756 39995
rect 36170 39992 36176 40004
rect 36228 39992 36234 40044
rect 36354 40032 36360 40044
rect 36315 40004 36360 40032
rect 36354 39992 36360 40004
rect 36412 39992 36418 40044
rect 37461 40035 37519 40041
rect 37461 40001 37473 40035
rect 37507 40032 37519 40035
rect 37550 40032 37556 40044
rect 37507 40004 37556 40032
rect 37507 40001 37519 40004
rect 37461 39995 37519 40001
rect 37550 39992 37556 40004
rect 37608 39992 37614 40044
rect 37645 40035 37703 40041
rect 37645 40001 37657 40035
rect 37691 40032 37703 40035
rect 38102 40032 38108 40044
rect 37691 40004 38108 40032
rect 37691 40001 37703 40004
rect 37645 39995 37703 40001
rect 38102 39992 38108 40004
rect 38160 39992 38166 40044
rect 38304 40041 38332 40072
rect 38654 40060 38660 40112
rect 38712 40100 38718 40112
rect 38712 40072 39804 40100
rect 38712 40060 38718 40072
rect 38289 40035 38347 40041
rect 38289 40001 38301 40035
rect 38335 40001 38347 40035
rect 38289 39995 38347 40001
rect 38565 40035 38623 40041
rect 38565 40001 38577 40035
rect 38611 40032 38623 40035
rect 38930 40032 38936 40044
rect 38611 40004 38700 40032
rect 38843 40004 38936 40032
rect 38611 40001 38623 40004
rect 38565 39995 38623 40001
rect 38672 39976 38700 40004
rect 38930 39992 38936 40004
rect 38988 40032 38994 40044
rect 39666 40032 39672 40044
rect 38988 40004 39528 40032
rect 39627 40004 39672 40032
rect 38988 39992 38994 40004
rect 36265 39967 36323 39973
rect 36265 39964 36277 39967
rect 35728 39936 36277 39964
rect 36265 39933 36277 39936
rect 36311 39933 36323 39967
rect 36265 39927 36323 39933
rect 38654 39924 38660 39976
rect 38712 39924 38718 39976
rect 39500 39964 39528 40004
rect 39666 39992 39672 40004
rect 39724 39992 39730 40044
rect 39776 40041 39804 40072
rect 39761 40035 39819 40041
rect 39761 40001 39773 40035
rect 39807 40001 39819 40035
rect 39761 39995 39819 40001
rect 39850 39992 39856 40044
rect 39908 40032 39914 40044
rect 40037 40035 40095 40041
rect 39908 40004 39953 40032
rect 39908 39992 39914 40004
rect 40037 40001 40049 40035
rect 40083 40032 40095 40035
rect 52917 40035 52975 40041
rect 40083 40004 49556 40032
rect 40083 40001 40095 40004
rect 40037 39995 40095 40001
rect 40052 39964 40080 39995
rect 39500 39936 40080 39964
rect 41046 39924 41052 39976
rect 41104 39964 41110 39976
rect 49528 39964 49556 40004
rect 52917 40001 52929 40035
rect 52963 40032 52975 40035
rect 53558 40032 53564 40044
rect 52963 40004 53564 40032
rect 52963 40001 52975 40004
rect 52917 39995 52975 40001
rect 53558 39992 53564 40004
rect 53616 39992 53622 40044
rect 53377 39967 53435 39973
rect 53377 39964 53389 39967
rect 41104 39936 45554 39964
rect 49528 39936 53389 39964
rect 41104 39924 41110 39936
rect 35802 39896 35808 39908
rect 35544 39868 35808 39896
rect 35802 39856 35808 39868
rect 35860 39856 35866 39908
rect 38286 39896 38292 39908
rect 38247 39868 38292 39896
rect 38286 39856 38292 39868
rect 38344 39856 38350 39908
rect 39850 39856 39856 39908
rect 39908 39896 39914 39908
rect 41601 39899 41659 39905
rect 41601 39896 41613 39899
rect 39908 39868 41613 39896
rect 39908 39856 39914 39868
rect 41601 39865 41613 39868
rect 41647 39865 41659 39899
rect 45526 39896 45554 39936
rect 53377 39933 53389 39936
rect 53423 39933 53435 39967
rect 53377 39927 53435 39933
rect 52822 39896 52828 39908
rect 45526 39868 52828 39896
rect 41601 39859 41659 39865
rect 52822 39856 52828 39868
rect 52880 39856 52886 39908
rect 35618 39828 35624 39840
rect 35360 39800 35624 39828
rect 33321 39791 33379 39797
rect 35618 39788 35624 39800
rect 35676 39828 35682 39840
rect 35713 39831 35771 39837
rect 35713 39828 35725 39831
rect 35676 39800 35725 39828
rect 35676 39788 35682 39800
rect 35713 39797 35725 39800
rect 35759 39797 35771 39831
rect 35713 39791 35771 39797
rect 37458 39788 37464 39840
rect 37516 39828 37522 39840
rect 37553 39831 37611 39837
rect 37553 39828 37565 39831
rect 37516 39800 37565 39828
rect 37516 39788 37522 39800
rect 37553 39797 37565 39800
rect 37599 39797 37611 39831
rect 37553 39791 37611 39797
rect 1104 39738 54372 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 54372 39738
rect 1104 39664 54372 39686
rect 21174 39624 21180 39636
rect 18616 39596 21180 39624
rect 18616 39565 18644 39596
rect 21174 39584 21180 39596
rect 21232 39584 21238 39636
rect 21361 39627 21419 39633
rect 21361 39593 21373 39627
rect 21407 39624 21419 39627
rect 22186 39624 22192 39636
rect 21407 39596 22192 39624
rect 21407 39593 21419 39596
rect 21361 39587 21419 39593
rect 22186 39584 22192 39596
rect 22244 39584 22250 39636
rect 22370 39624 22376 39636
rect 22331 39596 22376 39624
rect 22370 39584 22376 39596
rect 22428 39584 22434 39636
rect 22462 39584 22468 39636
rect 22520 39624 22526 39636
rect 23658 39624 23664 39636
rect 22520 39596 23664 39624
rect 22520 39584 22526 39596
rect 23658 39584 23664 39596
rect 23716 39624 23722 39636
rect 26878 39624 26884 39636
rect 23716 39596 26884 39624
rect 23716 39584 23722 39596
rect 26878 39584 26884 39596
rect 26936 39584 26942 39636
rect 31478 39584 31484 39636
rect 31536 39624 31542 39636
rect 31573 39627 31631 39633
rect 31573 39624 31585 39627
rect 31536 39596 31585 39624
rect 31536 39584 31542 39596
rect 31573 39593 31585 39596
rect 31619 39593 31631 39627
rect 32674 39624 32680 39636
rect 32635 39596 32680 39624
rect 31573 39587 31631 39593
rect 32674 39584 32680 39596
rect 32732 39624 32738 39636
rect 33134 39624 33140 39636
rect 32732 39596 33140 39624
rect 32732 39584 32738 39596
rect 33134 39584 33140 39596
rect 33192 39584 33198 39636
rect 33318 39584 33324 39636
rect 33376 39624 33382 39636
rect 33778 39624 33784 39636
rect 33376 39596 33784 39624
rect 33376 39584 33382 39596
rect 33778 39584 33784 39596
rect 33836 39584 33842 39636
rect 34146 39584 34152 39636
rect 34204 39624 34210 39636
rect 35342 39624 35348 39636
rect 34204 39596 35348 39624
rect 34204 39584 34210 39596
rect 35342 39584 35348 39596
rect 35400 39624 35406 39636
rect 38562 39624 38568 39636
rect 35400 39596 38568 39624
rect 35400 39584 35406 39596
rect 38562 39584 38568 39596
rect 38620 39584 38626 39636
rect 41506 39624 41512 39636
rect 41467 39596 41512 39624
rect 41506 39584 41512 39596
rect 41564 39584 41570 39636
rect 18601 39559 18659 39565
rect 18601 39556 18613 39559
rect 16546 39528 18613 39556
rect 15470 39448 15476 39500
rect 15528 39488 15534 39500
rect 16546 39488 16574 39528
rect 18601 39525 18613 39528
rect 18647 39525 18659 39559
rect 18601 39519 18659 39525
rect 19981 39559 20039 39565
rect 19981 39525 19993 39559
rect 20027 39525 20039 39559
rect 19981 39519 20039 39525
rect 15528 39460 16574 39488
rect 17681 39491 17739 39497
rect 15528 39448 15534 39460
rect 16132 39429 16160 39460
rect 17681 39457 17693 39491
rect 17727 39488 17739 39491
rect 18046 39488 18052 39500
rect 17727 39460 18052 39488
rect 17727 39457 17739 39460
rect 17681 39451 17739 39457
rect 18046 39448 18052 39460
rect 18104 39448 18110 39500
rect 18141 39491 18199 39497
rect 18141 39457 18153 39491
rect 18187 39488 18199 39491
rect 18782 39488 18788 39500
rect 18187 39460 18788 39488
rect 18187 39457 18199 39460
rect 18141 39451 18199 39457
rect 18782 39448 18788 39460
rect 18840 39448 18846 39500
rect 19996 39488 20024 39519
rect 19996 39460 20668 39488
rect 15933 39423 15991 39429
rect 15933 39389 15945 39423
rect 15979 39389 15991 39423
rect 15933 39383 15991 39389
rect 16117 39423 16175 39429
rect 16117 39389 16129 39423
rect 16163 39389 16175 39423
rect 16758 39420 16764 39432
rect 16719 39392 16764 39420
rect 16117 39383 16175 39389
rect 14921 39355 14979 39361
rect 14921 39321 14933 39355
rect 14967 39352 14979 39355
rect 15948 39352 15976 39383
rect 16758 39380 16764 39392
rect 16816 39380 16822 39432
rect 16942 39420 16948 39432
rect 16903 39392 16948 39420
rect 16942 39380 16948 39392
rect 17000 39380 17006 39432
rect 17037 39423 17095 39429
rect 17037 39389 17049 39423
rect 17083 39420 17095 39423
rect 17310 39420 17316 39432
rect 17083 39392 17316 39420
rect 17083 39389 17095 39392
rect 17037 39383 17095 39389
rect 17310 39380 17316 39392
rect 17368 39380 17374 39432
rect 17770 39380 17776 39432
rect 17828 39420 17834 39432
rect 17828 39392 17873 39420
rect 17828 39380 17834 39392
rect 19334 39380 19340 39432
rect 19392 39420 19398 39432
rect 19705 39423 19763 39429
rect 19705 39420 19717 39423
rect 19392 39392 19717 39420
rect 19392 39380 19398 39392
rect 19705 39389 19717 39392
rect 19751 39389 19763 39423
rect 20438 39420 20444 39432
rect 20399 39392 20444 39420
rect 19705 39383 19763 39389
rect 20438 39380 20444 39392
rect 20496 39380 20502 39432
rect 20640 39429 20668 39460
rect 20625 39423 20683 39429
rect 20625 39389 20637 39423
rect 20671 39389 20683 39423
rect 20625 39383 20683 39389
rect 16298 39352 16304 39364
rect 14967 39324 16304 39352
rect 14967 39321 14979 39324
rect 14921 39315 14979 39321
rect 16298 39312 16304 39324
rect 16356 39312 16362 39364
rect 16577 39355 16635 39361
rect 16577 39321 16589 39355
rect 16623 39352 16635 39355
rect 17402 39352 17408 39364
rect 16623 39324 17408 39352
rect 16623 39321 16635 39324
rect 16577 39315 16635 39321
rect 17402 39312 17408 39324
rect 17460 39312 17466 39364
rect 19981 39355 20039 39361
rect 19981 39321 19993 39355
rect 20027 39352 20039 39355
rect 20806 39352 20812 39364
rect 20027 39324 20812 39352
rect 20027 39321 20039 39324
rect 19981 39315 20039 39321
rect 20806 39312 20812 39324
rect 20864 39312 20870 39364
rect 21192 39352 21220 39584
rect 23569 39559 23627 39565
rect 23569 39525 23581 39559
rect 23615 39556 23627 39559
rect 25498 39556 25504 39568
rect 23615 39528 25504 39556
rect 23615 39525 23627 39528
rect 23569 39519 23627 39525
rect 25498 39516 25504 39528
rect 25556 39516 25562 39568
rect 26513 39559 26571 39565
rect 26513 39525 26525 39559
rect 26559 39525 26571 39559
rect 26513 39519 26571 39525
rect 23474 39488 23480 39500
rect 23435 39460 23480 39488
rect 23474 39448 23480 39460
rect 23532 39448 23538 39500
rect 23845 39491 23903 39497
rect 23845 39457 23857 39491
rect 23891 39488 23903 39491
rect 23891 39460 26280 39488
rect 23891 39457 23903 39460
rect 23845 39451 23903 39457
rect 22370 39380 22376 39432
rect 22428 39420 22434 39432
rect 23201 39423 23259 39429
rect 23201 39420 23213 39423
rect 22428 39392 23213 39420
rect 22428 39380 22434 39392
rect 23201 39389 23213 39392
rect 23247 39389 23259 39423
rect 23201 39383 23259 39389
rect 23385 39423 23443 39429
rect 23385 39389 23397 39423
rect 23431 39389 23443 39423
rect 23658 39420 23664 39432
rect 23619 39392 23664 39420
rect 23385 39383 23443 39389
rect 22554 39352 22560 39364
rect 21192 39324 22560 39352
rect 22554 39312 22560 39324
rect 22612 39312 22618 39364
rect 22738 39312 22744 39364
rect 22796 39352 22802 39364
rect 22796 39324 22889 39352
rect 22796 39312 22802 39324
rect 23106 39312 23112 39364
rect 23164 39352 23170 39364
rect 23400 39352 23428 39383
rect 23658 39380 23664 39392
rect 23716 39380 23722 39432
rect 23750 39380 23756 39432
rect 23808 39420 23814 39432
rect 24397 39423 24455 39429
rect 24397 39420 24409 39423
rect 23808 39392 24409 39420
rect 23808 39380 23814 39392
rect 24397 39389 24409 39392
rect 24443 39389 24455 39423
rect 24397 39383 24455 39389
rect 24486 39380 24492 39432
rect 24544 39420 24550 39432
rect 24581 39423 24639 39429
rect 24581 39420 24593 39423
rect 24544 39392 24593 39420
rect 24544 39380 24550 39392
rect 24581 39389 24593 39392
rect 24627 39389 24639 39423
rect 24581 39383 24639 39389
rect 24673 39423 24731 39429
rect 24673 39389 24685 39423
rect 24719 39389 24731 39423
rect 24673 39383 24731 39389
rect 24765 39423 24823 39429
rect 24765 39389 24777 39423
rect 24811 39420 24823 39423
rect 24854 39420 24860 39432
rect 24811 39392 24860 39420
rect 24811 39389 24823 39392
rect 24765 39383 24823 39389
rect 23164 39324 23428 39352
rect 23164 39312 23170 39324
rect 15470 39284 15476 39296
rect 15431 39256 15476 39284
rect 15470 39244 15476 39256
rect 15528 39244 15534 39296
rect 15930 39244 15936 39296
rect 15988 39284 15994 39296
rect 16025 39287 16083 39293
rect 16025 39284 16037 39287
rect 15988 39256 16037 39284
rect 15988 39244 15994 39256
rect 16025 39253 16037 39256
rect 16071 39253 16083 39287
rect 17494 39284 17500 39296
rect 17455 39256 17500 39284
rect 16025 39247 16083 39253
rect 17494 39244 17500 39256
rect 17552 39244 17558 39296
rect 19426 39244 19432 39296
rect 19484 39284 19490 39296
rect 19797 39287 19855 39293
rect 19797 39284 19809 39287
rect 19484 39256 19809 39284
rect 19484 39244 19490 39256
rect 19797 39253 19809 39256
rect 19843 39253 19855 39287
rect 19797 39247 19855 39253
rect 20533 39287 20591 39293
rect 20533 39253 20545 39287
rect 20579 39284 20591 39287
rect 20714 39284 20720 39296
rect 20579 39256 20720 39284
rect 20579 39253 20591 39256
rect 20533 39247 20591 39253
rect 20714 39244 20720 39256
rect 20772 39244 20778 39296
rect 21913 39287 21971 39293
rect 21913 39253 21925 39287
rect 21959 39284 21971 39287
rect 22462 39284 22468 39296
rect 21959 39256 22468 39284
rect 21959 39253 21971 39256
rect 21913 39247 21971 39253
rect 22462 39244 22468 39256
rect 22520 39244 22526 39296
rect 22756 39284 22784 39312
rect 23290 39284 23296 39296
rect 22756 39256 23296 39284
rect 23290 39244 23296 39256
rect 23348 39244 23354 39296
rect 24302 39244 24308 39296
rect 24360 39284 24366 39296
rect 24688 39284 24716 39383
rect 24854 39380 24860 39392
rect 24912 39380 24918 39432
rect 24946 39380 24952 39432
rect 25004 39420 25010 39432
rect 26252 39429 26280 39460
rect 26237 39423 26295 39429
rect 25004 39392 25049 39420
rect 25004 39380 25010 39392
rect 26237 39389 26249 39423
rect 26283 39389 26295 39423
rect 26528 39420 26556 39519
rect 30834 39516 30840 39568
rect 30892 39556 30898 39568
rect 30892 39528 31754 39556
rect 30892 39516 30898 39528
rect 26970 39488 26976 39500
rect 26931 39460 26976 39488
rect 26970 39448 26976 39460
rect 27028 39448 27034 39500
rect 29733 39491 29791 39497
rect 29733 39457 29745 39491
rect 29779 39488 29791 39491
rect 30285 39491 30343 39497
rect 30285 39488 30297 39491
rect 29779 39460 30297 39488
rect 29779 39457 29791 39460
rect 29733 39451 29791 39457
rect 30285 39457 30297 39460
rect 30331 39457 30343 39491
rect 31110 39488 31116 39500
rect 30285 39451 30343 39457
rect 30677 39460 31116 39488
rect 27249 39423 27307 39429
rect 27249 39420 27261 39423
rect 26528 39392 27261 39420
rect 26237 39383 26295 39389
rect 27249 39389 27261 39392
rect 27295 39389 27307 39423
rect 27249 39383 27307 39389
rect 29825 39423 29883 39429
rect 29825 39389 29837 39423
rect 29871 39420 29883 39423
rect 30677 39420 30705 39460
rect 31110 39448 31116 39460
rect 31168 39448 31174 39500
rect 31726 39488 31754 39528
rect 34422 39516 34428 39568
rect 34480 39556 34486 39568
rect 34977 39559 35035 39565
rect 34977 39556 34989 39559
rect 34480 39528 34989 39556
rect 34480 39516 34486 39528
rect 34977 39525 34989 39528
rect 35023 39525 35035 39559
rect 39853 39559 39911 39565
rect 39853 39556 39865 39559
rect 34977 39519 35035 39525
rect 36556 39528 39865 39556
rect 31726 39460 31800 39488
rect 29871 39392 30705 39420
rect 29871 39389 29883 39392
rect 29825 39383 29883 39389
rect 30742 39380 30748 39432
rect 30800 39420 30806 39432
rect 30800 39392 30880 39420
rect 30800 39380 30806 39392
rect 25777 39355 25835 39361
rect 25777 39321 25789 39355
rect 25823 39352 25835 39355
rect 26418 39352 26424 39364
rect 25823 39324 26424 39352
rect 25823 39321 25835 39324
rect 25777 39315 25835 39321
rect 26418 39312 26424 39324
rect 26476 39312 26482 39364
rect 26510 39312 26516 39364
rect 26568 39352 26574 39364
rect 26568 39324 26613 39352
rect 26568 39312 26574 39324
rect 29914 39312 29920 39364
rect 29972 39352 29978 39364
rect 30423 39355 30481 39361
rect 30423 39352 30435 39355
rect 29972 39324 30435 39352
rect 29972 39312 29978 39324
rect 30423 39321 30435 39324
rect 30469 39321 30481 39355
rect 30423 39315 30481 39321
rect 30561 39355 30619 39361
rect 30561 39321 30573 39355
rect 30607 39321 30619 39355
rect 30561 39315 30619 39321
rect 25130 39284 25136 39296
rect 24360 39256 24716 39284
rect 25091 39256 25136 39284
rect 24360 39244 24366 39256
rect 25130 39244 25136 39256
rect 25188 39244 25194 39296
rect 26326 39284 26332 39296
rect 26287 39256 26332 39284
rect 26326 39244 26332 39256
rect 26384 39244 26390 39296
rect 27246 39244 27252 39296
rect 27304 39284 27310 39296
rect 28353 39287 28411 39293
rect 28353 39284 28365 39287
rect 27304 39256 28365 39284
rect 27304 39244 27310 39256
rect 28353 39253 28365 39256
rect 28399 39253 28411 39287
rect 30576 39284 30604 39315
rect 30650 39312 30656 39364
rect 30708 39352 30714 39364
rect 30852 39352 30880 39392
rect 31772 39361 31800 39460
rect 32582 39448 32588 39500
rect 32640 39488 32646 39500
rect 33318 39488 33324 39500
rect 32640 39460 33324 39488
rect 32640 39448 32646 39460
rect 33318 39448 33324 39460
rect 33376 39448 33382 39500
rect 35342 39488 35348 39500
rect 34716 39460 35348 39488
rect 33410 39380 33416 39432
rect 33468 39420 33474 39432
rect 34716 39429 34744 39460
rect 35342 39448 35348 39460
rect 35400 39488 35406 39500
rect 35529 39491 35587 39497
rect 35529 39488 35541 39491
rect 35400 39460 35541 39488
rect 35400 39448 35406 39460
rect 35529 39457 35541 39460
rect 35575 39457 35587 39491
rect 35529 39451 35587 39457
rect 36170 39448 36176 39500
rect 36228 39488 36234 39500
rect 36556 39497 36584 39528
rect 39853 39525 39865 39528
rect 39899 39556 39911 39559
rect 40034 39556 40040 39568
rect 39899 39528 40040 39556
rect 39899 39525 39911 39528
rect 39853 39519 39911 39525
rect 40034 39516 40040 39528
rect 40092 39516 40098 39568
rect 36541 39491 36599 39497
rect 36541 39488 36553 39491
rect 36228 39460 36553 39488
rect 36228 39448 36234 39460
rect 36541 39457 36553 39460
rect 36587 39457 36599 39491
rect 36541 39451 36599 39457
rect 38286 39448 38292 39500
rect 38344 39488 38350 39500
rect 38381 39491 38439 39497
rect 38381 39488 38393 39491
rect 38344 39460 38393 39488
rect 38344 39448 38350 39460
rect 38381 39457 38393 39460
rect 38427 39457 38439 39491
rect 38381 39451 38439 39457
rect 34701 39423 34759 39429
rect 34701 39420 34713 39423
rect 33468 39392 34713 39420
rect 33468 39380 33474 39392
rect 34701 39389 34713 39392
rect 34747 39389 34759 39423
rect 34701 39383 34759 39389
rect 34790 39380 34796 39432
rect 34848 39420 34854 39432
rect 35250 39420 35256 39432
rect 34848 39392 35256 39420
rect 34848 39380 34854 39392
rect 35250 39380 35256 39392
rect 35308 39420 35314 39432
rect 35437 39423 35495 39429
rect 35437 39420 35449 39423
rect 35308 39392 35449 39420
rect 35308 39380 35314 39392
rect 35437 39389 35449 39392
rect 35483 39389 35495 39423
rect 35618 39420 35624 39432
rect 35579 39392 35624 39420
rect 35437 39383 35495 39389
rect 35618 39380 35624 39392
rect 35676 39380 35682 39432
rect 36354 39420 36360 39432
rect 36315 39392 36360 39420
rect 36354 39380 36360 39392
rect 36412 39380 36418 39432
rect 37366 39380 37372 39432
rect 37424 39420 37430 39432
rect 37461 39423 37519 39429
rect 37461 39420 37473 39423
rect 37424 39392 37473 39420
rect 37424 39380 37430 39392
rect 37461 39389 37473 39392
rect 37507 39389 37519 39423
rect 37461 39383 37519 39389
rect 37550 39380 37556 39432
rect 37608 39420 37614 39432
rect 37737 39423 37795 39429
rect 37737 39420 37749 39423
rect 37608 39392 37749 39420
rect 37608 39380 37614 39392
rect 37737 39389 37749 39392
rect 37783 39389 37795 39423
rect 38470 39420 38476 39432
rect 38431 39392 38476 39420
rect 37737 39383 37795 39389
rect 38470 39380 38476 39392
rect 38528 39380 38534 39432
rect 31541 39355 31599 39361
rect 31541 39352 31553 39355
rect 30708 39324 30753 39352
rect 30852 39324 31553 39352
rect 30708 39312 30714 39324
rect 31541 39321 31553 39324
rect 31587 39321 31599 39355
rect 31541 39315 31599 39321
rect 31757 39355 31815 39361
rect 31757 39321 31769 39355
rect 31803 39321 31815 39355
rect 31757 39315 31815 39321
rect 32950 39312 32956 39364
rect 33008 39352 33014 39364
rect 33289 39355 33347 39361
rect 33289 39352 33301 39355
rect 33008 39324 33301 39352
rect 33008 39312 33014 39324
rect 33289 39321 33301 39324
rect 33335 39321 33347 39355
rect 33502 39352 33508 39364
rect 33463 39324 33508 39352
rect 33289 39315 33347 39321
rect 33502 39312 33508 39324
rect 33560 39312 33566 39364
rect 34974 39352 34980 39364
rect 34935 39324 34980 39352
rect 34974 39312 34980 39324
rect 35032 39312 35038 39364
rect 37645 39355 37703 39361
rect 37645 39321 37657 39355
rect 37691 39352 37703 39355
rect 38194 39352 38200 39364
rect 37691 39324 38200 39352
rect 37691 39321 37703 39324
rect 37645 39315 37703 39321
rect 38194 39312 38200 39324
rect 38252 39312 38258 39364
rect 39850 39312 39856 39364
rect 39908 39352 39914 39364
rect 40957 39355 41015 39361
rect 40957 39352 40969 39355
rect 39908 39324 40969 39352
rect 39908 39312 39914 39324
rect 40957 39321 40969 39324
rect 41003 39321 41015 39355
rect 40957 39315 41015 39321
rect 30834 39284 30840 39296
rect 30576 39256 30840 39284
rect 28353 39247 28411 39253
rect 30834 39244 30840 39256
rect 30892 39244 30898 39296
rect 30929 39287 30987 39293
rect 30929 39253 30941 39287
rect 30975 39284 30987 39287
rect 31018 39284 31024 39296
rect 30975 39256 31024 39284
rect 30975 39253 30987 39256
rect 30929 39247 30987 39253
rect 31018 39244 31024 39256
rect 31076 39244 31082 39296
rect 31386 39284 31392 39296
rect 31347 39256 31392 39284
rect 31386 39244 31392 39256
rect 31444 39244 31450 39296
rect 33042 39244 33048 39296
rect 33100 39284 33106 39296
rect 33137 39287 33195 39293
rect 33137 39284 33149 39287
rect 33100 39256 33149 39284
rect 33100 39244 33106 39256
rect 33137 39253 33149 39256
rect 33183 39253 33195 39287
rect 33137 39247 33195 39253
rect 33778 39244 33784 39296
rect 33836 39284 33842 39296
rect 33965 39287 34023 39293
rect 33965 39284 33977 39287
rect 33836 39256 33977 39284
rect 33836 39244 33842 39256
rect 33965 39253 33977 39256
rect 34011 39253 34023 39287
rect 33965 39247 34023 39253
rect 34698 39244 34704 39296
rect 34756 39284 34762 39296
rect 34793 39287 34851 39293
rect 34793 39284 34805 39287
rect 34756 39256 34805 39284
rect 34756 39244 34762 39256
rect 34793 39253 34805 39256
rect 34839 39253 34851 39287
rect 34793 39247 34851 39253
rect 35802 39244 35808 39296
rect 35860 39284 35866 39296
rect 36173 39287 36231 39293
rect 36173 39284 36185 39287
rect 35860 39256 36185 39284
rect 35860 39244 35866 39256
rect 36173 39253 36185 39256
rect 36219 39253 36231 39287
rect 37274 39284 37280 39296
rect 37235 39256 37280 39284
rect 36173 39247 36231 39253
rect 37274 39244 37280 39256
rect 37332 39244 37338 39296
rect 39022 39244 39028 39296
rect 39080 39284 39086 39296
rect 39301 39287 39359 39293
rect 39301 39284 39313 39287
rect 39080 39256 39313 39284
rect 39080 39244 39086 39256
rect 39301 39253 39313 39256
rect 39347 39253 39359 39287
rect 40402 39284 40408 39296
rect 40363 39256 40408 39284
rect 39301 39247 39359 39253
rect 40402 39244 40408 39256
rect 40460 39244 40466 39296
rect 1104 39194 54372 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 54372 39194
rect 1104 39120 54372 39142
rect 15930 39040 15936 39092
rect 15988 39080 15994 39092
rect 17589 39083 17647 39089
rect 17589 39080 17601 39083
rect 15988 39052 17601 39080
rect 15988 39040 15994 39052
rect 17589 39049 17601 39052
rect 17635 39080 17647 39083
rect 17770 39080 17776 39092
rect 17635 39052 17776 39080
rect 17635 39049 17647 39052
rect 17589 39043 17647 39049
rect 17770 39040 17776 39052
rect 17828 39040 17834 39092
rect 17957 39083 18015 39089
rect 17957 39049 17969 39083
rect 18003 39080 18015 39083
rect 19334 39080 19340 39092
rect 18003 39052 19340 39080
rect 18003 39049 18015 39052
rect 17957 39043 18015 39049
rect 19334 39040 19340 39052
rect 19392 39080 19398 39092
rect 20162 39080 20168 39092
rect 19392 39052 20040 39080
rect 20075 39052 20168 39080
rect 19392 39040 19398 39052
rect 16025 39015 16083 39021
rect 16025 38981 16037 39015
rect 16071 39012 16083 39015
rect 16758 39012 16764 39024
rect 16071 38984 16764 39012
rect 16071 38981 16083 38984
rect 16025 38975 16083 38981
rect 16758 38972 16764 38984
rect 16816 39012 16822 39024
rect 16853 39015 16911 39021
rect 16853 39012 16865 39015
rect 16816 38984 16865 39012
rect 16816 38972 16822 38984
rect 16853 38981 16865 38984
rect 16899 38981 16911 39015
rect 16853 38975 16911 38981
rect 17037 39015 17095 39021
rect 17037 38981 17049 39015
rect 17083 39012 17095 39015
rect 17788 39012 17816 39040
rect 18690 39012 18696 39024
rect 17083 38984 17724 39012
rect 17788 38984 18460 39012
rect 18651 38984 18696 39012
rect 17083 38981 17095 38984
rect 17037 38975 17095 38981
rect 1578 38904 1584 38956
rect 1636 38944 1642 38956
rect 1857 38947 1915 38953
rect 1857 38944 1869 38947
rect 1636 38916 1869 38944
rect 1636 38904 1642 38916
rect 1857 38913 1869 38916
rect 1903 38913 1915 38947
rect 15930 38944 15936 38956
rect 15891 38916 15936 38944
rect 1857 38907 1915 38913
rect 15930 38904 15936 38916
rect 15988 38904 15994 38956
rect 16117 38947 16175 38953
rect 16117 38913 16129 38947
rect 16163 38944 16175 38947
rect 16666 38944 16672 38956
rect 16163 38916 16672 38944
rect 16163 38913 16175 38916
rect 16117 38907 16175 38913
rect 16666 38904 16672 38916
rect 16724 38904 16730 38956
rect 17402 38904 17408 38956
rect 17460 38944 17466 38956
rect 17497 38947 17555 38953
rect 17497 38944 17509 38947
rect 17460 38916 17509 38944
rect 17460 38904 17466 38916
rect 17497 38913 17509 38916
rect 17543 38913 17555 38947
rect 17696 38944 17724 38984
rect 17773 38947 17831 38953
rect 17773 38944 17785 38947
rect 17696 38916 17785 38944
rect 17497 38907 17555 38913
rect 17773 38913 17785 38916
rect 17819 38944 17831 38947
rect 18322 38944 18328 38956
rect 17819 38916 18328 38944
rect 17819 38913 17831 38916
rect 17773 38907 17831 38913
rect 17512 38876 17540 38907
rect 18322 38904 18328 38916
rect 18380 38904 18386 38956
rect 18432 38953 18460 38984
rect 18690 38972 18696 38984
rect 18748 38972 18754 39024
rect 20012 39021 20040 39052
rect 20162 39040 20168 39052
rect 20220 39080 20226 39092
rect 20438 39080 20444 39092
rect 20220 39052 20444 39080
rect 20220 39040 20226 39052
rect 20438 39040 20444 39052
rect 20496 39040 20502 39092
rect 20622 39080 20628 39092
rect 20583 39052 20628 39080
rect 20622 39040 20628 39052
rect 20680 39040 20686 39092
rect 22370 39080 22376 39092
rect 22331 39052 22376 39080
rect 22370 39040 22376 39052
rect 22428 39040 22434 39092
rect 22830 39040 22836 39092
rect 22888 39080 22894 39092
rect 23201 39083 23259 39089
rect 23201 39080 23213 39083
rect 22888 39052 23213 39080
rect 22888 39040 22894 39052
rect 23201 39049 23213 39052
rect 23247 39049 23259 39083
rect 23201 39043 23259 39049
rect 19797 39015 19855 39021
rect 19797 38981 19809 39015
rect 19843 38981 19855 39015
rect 19797 38975 19855 38981
rect 19997 39015 20055 39021
rect 19997 38981 20009 39015
rect 20043 38981 20055 39015
rect 19997 38975 20055 38981
rect 18417 38947 18475 38953
rect 18417 38913 18429 38947
rect 18463 38913 18475 38947
rect 18417 38907 18475 38913
rect 18509 38947 18567 38953
rect 18509 38913 18521 38947
rect 18555 38913 18567 38947
rect 19812 38944 19840 38975
rect 20714 38972 20720 39024
rect 20772 39012 20778 39024
rect 23216 39012 23244 39043
rect 23750 39040 23756 39092
rect 23808 39080 23814 39092
rect 23845 39083 23903 39089
rect 23845 39080 23857 39083
rect 23808 39052 23857 39080
rect 23808 39040 23814 39052
rect 23845 39049 23857 39052
rect 23891 39049 23903 39083
rect 23845 39043 23903 39049
rect 24765 39083 24823 39089
rect 24765 39049 24777 39083
rect 24811 39080 24823 39083
rect 25317 39083 25375 39089
rect 24811 39052 25268 39080
rect 24811 39049 24823 39052
rect 24765 39043 24823 39049
rect 24946 39012 24952 39024
rect 20772 38984 22048 39012
rect 23216 38984 24952 39012
rect 20772 38972 20778 38984
rect 22020 38956 22048 38984
rect 24946 38972 24952 38984
rect 25004 38972 25010 39024
rect 25240 39012 25268 39052
rect 25317 39049 25329 39083
rect 25363 39080 25375 39083
rect 26234 39080 26240 39092
rect 25363 39052 26240 39080
rect 25363 39049 25375 39052
rect 25317 39043 25375 39049
rect 26234 39040 26240 39052
rect 26292 39040 26298 39092
rect 26326 39040 26332 39092
rect 26384 39080 26390 39092
rect 26973 39083 27031 39089
rect 26973 39080 26985 39083
rect 26384 39052 26985 39080
rect 26384 39040 26390 39052
rect 26973 39049 26985 39052
rect 27019 39049 27031 39083
rect 26973 39043 27031 39049
rect 28997 39083 29055 39089
rect 28997 39049 29009 39083
rect 29043 39080 29055 39083
rect 29546 39080 29552 39092
rect 29043 39052 29552 39080
rect 29043 39049 29055 39052
rect 28997 39043 29055 39049
rect 29546 39040 29552 39052
rect 29604 39040 29610 39092
rect 29914 39080 29920 39092
rect 29875 39052 29920 39080
rect 29914 39040 29920 39052
rect 29972 39040 29978 39092
rect 35069 39083 35127 39089
rect 30576 39052 33364 39080
rect 26510 39012 26516 39024
rect 25240 38984 26516 39012
rect 26510 38972 26516 38984
rect 26568 38972 26574 39024
rect 30576 39012 30604 39052
rect 31386 39012 31392 39024
rect 26620 38984 30604 39012
rect 30668 38984 31392 39012
rect 20806 38944 20812 38956
rect 19812 38916 20812 38944
rect 18509 38907 18567 38913
rect 18524 38876 18552 38907
rect 20806 38904 20812 38916
rect 20864 38904 20870 38956
rect 21082 38944 21088 38956
rect 21043 38916 21088 38944
rect 21082 38904 21088 38916
rect 21140 38944 21146 38956
rect 21818 38944 21824 38956
rect 21140 38916 21824 38944
rect 21140 38904 21146 38916
rect 21818 38904 21824 38916
rect 21876 38904 21882 38956
rect 22002 38904 22008 38956
rect 22060 38944 22066 38956
rect 22060 38916 22153 38944
rect 22060 38904 22066 38916
rect 22554 38904 22560 38956
rect 22612 38944 22618 38956
rect 23109 38947 23167 38953
rect 23109 38944 23121 38947
rect 22612 38916 23121 38944
rect 22612 38904 22618 38916
rect 23109 38913 23121 38916
rect 23155 38913 23167 38947
rect 23290 38944 23296 38956
rect 23251 38916 23296 38944
rect 23109 38907 23167 38913
rect 23290 38904 23296 38916
rect 23348 38904 23354 38956
rect 23753 38947 23811 38953
rect 23753 38913 23765 38947
rect 23799 38944 23811 38947
rect 23934 38944 23940 38956
rect 23799 38916 23940 38944
rect 23799 38913 23811 38916
rect 23753 38907 23811 38913
rect 23934 38904 23940 38916
rect 23992 38904 23998 38956
rect 24029 38947 24087 38953
rect 24029 38913 24041 38947
rect 24075 38944 24087 38947
rect 24854 38944 24860 38956
rect 24075 38916 24860 38944
rect 24075 38913 24087 38916
rect 24029 38907 24087 38913
rect 24854 38904 24860 38916
rect 24912 38904 24918 38956
rect 25222 38904 25228 38956
rect 25280 38944 25286 38956
rect 26620 38944 26648 38984
rect 27154 38944 27160 38956
rect 25280 38916 26648 38944
rect 27115 38916 27160 38944
rect 25280 38904 25286 38916
rect 27154 38904 27160 38916
rect 27212 38904 27218 38956
rect 27246 38904 27252 38956
rect 27304 38944 27310 38956
rect 27341 38947 27399 38953
rect 27341 38944 27353 38947
rect 27304 38916 27353 38944
rect 27304 38904 27310 38916
rect 27341 38913 27353 38916
rect 27387 38913 27399 38947
rect 27341 38907 27399 38913
rect 27430 38904 27436 38956
rect 27488 38944 27494 38956
rect 29457 38947 29515 38953
rect 27488 38916 27533 38944
rect 27488 38904 27494 38916
rect 29457 38913 29469 38947
rect 29503 38913 29515 38947
rect 29457 38907 29515 38913
rect 29733 38947 29791 38953
rect 29733 38913 29745 38947
rect 29779 38944 29791 38947
rect 30558 38944 30564 38956
rect 29779 38916 30564 38944
rect 29779 38913 29791 38916
rect 29733 38907 29791 38913
rect 17512 38848 18552 38876
rect 19337 38879 19395 38885
rect 19337 38845 19349 38879
rect 19383 38876 19395 38879
rect 19518 38876 19524 38888
rect 19383 38848 19524 38876
rect 19383 38845 19395 38848
rect 19337 38839 19395 38845
rect 19518 38836 19524 38848
rect 19576 38876 19582 38888
rect 20990 38876 20996 38888
rect 19576 38848 20852 38876
rect 20951 38848 20996 38876
rect 19576 38836 19582 38848
rect 18601 38811 18659 38817
rect 18601 38777 18613 38811
rect 18647 38808 18659 38811
rect 19426 38808 19432 38820
rect 18647 38780 19432 38808
rect 18647 38777 18659 38780
rect 18601 38771 18659 38777
rect 19426 38768 19432 38780
rect 19484 38808 19490 38820
rect 20824 38808 20852 38848
rect 20990 38836 20996 38848
rect 21048 38836 21054 38888
rect 21266 38836 21272 38888
rect 21324 38876 21330 38888
rect 21913 38879 21971 38885
rect 21913 38876 21925 38879
rect 21324 38848 21925 38876
rect 21324 38836 21330 38848
rect 21913 38845 21925 38848
rect 21959 38845 21971 38879
rect 21913 38839 21971 38845
rect 22186 38836 22192 38888
rect 22244 38876 22250 38888
rect 29472 38876 29500 38907
rect 30558 38904 30564 38916
rect 30616 38904 30622 38956
rect 30668 38953 30696 38984
rect 31386 38972 31392 38984
rect 31444 38972 31450 39024
rect 31570 39012 31576 39024
rect 31531 38984 31576 39012
rect 31570 38972 31576 38984
rect 31628 38972 31634 39024
rect 30653 38947 30711 38953
rect 30653 38913 30665 38947
rect 30699 38913 30711 38947
rect 30653 38907 30711 38913
rect 30745 38947 30803 38953
rect 30745 38913 30757 38947
rect 30791 38913 30803 38947
rect 30926 38944 30932 38956
rect 30887 38916 30932 38944
rect 30745 38907 30803 38913
rect 30466 38876 30472 38888
rect 22244 38848 28994 38876
rect 29472 38848 30472 38876
rect 22244 38836 22250 38848
rect 25222 38808 25228 38820
rect 19484 38780 20024 38808
rect 20824 38780 25228 38808
rect 19484 38768 19490 38780
rect 1949 38743 2007 38749
rect 1949 38709 1961 38743
rect 1995 38740 2007 38743
rect 15378 38740 15384 38752
rect 1995 38712 15384 38740
rect 1995 38709 2007 38712
rect 1949 38703 2007 38709
rect 15378 38700 15384 38712
rect 15436 38700 15442 38752
rect 16669 38743 16727 38749
rect 16669 38709 16681 38743
rect 16715 38740 16727 38743
rect 17494 38740 17500 38752
rect 16715 38712 17500 38740
rect 16715 38709 16727 38712
rect 16669 38703 16727 38709
rect 17494 38700 17500 38712
rect 17552 38700 17558 38752
rect 19996 38749 20024 38780
rect 25222 38768 25228 38780
rect 25280 38768 25286 38820
rect 27246 38768 27252 38820
rect 27304 38808 27310 38820
rect 27893 38811 27951 38817
rect 27893 38808 27905 38811
rect 27304 38780 27905 38808
rect 27304 38768 27310 38780
rect 27893 38777 27905 38780
rect 27939 38777 27951 38811
rect 27893 38771 27951 38777
rect 19981 38743 20039 38749
rect 19981 38709 19993 38743
rect 20027 38709 20039 38743
rect 19981 38703 20039 38709
rect 20990 38700 20996 38752
rect 21048 38740 21054 38752
rect 21450 38740 21456 38752
rect 21048 38712 21456 38740
rect 21048 38700 21054 38712
rect 21450 38700 21456 38712
rect 21508 38740 21514 38752
rect 22186 38740 22192 38752
rect 21508 38712 22192 38740
rect 21508 38700 21514 38712
rect 22186 38700 22192 38712
rect 22244 38700 22250 38752
rect 24213 38743 24271 38749
rect 24213 38709 24225 38743
rect 24259 38740 24271 38743
rect 24394 38740 24400 38752
rect 24259 38712 24400 38740
rect 24259 38709 24271 38712
rect 24213 38703 24271 38709
rect 24394 38700 24400 38712
rect 24452 38700 24458 38752
rect 24670 38700 24676 38752
rect 24728 38740 24734 38752
rect 25777 38743 25835 38749
rect 25777 38740 25789 38743
rect 24728 38712 25789 38740
rect 24728 38700 24734 38712
rect 25777 38709 25789 38712
rect 25823 38709 25835 38743
rect 26326 38740 26332 38752
rect 26287 38712 26332 38740
rect 25777 38703 25835 38709
rect 26326 38700 26332 38712
rect 26384 38700 26390 38752
rect 28966 38740 28994 38848
rect 30466 38836 30472 38848
rect 30524 38836 30530 38888
rect 30760 38876 30788 38907
rect 30926 38904 30932 38916
rect 30984 38904 30990 38956
rect 31018 38904 31024 38956
rect 31076 38944 31082 38956
rect 32392 38947 32450 38953
rect 31076 38916 31121 38944
rect 31076 38904 31082 38916
rect 32392 38913 32404 38947
rect 32438 38944 32450 38947
rect 32950 38944 32956 38956
rect 32438 38916 32956 38944
rect 32438 38913 32450 38916
rect 32392 38907 32450 38913
rect 32950 38904 32956 38916
rect 33008 38904 33014 38956
rect 31202 38876 31208 38888
rect 30760 38848 31208 38876
rect 31202 38836 31208 38848
rect 31260 38836 31266 38888
rect 32125 38879 32183 38885
rect 32125 38845 32137 38879
rect 32171 38845 32183 38879
rect 32125 38839 32183 38845
rect 30282 38768 30288 38820
rect 30340 38808 30346 38820
rect 32140 38808 32168 38839
rect 30340 38780 32168 38808
rect 33336 38808 33364 39052
rect 35069 39049 35081 39083
rect 35115 39080 35127 39083
rect 36354 39080 36360 39092
rect 35115 39052 36360 39080
rect 35115 39049 35127 39052
rect 35069 39043 35127 39049
rect 36354 39040 36360 39052
rect 36412 39040 36418 39092
rect 37274 39040 37280 39092
rect 37332 39080 37338 39092
rect 37435 39083 37493 39089
rect 37435 39080 37447 39083
rect 37332 39052 37447 39080
rect 37332 39040 37338 39052
rect 37435 39049 37447 39052
rect 37481 39049 37493 39083
rect 37435 39043 37493 39049
rect 38378 39040 38384 39092
rect 38436 39080 38442 39092
rect 38473 39083 38531 39089
rect 38473 39080 38485 39083
rect 38436 39052 38485 39080
rect 38436 39040 38442 39052
rect 38473 39049 38485 39052
rect 38519 39049 38531 39083
rect 38473 39043 38531 39049
rect 38562 39040 38568 39092
rect 38620 39080 38626 39092
rect 39485 39083 39543 39089
rect 39485 39080 39497 39083
rect 38620 39052 39497 39080
rect 38620 39040 38626 39052
rect 39485 39049 39497 39052
rect 39531 39049 39543 39083
rect 40034 39080 40040 39092
rect 39995 39052 40040 39080
rect 39485 39043 39543 39049
rect 40034 39040 40040 39052
rect 40092 39040 40098 39092
rect 34974 38972 34980 39024
rect 35032 39012 35038 39024
rect 35161 39015 35219 39021
rect 35161 39012 35173 39015
rect 35032 38984 35173 39012
rect 35032 38972 35038 38984
rect 35161 38981 35173 38984
rect 35207 39012 35219 39015
rect 35526 39012 35532 39024
rect 35207 38984 35532 39012
rect 35207 38981 35219 38984
rect 35161 38975 35219 38981
rect 35526 38972 35532 38984
rect 35584 38972 35590 39024
rect 36449 39015 36507 39021
rect 36449 38981 36461 39015
rect 36495 39012 36507 39015
rect 37645 39015 37703 39021
rect 37645 39012 37657 39015
rect 36495 38984 37657 39012
rect 36495 38981 36507 38984
rect 36449 38975 36507 38981
rect 37645 38981 37657 38984
rect 37691 38981 37703 39015
rect 37645 38975 37703 38981
rect 34146 38904 34152 38956
rect 34204 38944 34210 38956
rect 34241 38947 34299 38953
rect 34241 38944 34253 38947
rect 34204 38916 34253 38944
rect 34204 38904 34210 38916
rect 34241 38913 34253 38916
rect 34287 38913 34299 38947
rect 34422 38944 34428 38956
rect 34383 38916 34428 38944
rect 34241 38907 34299 38913
rect 34422 38904 34428 38916
rect 34480 38904 34486 38956
rect 35250 38944 35256 38956
rect 35211 38916 35256 38944
rect 35250 38904 35256 38916
rect 35308 38904 35314 38956
rect 35437 38947 35495 38953
rect 35437 38913 35449 38947
rect 35483 38944 35495 38947
rect 35618 38944 35624 38956
rect 35483 38916 35624 38944
rect 35483 38913 35495 38916
rect 35437 38907 35495 38913
rect 35618 38904 35624 38916
rect 35676 38904 35682 38956
rect 36633 38947 36691 38953
rect 36633 38913 36645 38947
rect 36679 38913 36691 38947
rect 36633 38907 36691 38913
rect 36725 38947 36783 38953
rect 36725 38913 36737 38947
rect 36771 38944 36783 38947
rect 37274 38944 37280 38956
rect 36771 38916 37280 38944
rect 36771 38913 36783 38916
rect 36725 38907 36783 38913
rect 33410 38836 33416 38888
rect 33468 38876 33474 38888
rect 34885 38879 34943 38885
rect 34885 38876 34897 38879
rect 33468 38848 34897 38876
rect 33468 38836 33474 38848
rect 34885 38845 34897 38848
rect 34931 38845 34943 38879
rect 36648 38876 36676 38907
rect 37274 38904 37280 38916
rect 37332 38904 37338 38956
rect 37660 38944 37688 38975
rect 38378 38944 38384 38956
rect 37660 38916 38384 38944
rect 38378 38904 38384 38916
rect 38436 38904 38442 38956
rect 38654 38904 38660 38956
rect 38712 38944 38718 38956
rect 38841 38947 38899 38953
rect 38841 38944 38853 38947
rect 38712 38916 38853 38944
rect 38712 38904 38718 38916
rect 38841 38913 38853 38916
rect 38887 38913 38899 38947
rect 38841 38907 38899 38913
rect 37458 38876 37464 38888
rect 36648 38848 37464 38876
rect 34885 38839 34943 38845
rect 37458 38836 37464 38848
rect 37516 38836 37522 38888
rect 38930 38876 38936 38888
rect 38891 38848 38936 38876
rect 38930 38836 38936 38848
rect 38988 38836 38994 38888
rect 38838 38808 38844 38820
rect 33336 38780 38844 38808
rect 30340 38768 30346 38780
rect 38838 38768 38844 38780
rect 38896 38768 38902 38820
rect 30469 38743 30527 38749
rect 30469 38740 30481 38743
rect 28966 38712 30481 38740
rect 30469 38709 30481 38712
rect 30515 38709 30527 38743
rect 30469 38703 30527 38709
rect 31202 38700 31208 38752
rect 31260 38740 31266 38752
rect 32490 38740 32496 38752
rect 31260 38712 32496 38740
rect 31260 38700 31266 38712
rect 32490 38700 32496 38712
rect 32548 38740 32554 38752
rect 33410 38740 33416 38752
rect 32548 38712 33416 38740
rect 32548 38700 32554 38712
rect 33410 38700 33416 38712
rect 33468 38700 33474 38752
rect 33505 38743 33563 38749
rect 33505 38709 33517 38743
rect 33551 38740 33563 38743
rect 33778 38740 33784 38752
rect 33551 38712 33784 38740
rect 33551 38709 33563 38712
rect 33505 38703 33563 38709
rect 33778 38700 33784 38712
rect 33836 38700 33842 38752
rect 34054 38740 34060 38752
rect 34015 38712 34060 38740
rect 34054 38700 34060 38712
rect 34112 38700 34118 38752
rect 34425 38743 34483 38749
rect 34425 38709 34437 38743
rect 34471 38740 34483 38743
rect 34790 38740 34796 38752
rect 34471 38712 34796 38740
rect 34471 38709 34483 38712
rect 34425 38703 34483 38709
rect 34790 38700 34796 38712
rect 34848 38700 34854 38752
rect 35986 38740 35992 38752
rect 35947 38712 35992 38740
rect 35986 38700 35992 38712
rect 36044 38700 36050 38752
rect 36446 38740 36452 38752
rect 36407 38712 36452 38740
rect 36446 38700 36452 38712
rect 36504 38700 36510 38752
rect 37274 38740 37280 38752
rect 37235 38712 37280 38740
rect 37274 38700 37280 38712
rect 37332 38700 37338 38752
rect 37458 38740 37464 38752
rect 37419 38712 37464 38740
rect 37458 38700 37464 38712
rect 37516 38700 37522 38752
rect 40034 38700 40040 38752
rect 40092 38740 40098 38752
rect 40402 38740 40408 38752
rect 40092 38712 40408 38740
rect 40092 38700 40098 38712
rect 40402 38700 40408 38712
rect 40460 38740 40466 38752
rect 40589 38743 40647 38749
rect 40589 38740 40601 38743
rect 40460 38712 40601 38740
rect 40460 38700 40466 38712
rect 40589 38709 40601 38712
rect 40635 38709 40647 38743
rect 40589 38703 40647 38709
rect 1104 38650 54372 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 54372 38650
rect 1104 38576 54372 38598
rect 1578 38536 1584 38548
rect 1539 38508 1584 38536
rect 1578 38496 1584 38508
rect 1636 38496 1642 38548
rect 16666 38536 16672 38548
rect 16627 38508 16672 38536
rect 16666 38496 16672 38508
rect 16724 38496 16730 38548
rect 26510 38536 26516 38548
rect 26423 38508 26516 38536
rect 26510 38496 26516 38508
rect 26568 38536 26574 38548
rect 27706 38536 27712 38548
rect 26568 38508 27712 38536
rect 26568 38496 26574 38508
rect 27706 38496 27712 38508
rect 27764 38496 27770 38548
rect 28997 38539 29055 38545
rect 28997 38505 29009 38539
rect 29043 38536 29055 38539
rect 30006 38536 30012 38548
rect 29043 38508 30012 38536
rect 29043 38505 29055 38508
rect 28997 38499 29055 38505
rect 30006 38496 30012 38508
rect 30064 38496 30070 38548
rect 30653 38539 30711 38545
rect 30653 38505 30665 38539
rect 30699 38536 30711 38539
rect 30926 38536 30932 38548
rect 30699 38508 30932 38536
rect 30699 38505 30711 38508
rect 30653 38499 30711 38505
rect 30926 38496 30932 38508
rect 30984 38496 30990 38548
rect 32950 38536 32956 38548
rect 32911 38508 32956 38536
rect 32950 38496 32956 38508
rect 33008 38496 33014 38548
rect 34790 38536 34796 38548
rect 34751 38508 34796 38536
rect 34790 38496 34796 38508
rect 34848 38496 34854 38548
rect 34977 38539 35035 38545
rect 34977 38505 34989 38539
rect 35023 38536 35035 38539
rect 35342 38536 35348 38548
rect 35023 38508 35348 38536
rect 35023 38505 35035 38508
rect 34977 38499 35035 38505
rect 35342 38496 35348 38508
rect 35400 38496 35406 38548
rect 36219 38539 36277 38545
rect 36219 38505 36231 38539
rect 36265 38536 36277 38539
rect 36446 38536 36452 38548
rect 36265 38508 36452 38536
rect 36265 38505 36277 38508
rect 36219 38499 36277 38505
rect 36446 38496 36452 38508
rect 36504 38536 36510 38548
rect 37001 38539 37059 38545
rect 37001 38536 37013 38539
rect 36504 38508 37013 38536
rect 36504 38496 36510 38508
rect 37001 38505 37013 38508
rect 37047 38505 37059 38539
rect 37001 38499 37059 38505
rect 23845 38471 23903 38477
rect 23845 38437 23857 38471
rect 23891 38468 23903 38471
rect 25314 38468 25320 38480
rect 23891 38440 25320 38468
rect 23891 38437 23903 38440
rect 23845 38431 23903 38437
rect 25314 38428 25320 38440
rect 25372 38428 25378 38480
rect 21266 38400 21272 38412
rect 16868 38372 19288 38400
rect 15289 38335 15347 38341
rect 15289 38301 15301 38335
rect 15335 38332 15347 38335
rect 15470 38332 15476 38344
rect 15335 38304 15476 38332
rect 15335 38301 15347 38304
rect 15289 38295 15347 38301
rect 15470 38292 15476 38304
rect 15528 38332 15534 38344
rect 15528 38304 16528 38332
rect 15528 38292 15534 38304
rect 16500 38276 16528 38304
rect 16298 38264 16304 38276
rect 16259 38236 16304 38264
rect 16298 38224 16304 38236
rect 16356 38224 16362 38276
rect 16482 38264 16488 38276
rect 16443 38236 16488 38264
rect 16482 38224 16488 38236
rect 16540 38224 16546 38276
rect 15841 38199 15899 38205
rect 15841 38165 15853 38199
rect 15887 38196 15899 38199
rect 16390 38196 16396 38208
rect 15887 38168 16396 38196
rect 15887 38165 15899 38168
rect 15841 38159 15899 38165
rect 16390 38156 16396 38168
rect 16448 38196 16454 38208
rect 16868 38196 16896 38372
rect 19260 38344 19288 38372
rect 20456 38372 21272 38400
rect 17218 38332 17224 38344
rect 17179 38304 17224 38332
rect 17218 38292 17224 38304
rect 17276 38292 17282 38344
rect 17494 38332 17500 38344
rect 17455 38304 17500 38332
rect 17494 38292 17500 38304
rect 17552 38292 17558 38344
rect 18138 38332 18144 38344
rect 18051 38304 18144 38332
rect 18138 38292 18144 38304
rect 18196 38292 18202 38344
rect 18322 38332 18328 38344
rect 18283 38304 18328 38332
rect 18322 38292 18328 38304
rect 18380 38292 18386 38344
rect 19242 38332 19248 38344
rect 19203 38304 19248 38332
rect 19242 38292 19248 38304
rect 19300 38292 19306 38344
rect 19429 38335 19487 38341
rect 19429 38301 19441 38335
rect 19475 38332 19487 38335
rect 19518 38332 19524 38344
rect 19475 38304 19524 38332
rect 19475 38301 19487 38304
rect 19429 38295 19487 38301
rect 19518 38292 19524 38304
rect 19576 38292 19582 38344
rect 20162 38332 20168 38344
rect 20123 38304 20168 38332
rect 20162 38292 20168 38304
rect 20220 38292 20226 38344
rect 20456 38341 20484 38372
rect 21266 38360 21272 38372
rect 21324 38360 21330 38412
rect 22002 38360 22008 38412
rect 22060 38400 22066 38412
rect 23017 38403 23075 38409
rect 23017 38400 23029 38403
rect 22060 38372 23029 38400
rect 22060 38360 22066 38372
rect 23017 38369 23029 38372
rect 23063 38369 23075 38403
rect 23017 38363 23075 38369
rect 24412 38372 25452 38400
rect 24412 38344 24440 38372
rect 20441 38335 20499 38341
rect 20441 38301 20453 38335
rect 20487 38301 20499 38335
rect 20898 38332 20904 38344
rect 20811 38304 20904 38332
rect 20441 38295 20499 38301
rect 16942 38224 16948 38276
rect 17000 38264 17006 38276
rect 17313 38267 17371 38273
rect 17313 38264 17325 38267
rect 17000 38236 17325 38264
rect 17000 38224 17006 38236
rect 17313 38233 17325 38236
rect 17359 38233 17371 38267
rect 18156 38264 18184 38292
rect 19337 38267 19395 38273
rect 19337 38264 19349 38267
rect 18156 38236 19349 38264
rect 17313 38227 17371 38233
rect 19337 38233 19349 38236
rect 19383 38233 19395 38267
rect 19337 38227 19395 38233
rect 19981 38267 20039 38273
rect 19981 38233 19993 38267
rect 20027 38264 20039 38267
rect 20824 38264 20852 38304
rect 20898 38292 20904 38304
rect 20956 38292 20962 38344
rect 21174 38332 21180 38344
rect 21135 38304 21180 38332
rect 21174 38292 21180 38304
rect 21232 38292 21238 38344
rect 21634 38292 21640 38344
rect 21692 38332 21698 38344
rect 21821 38335 21879 38341
rect 21821 38332 21833 38335
rect 21692 38304 21833 38332
rect 21692 38292 21698 38304
rect 21821 38301 21833 38304
rect 21867 38301 21879 38335
rect 22186 38332 22192 38344
rect 22147 38304 22192 38332
rect 21821 38295 21879 38301
rect 22186 38292 22192 38304
rect 22244 38292 22250 38344
rect 22830 38332 22836 38344
rect 22791 38304 22836 38332
rect 22830 38292 22836 38304
rect 22888 38292 22894 38344
rect 24394 38332 24400 38344
rect 24355 38304 24400 38332
rect 24394 38292 24400 38304
rect 24452 38292 24458 38344
rect 25424 38341 25452 38372
rect 25225 38335 25283 38341
rect 25225 38332 25237 38335
rect 24596 38304 25237 38332
rect 20027 38236 20852 38264
rect 20027 38233 20039 38236
rect 19981 38227 20039 38233
rect 21082 38224 21088 38276
rect 21140 38264 21146 38276
rect 21913 38267 21971 38273
rect 21913 38264 21925 38267
rect 21140 38236 21925 38264
rect 21140 38224 21146 38236
rect 21913 38233 21925 38236
rect 21959 38264 21971 38267
rect 22649 38267 22707 38273
rect 22649 38264 22661 38267
rect 21959 38236 22661 38264
rect 21959 38233 21971 38236
rect 21913 38227 21971 38233
rect 22649 38233 22661 38236
rect 22695 38233 22707 38267
rect 22649 38227 22707 38233
rect 24026 38224 24032 38276
rect 24084 38264 24090 38276
rect 24596 38273 24624 38304
rect 25225 38301 25237 38304
rect 25271 38301 25283 38335
rect 25225 38295 25283 38301
rect 25409 38335 25467 38341
rect 25409 38301 25421 38335
rect 25455 38301 25467 38335
rect 26050 38332 26056 38344
rect 26011 38304 26056 38332
rect 25409 38295 25467 38301
rect 26050 38292 26056 38304
rect 26108 38292 26114 38344
rect 26237 38335 26295 38341
rect 26237 38301 26249 38335
rect 26283 38332 26295 38335
rect 26528 38332 26556 38496
rect 26694 38468 26700 38480
rect 26655 38440 26700 38468
rect 26694 38428 26700 38440
rect 26752 38428 26758 38480
rect 27338 38428 27344 38480
rect 27396 38468 27402 38480
rect 27433 38471 27491 38477
rect 27433 38468 27445 38471
rect 27396 38440 27445 38468
rect 27396 38428 27402 38440
rect 27433 38437 27445 38440
rect 27479 38437 27491 38471
rect 30834 38468 30840 38480
rect 27433 38431 27491 38437
rect 30300 38440 30840 38468
rect 27985 38403 28043 38409
rect 27985 38400 27997 38403
rect 26712 38372 27997 38400
rect 26712 38341 26740 38372
rect 27985 38369 27997 38372
rect 28031 38369 28043 38403
rect 29914 38400 29920 38412
rect 27985 38363 28043 38369
rect 28736 38372 29920 38400
rect 26283 38304 26556 38332
rect 26697 38335 26755 38341
rect 26283 38301 26295 38304
rect 26237 38295 26295 38301
rect 26697 38301 26709 38335
rect 26743 38301 26755 38335
rect 26697 38295 26755 38301
rect 24581 38267 24639 38273
rect 24581 38264 24593 38267
rect 24084 38236 24593 38264
rect 24084 38224 24090 38236
rect 24581 38233 24593 38236
rect 24627 38233 24639 38267
rect 24581 38227 24639 38233
rect 24670 38224 24676 38276
rect 24728 38264 24734 38276
rect 26602 38264 26608 38276
rect 24728 38236 26608 38264
rect 24728 38224 24734 38236
rect 26602 38224 26608 38236
rect 26660 38264 26666 38276
rect 26712 38264 26740 38295
rect 26878 38292 26884 38344
rect 26936 38332 26942 38344
rect 26973 38335 27031 38341
rect 26973 38332 26985 38335
rect 26936 38304 26985 38332
rect 26936 38292 26942 38304
rect 26973 38301 26985 38304
rect 27019 38332 27031 38335
rect 27430 38332 27436 38344
rect 27019 38304 27436 38332
rect 27019 38301 27031 38304
rect 26973 38295 27031 38301
rect 27430 38292 27436 38304
rect 27488 38292 27494 38344
rect 28736 38341 28764 38372
rect 29914 38360 29920 38372
rect 29972 38360 29978 38412
rect 28721 38335 28779 38341
rect 28721 38301 28733 38335
rect 28767 38301 28779 38335
rect 28721 38295 28779 38301
rect 28813 38335 28871 38341
rect 28813 38301 28825 38335
rect 28859 38332 28871 38335
rect 29825 38335 29883 38341
rect 29825 38332 29837 38335
rect 28859 38304 29837 38332
rect 28859 38301 28871 38304
rect 28813 38295 28871 38301
rect 29825 38301 29837 38304
rect 29871 38332 29883 38335
rect 30300 38332 30328 38440
rect 30834 38428 30840 38440
rect 30892 38468 30898 38480
rect 30892 38440 31064 38468
rect 30892 38428 30898 38440
rect 31036 38409 31064 38440
rect 35802 38428 35808 38480
rect 35860 38468 35866 38480
rect 35860 38440 37504 38468
rect 35860 38428 35866 38440
rect 31021 38403 31079 38409
rect 31021 38369 31033 38403
rect 31067 38369 31079 38403
rect 31021 38363 31079 38369
rect 36357 38403 36415 38409
rect 36357 38369 36369 38403
rect 36403 38400 36415 38403
rect 36403 38372 37320 38400
rect 36403 38369 36415 38372
rect 36357 38363 36415 38369
rect 37292 38344 37320 38372
rect 31297 38335 31355 38341
rect 30827 38332 30972 38334
rect 29871 38304 30328 38332
rect 30392 38306 31064 38332
rect 30392 38304 30855 38306
rect 30944 38304 31064 38306
rect 29871 38301 29883 38304
rect 29825 38295 29883 38301
rect 27062 38264 27068 38276
rect 26660 38236 26740 38264
rect 26804 38236 27068 38264
rect 26660 38224 26666 38236
rect 17678 38196 17684 38208
rect 16448 38168 16896 38196
rect 17639 38168 17684 38196
rect 16448 38156 16454 38168
rect 17678 38156 17684 38168
rect 17736 38156 17742 38208
rect 17770 38156 17776 38208
rect 17828 38196 17834 38208
rect 18141 38199 18199 38205
rect 18141 38196 18153 38199
rect 17828 38168 18153 38196
rect 17828 38156 17834 38168
rect 18141 38165 18153 38168
rect 18187 38165 18199 38199
rect 18141 38159 18199 38165
rect 20349 38199 20407 38205
rect 20349 38165 20361 38199
rect 20395 38196 20407 38199
rect 20714 38196 20720 38208
rect 20395 38168 20720 38196
rect 20395 38165 20407 38168
rect 20349 38159 20407 38165
rect 20714 38156 20720 38168
rect 20772 38156 20778 38208
rect 20990 38196 20996 38208
rect 20951 38168 20996 38196
rect 20990 38156 20996 38168
rect 21048 38156 21054 38208
rect 21358 38196 21364 38208
rect 21319 38168 21364 38196
rect 21358 38156 21364 38168
rect 21416 38156 21422 38208
rect 21818 38156 21824 38208
rect 21876 38196 21882 38208
rect 22005 38199 22063 38205
rect 22005 38196 22017 38199
rect 21876 38168 22017 38196
rect 21876 38156 21882 38168
rect 22005 38165 22017 38168
rect 22051 38165 22063 38199
rect 22005 38159 22063 38165
rect 22094 38156 22100 38208
rect 22152 38196 22158 38208
rect 24762 38196 24768 38208
rect 22152 38168 22197 38196
rect 24723 38168 24768 38196
rect 22152 38156 22158 38168
rect 24762 38156 24768 38168
rect 24820 38156 24826 38208
rect 25222 38196 25228 38208
rect 25183 38168 25228 38196
rect 25222 38156 25228 38168
rect 25280 38156 25286 38208
rect 26145 38199 26203 38205
rect 26145 38165 26157 38199
rect 26191 38196 26203 38199
rect 26804 38196 26832 38236
rect 27062 38224 27068 38236
rect 27120 38224 27126 38276
rect 28997 38267 29055 38273
rect 28997 38233 29009 38267
rect 29043 38264 29055 38267
rect 30392 38264 30420 38304
rect 29043 38236 30420 38264
rect 30812 38267 30870 38273
rect 29043 38233 29055 38236
rect 28997 38227 29055 38233
rect 30812 38233 30824 38267
rect 30858 38233 30870 38267
rect 30812 38227 30870 38233
rect 26191 38168 26832 38196
rect 26881 38199 26939 38205
rect 26191 38165 26203 38168
rect 26145 38159 26203 38165
rect 26881 38165 26893 38199
rect 26927 38196 26939 38199
rect 27154 38196 27160 38208
rect 26927 38168 27160 38196
rect 26927 38165 26939 38168
rect 26881 38159 26939 38165
rect 27154 38156 27160 38168
rect 27212 38156 27218 38208
rect 30098 38156 30104 38208
rect 30156 38196 30162 38208
rect 30193 38199 30251 38205
rect 30193 38196 30205 38199
rect 30156 38168 30205 38196
rect 30156 38156 30162 38168
rect 30193 38165 30205 38168
rect 30239 38165 30251 38199
rect 30193 38159 30251 38165
rect 30558 38156 30564 38208
rect 30616 38196 30622 38208
rect 30827 38196 30855 38227
rect 30926 38196 30932 38208
rect 30616 38168 30855 38196
rect 30887 38168 30932 38196
rect 30616 38156 30622 38168
rect 30926 38156 30932 38168
rect 30984 38156 30990 38208
rect 31036 38196 31064 38304
rect 31297 38301 31309 38335
rect 31343 38332 31355 38335
rect 31938 38332 31944 38344
rect 31343 38304 31754 38332
rect 31899 38304 31944 38332
rect 31343 38301 31355 38304
rect 31297 38295 31355 38301
rect 31726 38264 31754 38304
rect 31938 38292 31944 38304
rect 31996 38292 32002 38344
rect 32030 38292 32036 38344
rect 32088 38332 32094 38344
rect 33229 38335 33287 38341
rect 32088 38304 32133 38332
rect 32088 38292 32094 38304
rect 33229 38301 33241 38335
rect 33275 38332 33287 38335
rect 33410 38332 33416 38344
rect 33275 38304 33416 38332
rect 33275 38301 33287 38304
rect 33229 38295 33287 38301
rect 33410 38292 33416 38304
rect 33468 38292 33474 38344
rect 33594 38332 33600 38344
rect 33555 38304 33600 38332
rect 33594 38292 33600 38304
rect 33652 38292 33658 38344
rect 33686 38292 33692 38344
rect 33744 38332 33750 38344
rect 33744 38304 35296 38332
rect 33744 38292 33750 38304
rect 32582 38264 32588 38276
rect 31726 38236 32588 38264
rect 32582 38224 32588 38236
rect 32640 38224 32646 38276
rect 33321 38267 33379 38273
rect 33321 38233 33333 38267
rect 33367 38264 33379 38267
rect 34054 38264 34060 38276
rect 33367 38236 34060 38264
rect 33367 38233 33379 38236
rect 33321 38227 33379 38233
rect 34054 38224 34060 38236
rect 34112 38224 34118 38276
rect 34698 38224 34704 38276
rect 34756 38264 34762 38276
rect 35158 38264 35164 38276
rect 34756 38236 35164 38264
rect 34756 38224 34762 38236
rect 35158 38224 35164 38236
rect 35216 38224 35222 38276
rect 35268 38264 35296 38304
rect 35342 38292 35348 38344
rect 35400 38332 35406 38344
rect 36081 38335 36139 38341
rect 36081 38332 36093 38335
rect 35400 38304 36093 38332
rect 35400 38292 35406 38304
rect 36081 38301 36093 38304
rect 36127 38301 36139 38335
rect 36081 38295 36139 38301
rect 36541 38335 36599 38341
rect 36541 38301 36553 38335
rect 36587 38332 36599 38335
rect 37182 38332 37188 38344
rect 36587 38304 37188 38332
rect 36587 38301 36599 38304
rect 36541 38295 36599 38301
rect 37182 38292 37188 38304
rect 37240 38292 37246 38344
rect 37274 38292 37280 38344
rect 37332 38332 37338 38344
rect 37476 38341 37504 38440
rect 37461 38335 37519 38341
rect 37332 38304 37377 38332
rect 37332 38292 37338 38304
rect 37461 38301 37473 38335
rect 37507 38301 37519 38335
rect 38470 38332 38476 38344
rect 38431 38304 38476 38332
rect 37461 38295 37519 38301
rect 38470 38292 38476 38304
rect 38528 38292 38534 38344
rect 35894 38264 35900 38276
rect 35268 38236 35900 38264
rect 35894 38224 35900 38236
rect 35952 38264 35958 38276
rect 37921 38267 37979 38273
rect 37921 38264 37933 38267
rect 35952 38236 37933 38264
rect 35952 38224 35958 38236
rect 37921 38233 37933 38236
rect 37967 38233 37979 38267
rect 37921 38227 37979 38233
rect 38378 38224 38384 38276
rect 38436 38264 38442 38276
rect 39025 38267 39083 38273
rect 39025 38264 39037 38267
rect 38436 38236 39037 38264
rect 38436 38224 38442 38236
rect 39025 38233 39037 38236
rect 39071 38264 39083 38267
rect 40034 38264 40040 38276
rect 39071 38236 40040 38264
rect 39071 38233 39083 38236
rect 39025 38227 39083 38233
rect 40034 38224 40040 38236
rect 40092 38224 40098 38276
rect 31757 38199 31815 38205
rect 31757 38196 31769 38199
rect 31036 38168 31769 38196
rect 31757 38165 31769 38168
rect 31803 38165 31815 38199
rect 31757 38159 31815 38165
rect 33410 38156 33416 38208
rect 33468 38196 33474 38208
rect 34961 38199 35019 38205
rect 33468 38168 33513 38196
rect 33468 38156 33474 38168
rect 34961 38165 34973 38199
rect 35007 38196 35019 38199
rect 35526 38196 35532 38208
rect 35007 38168 35532 38196
rect 35007 38165 35019 38168
rect 34961 38159 35019 38165
rect 35526 38156 35532 38168
rect 35584 38156 35590 38208
rect 36541 38199 36599 38205
rect 36541 38165 36553 38199
rect 36587 38196 36599 38199
rect 36630 38196 36636 38208
rect 36587 38168 36636 38196
rect 36587 38165 36599 38168
rect 36541 38159 36599 38165
rect 36630 38156 36636 38168
rect 36688 38156 36694 38208
rect 37182 38196 37188 38208
rect 37143 38168 37188 38196
rect 37182 38156 37188 38168
rect 37240 38156 37246 38208
rect 38654 38156 38660 38208
rect 38712 38196 38718 38208
rect 39850 38196 39856 38208
rect 38712 38168 39856 38196
rect 38712 38156 38718 38168
rect 39850 38156 39856 38168
rect 39908 38156 39914 38208
rect 1104 38106 54372 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 54372 38106
rect 1104 38032 54372 38054
rect 15565 37995 15623 38001
rect 15565 37961 15577 37995
rect 15611 37992 15623 37995
rect 16298 37992 16304 38004
rect 15611 37964 16304 37992
rect 15611 37961 15623 37964
rect 15565 37955 15623 37961
rect 16298 37952 16304 37964
rect 16356 37952 16362 38004
rect 17497 37995 17555 38001
rect 17497 37961 17509 37995
rect 17543 37992 17555 37995
rect 17678 37992 17684 38004
rect 17543 37964 17684 37992
rect 17543 37961 17555 37964
rect 17497 37955 17555 37961
rect 17678 37952 17684 37964
rect 17736 37952 17742 38004
rect 19426 37992 19432 38004
rect 18340 37964 19432 37992
rect 16945 37927 17003 37933
rect 16945 37893 16957 37927
rect 16991 37924 17003 37927
rect 18340 37924 18368 37964
rect 19426 37952 19432 37964
rect 19484 37952 19490 38004
rect 21174 37952 21180 38004
rect 21232 37992 21238 38004
rect 21821 37995 21879 38001
rect 21821 37992 21833 37995
rect 21232 37964 21833 37992
rect 21232 37952 21238 37964
rect 21821 37961 21833 37964
rect 21867 37961 21879 37995
rect 25222 37992 25228 38004
rect 25183 37964 25228 37992
rect 21821 37955 21879 37961
rect 25222 37952 25228 37964
rect 25280 37952 25286 38004
rect 25409 37995 25467 38001
rect 25409 37961 25421 37995
rect 25455 37992 25467 37995
rect 26050 37992 26056 38004
rect 25455 37964 26056 37992
rect 25455 37961 25467 37964
rect 25409 37955 25467 37961
rect 26050 37952 26056 37964
rect 26108 37952 26114 38004
rect 30282 37992 30288 38004
rect 26988 37964 30288 37992
rect 16991 37896 18368 37924
rect 18417 37927 18475 37933
rect 16991 37893 17003 37896
rect 16945 37887 17003 37893
rect 18417 37893 18429 37927
rect 18463 37893 18475 37927
rect 18417 37887 18475 37893
rect 17402 37856 17408 37868
rect 17363 37828 17408 37856
rect 17402 37816 17408 37828
rect 17460 37816 17466 37868
rect 17681 37859 17739 37865
rect 17681 37825 17693 37859
rect 17727 37856 17739 37859
rect 17770 37856 17776 37868
rect 17727 37828 17776 37856
rect 17727 37825 17739 37828
rect 17681 37819 17739 37825
rect 17770 37816 17776 37828
rect 17828 37816 17834 37868
rect 18432 37788 18460 37887
rect 18506 37884 18512 37936
rect 18564 37924 18570 37936
rect 18617 37927 18675 37933
rect 18617 37924 18629 37927
rect 18564 37896 18629 37924
rect 18564 37884 18570 37896
rect 18617 37893 18629 37896
rect 18663 37893 18675 37927
rect 18617 37887 18675 37893
rect 20898 37884 20904 37936
rect 20956 37924 20962 37936
rect 20956 37896 21220 37924
rect 20956 37884 20962 37896
rect 19981 37859 20039 37865
rect 19981 37856 19993 37859
rect 18800 37828 19993 37856
rect 18690 37788 18696 37800
rect 16546 37760 18696 37788
rect 16022 37652 16028 37664
rect 15983 37624 16028 37652
rect 16022 37612 16028 37624
rect 16080 37652 16086 37664
rect 16546 37652 16574 37760
rect 18690 37748 18696 37760
rect 18748 37748 18754 37800
rect 18800 37729 18828 37828
rect 19981 37825 19993 37828
rect 20027 37856 20039 37859
rect 20070 37856 20076 37868
rect 20027 37828 20076 37856
rect 20027 37825 20039 37828
rect 19981 37819 20039 37825
rect 20070 37816 20076 37828
rect 20128 37816 20134 37868
rect 20162 37816 20168 37868
rect 20220 37856 20226 37868
rect 21082 37856 21088 37868
rect 20220 37828 20265 37856
rect 21043 37828 21088 37856
rect 20220 37816 20226 37828
rect 21082 37816 21088 37828
rect 21140 37816 21146 37868
rect 21192 37856 21220 37896
rect 21358 37884 21364 37936
rect 21416 37924 21422 37936
rect 21416 37896 26004 37924
rect 21416 37884 21422 37896
rect 22005 37859 22063 37865
rect 22005 37856 22017 37859
rect 21192 37828 22017 37856
rect 22005 37825 22017 37828
rect 22051 37825 22063 37859
rect 22005 37819 22063 37825
rect 22097 37859 22155 37865
rect 22097 37825 22109 37859
rect 22143 37856 22155 37859
rect 22830 37856 22836 37868
rect 22143 37828 22836 37856
rect 22143 37825 22155 37828
rect 22097 37819 22155 37825
rect 20625 37791 20683 37797
rect 20625 37788 20637 37791
rect 19996 37760 20637 37788
rect 19996 37729 20024 37760
rect 20625 37757 20637 37760
rect 20671 37788 20683 37791
rect 20714 37788 20720 37800
rect 20671 37760 20720 37788
rect 20671 37757 20683 37760
rect 20625 37751 20683 37757
rect 20714 37748 20720 37760
rect 20772 37748 20778 37800
rect 20993 37791 21051 37797
rect 20993 37757 21005 37791
rect 21039 37788 21051 37791
rect 21266 37788 21272 37800
rect 21039 37760 21272 37788
rect 21039 37757 21051 37760
rect 20993 37751 21051 37757
rect 21266 37748 21272 37760
rect 21324 37748 21330 37800
rect 21818 37788 21824 37800
rect 21779 37760 21824 37788
rect 21818 37748 21824 37760
rect 21876 37748 21882 37800
rect 18785 37723 18843 37729
rect 18785 37689 18797 37723
rect 18831 37689 18843 37723
rect 18785 37683 18843 37689
rect 19981 37723 20039 37729
rect 19981 37689 19993 37723
rect 20027 37689 20039 37723
rect 19981 37683 20039 37689
rect 21082 37680 21088 37732
rect 21140 37720 21146 37732
rect 22112 37720 22140 37819
rect 22830 37816 22836 37828
rect 22888 37816 22894 37868
rect 23382 37856 23388 37868
rect 23343 37828 23388 37856
rect 23382 37816 23388 37828
rect 23440 37816 23446 37868
rect 23569 37859 23627 37865
rect 23569 37825 23581 37859
rect 23615 37825 23627 37859
rect 23569 37819 23627 37825
rect 22462 37748 22468 37800
rect 22520 37788 22526 37800
rect 23584 37788 23612 37819
rect 24302 37816 24308 37868
rect 24360 37856 24366 37868
rect 24489 37859 24547 37865
rect 24489 37856 24501 37859
rect 24360 37828 24501 37856
rect 24360 37816 24366 37828
rect 24489 37825 24501 37828
rect 24535 37825 24547 37859
rect 24489 37819 24547 37825
rect 24762 37816 24768 37868
rect 24820 37856 24826 37868
rect 25133 37859 25191 37865
rect 25133 37856 25145 37859
rect 24820 37828 25145 37856
rect 24820 37816 24826 37828
rect 25133 37825 25145 37828
rect 25179 37856 25191 37859
rect 25406 37856 25412 37868
rect 25179 37828 25412 37856
rect 25179 37825 25191 37828
rect 25133 37819 25191 37825
rect 25406 37816 25412 37828
rect 25464 37816 25470 37868
rect 25976 37865 26004 37896
rect 25501 37859 25559 37865
rect 25501 37825 25513 37859
rect 25547 37825 25559 37859
rect 25501 37819 25559 37825
rect 25961 37859 26019 37865
rect 25961 37825 25973 37859
rect 26007 37825 26019 37859
rect 26418 37856 26424 37868
rect 26379 37828 26424 37856
rect 25961 37819 26019 37825
rect 24670 37788 24676 37800
rect 22520 37760 24676 37788
rect 22520 37748 22526 37760
rect 24670 37748 24676 37760
rect 24728 37748 24734 37800
rect 25314 37788 25320 37800
rect 25275 37760 25320 37788
rect 25314 37748 25320 37760
rect 25372 37748 25378 37800
rect 25516 37788 25544 37819
rect 26418 37816 26424 37828
rect 26476 37816 26482 37868
rect 26988 37865 27016 37964
rect 30282 37952 30288 37964
rect 30340 37952 30346 38004
rect 30834 37992 30840 38004
rect 30392 37964 30840 37992
rect 30101 37927 30159 37933
rect 30101 37893 30113 37927
rect 30147 37924 30159 37927
rect 30392 37924 30420 37964
rect 30834 37952 30840 37964
rect 30892 37952 30898 38004
rect 33321 37995 33379 38001
rect 33321 37961 33333 37995
rect 33367 37992 33379 37995
rect 33410 37992 33416 38004
rect 33367 37964 33416 37992
rect 33367 37961 33379 37964
rect 33321 37955 33379 37961
rect 33410 37952 33416 37964
rect 33468 37952 33474 38004
rect 33594 37952 33600 38004
rect 33652 37992 33658 38004
rect 34057 37995 34115 38001
rect 34057 37992 34069 37995
rect 33652 37964 34069 37992
rect 33652 37952 33658 37964
rect 34057 37961 34069 37964
rect 34103 37961 34115 37995
rect 34057 37955 34115 37961
rect 35158 37952 35164 38004
rect 35216 37992 35222 38004
rect 35437 37995 35495 38001
rect 35437 37992 35449 37995
rect 35216 37964 35449 37992
rect 35216 37952 35222 37964
rect 35437 37961 35449 37964
rect 35483 37961 35495 37995
rect 35437 37955 35495 37961
rect 35526 37952 35532 38004
rect 35584 37992 35590 38004
rect 36173 37995 36231 38001
rect 36173 37992 36185 37995
rect 35584 37964 36185 37992
rect 35584 37952 35590 37964
rect 36173 37961 36185 37964
rect 36219 37961 36231 37995
rect 36173 37955 36231 37961
rect 37274 37924 37280 37936
rect 30147 37896 30420 37924
rect 36096 37896 37280 37924
rect 30147 37893 30159 37896
rect 30101 37887 30159 37893
rect 26973 37859 27031 37865
rect 26973 37825 26985 37859
rect 27019 37825 27031 37859
rect 26973 37819 27031 37825
rect 27062 37816 27068 37868
rect 27120 37856 27126 37868
rect 27229 37859 27287 37865
rect 27229 37856 27241 37859
rect 27120 37828 27241 37856
rect 27120 37816 27126 37828
rect 27229 37825 27241 37828
rect 27275 37825 27287 37859
rect 30837 37859 30895 37865
rect 27229 37819 27287 37825
rect 26053 37791 26111 37797
rect 26053 37788 26065 37791
rect 25516 37760 26065 37788
rect 26053 37757 26065 37760
rect 26099 37757 26111 37791
rect 26053 37751 26111 37757
rect 26283 37791 26341 37797
rect 26283 37757 26295 37791
rect 26329 37788 26341 37791
rect 26694 37788 26700 37800
rect 26329 37760 26700 37788
rect 26329 37757 26341 37760
rect 26283 37751 26341 37757
rect 26694 37748 26700 37760
rect 26752 37748 26758 37800
rect 28350 37748 28356 37800
rect 28408 37788 28414 37800
rect 28997 37791 29055 37797
rect 28997 37788 29009 37791
rect 28408 37760 29009 37788
rect 28408 37748 28414 37760
rect 28997 37757 29009 37760
rect 29043 37757 29055 37791
rect 28997 37751 29055 37757
rect 30466 37748 30472 37800
rect 30524 37788 30530 37800
rect 30760 37788 30788 37842
rect 30837 37825 30849 37859
rect 30883 37856 30895 37859
rect 31018 37856 31024 37868
rect 30883 37828 31024 37856
rect 30883 37825 30895 37828
rect 30837 37819 30895 37825
rect 31018 37816 31024 37828
rect 31076 37856 31082 37868
rect 31389 37859 31447 37865
rect 31389 37856 31401 37859
rect 31076 37828 31401 37856
rect 31076 37816 31082 37828
rect 31389 37825 31401 37828
rect 31435 37856 31447 37859
rect 31570 37856 31576 37868
rect 31435 37828 31576 37856
rect 31435 37825 31447 37828
rect 31389 37819 31447 37825
rect 31570 37816 31576 37828
rect 31628 37856 31634 37868
rect 32030 37856 32036 37868
rect 31628 37828 32036 37856
rect 31628 37816 31634 37828
rect 32030 37816 32036 37828
rect 32088 37816 32094 37868
rect 32582 37856 32588 37868
rect 32543 37828 32588 37856
rect 32582 37816 32588 37828
rect 32640 37816 32646 37868
rect 33042 37856 33048 37868
rect 33003 37828 33048 37856
rect 33042 37816 33048 37828
rect 33100 37816 33106 37868
rect 33137 37859 33195 37865
rect 33137 37825 33149 37859
rect 33183 37856 33195 37859
rect 33226 37856 33232 37868
rect 33183 37828 33232 37856
rect 33183 37825 33195 37828
rect 33137 37819 33195 37825
rect 33226 37816 33232 37828
rect 33284 37816 33290 37868
rect 33962 37856 33968 37868
rect 33923 37828 33968 37856
rect 33962 37816 33968 37828
rect 34020 37816 34026 37868
rect 34149 37859 34207 37865
rect 34149 37825 34161 37859
rect 34195 37856 34207 37859
rect 34606 37856 34612 37868
rect 34195 37828 34612 37856
rect 34195 37825 34207 37828
rect 34149 37819 34207 37825
rect 34606 37816 34612 37828
rect 34664 37816 34670 37868
rect 35529 37859 35587 37865
rect 35529 37825 35541 37859
rect 35575 37856 35587 37859
rect 35802 37856 35808 37868
rect 35575 37828 35808 37856
rect 35575 37825 35587 37828
rect 35529 37819 35587 37825
rect 35802 37816 35808 37828
rect 35860 37816 35866 37868
rect 36096 37865 36124 37896
rect 37274 37884 37280 37896
rect 37332 37884 37338 37936
rect 36081 37859 36139 37865
rect 36081 37825 36093 37859
rect 36127 37825 36139 37859
rect 36081 37819 36139 37825
rect 36265 37859 36323 37865
rect 36265 37825 36277 37859
rect 36311 37856 36323 37859
rect 36446 37856 36452 37868
rect 36311 37828 36452 37856
rect 36311 37825 36323 37828
rect 36265 37819 36323 37825
rect 36446 37816 36452 37828
rect 36504 37816 36510 37868
rect 37734 37816 37740 37868
rect 37792 37865 37798 37868
rect 37792 37859 37825 37865
rect 37813 37825 37825 37859
rect 37792 37819 37825 37825
rect 37921 37859 37979 37865
rect 37921 37825 37933 37859
rect 37967 37856 37979 37859
rect 38746 37856 38752 37868
rect 37967 37828 38752 37856
rect 37967 37825 37979 37828
rect 37921 37819 37979 37825
rect 37792 37816 37798 37819
rect 38746 37816 38752 37828
rect 38804 37816 38810 37868
rect 31938 37788 31944 37800
rect 30524 37760 31944 37788
rect 30524 37748 30530 37760
rect 31938 37748 31944 37760
rect 31996 37748 32002 37800
rect 33321 37791 33379 37797
rect 33321 37788 33333 37791
rect 33152 37760 33333 37788
rect 33152 37732 33180 37760
rect 33321 37757 33333 37760
rect 33367 37757 33379 37791
rect 33321 37751 33379 37757
rect 21140 37692 22140 37720
rect 23569 37723 23627 37729
rect 21140 37680 21146 37692
rect 23569 37689 23581 37723
rect 23615 37720 23627 37723
rect 23615 37692 24256 37720
rect 23615 37689 23627 37692
rect 23569 37683 23627 37689
rect 16080 37624 16574 37652
rect 17865 37655 17923 37661
rect 16080 37612 16086 37624
rect 17865 37621 17877 37655
rect 17911 37652 17923 37655
rect 18506 37652 18512 37664
rect 17911 37624 18512 37652
rect 17911 37621 17923 37624
rect 17865 37615 17923 37621
rect 18506 37612 18512 37624
rect 18564 37652 18570 37664
rect 18601 37655 18659 37661
rect 18601 37652 18613 37655
rect 18564 37624 18613 37652
rect 18564 37612 18570 37624
rect 18601 37621 18613 37624
rect 18647 37621 18659 37655
rect 19702 37652 19708 37664
rect 19663 37624 19708 37652
rect 18601 37615 18659 37621
rect 19702 37612 19708 37624
rect 19760 37612 19766 37664
rect 21269 37655 21327 37661
rect 21269 37621 21281 37655
rect 21315 37652 21327 37655
rect 21450 37652 21456 37664
rect 21315 37624 21456 37652
rect 21315 37621 21327 37624
rect 21269 37615 21327 37621
rect 21450 37612 21456 37624
rect 21508 37612 21514 37664
rect 22925 37655 22983 37661
rect 22925 37621 22937 37655
rect 22971 37652 22983 37655
rect 23842 37652 23848 37664
rect 22971 37624 23848 37652
rect 22971 37621 22983 37624
rect 22925 37615 22983 37621
rect 23842 37612 23848 37624
rect 23900 37612 23906 37664
rect 24026 37652 24032 37664
rect 23987 37624 24032 37652
rect 24026 37612 24032 37624
rect 24084 37612 24090 37664
rect 24228 37661 24256 37692
rect 26602 37680 26608 37732
rect 26660 37720 26666 37732
rect 26660 37692 26832 37720
rect 26660 37680 26666 37692
rect 24213 37655 24271 37661
rect 24213 37621 24225 37655
rect 24259 37652 24271 37655
rect 24670 37652 24676 37664
rect 24259 37624 24676 37652
rect 24259 37621 24271 37624
rect 24213 37615 24271 37621
rect 24670 37612 24676 37624
rect 24728 37612 24734 37664
rect 26145 37655 26203 37661
rect 26145 37621 26157 37655
rect 26191 37652 26203 37655
rect 26694 37652 26700 37664
rect 26191 37624 26700 37652
rect 26191 37621 26203 37624
rect 26145 37615 26203 37621
rect 26694 37612 26700 37624
rect 26752 37612 26758 37664
rect 26804 37652 26832 37692
rect 31662 37680 31668 37732
rect 31720 37720 31726 37732
rect 33134 37720 33140 37732
rect 31720 37692 33140 37720
rect 31720 37680 31726 37692
rect 33134 37680 33140 37692
rect 33192 37680 33198 37732
rect 37550 37720 37556 37732
rect 37511 37692 37556 37720
rect 37550 37680 37556 37692
rect 37608 37680 37614 37732
rect 28353 37655 28411 37661
rect 28353 37652 28365 37655
rect 26804 37624 28365 37652
rect 28353 37621 28365 37624
rect 28399 37621 28411 37655
rect 32122 37652 32128 37664
rect 32083 37624 32128 37652
rect 28353 37615 28411 37621
rect 32122 37612 32128 37624
rect 32180 37612 32186 37664
rect 32490 37652 32496 37664
rect 32451 37624 32496 37652
rect 32490 37612 32496 37624
rect 32548 37612 32554 37664
rect 33594 37612 33600 37664
rect 33652 37652 33658 37664
rect 34146 37652 34152 37664
rect 33652 37624 34152 37652
rect 33652 37612 33658 37624
rect 34146 37612 34152 37624
rect 34204 37652 34210 37664
rect 34609 37655 34667 37661
rect 34609 37652 34621 37655
rect 34204 37624 34621 37652
rect 34204 37612 34210 37624
rect 34609 37621 34621 37624
rect 34655 37621 34667 37655
rect 38378 37652 38384 37664
rect 38339 37624 38384 37652
rect 34609 37615 34667 37621
rect 38378 37612 38384 37624
rect 38436 37652 38442 37664
rect 38933 37655 38991 37661
rect 38933 37652 38945 37655
rect 38436 37624 38945 37652
rect 38436 37612 38442 37624
rect 38933 37621 38945 37624
rect 38979 37621 38991 37655
rect 38933 37615 38991 37621
rect 1104 37562 54372 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 54372 37562
rect 1104 37488 54372 37510
rect 16390 37408 16396 37460
rect 16448 37448 16454 37460
rect 16577 37451 16635 37457
rect 16577 37448 16589 37451
rect 16448 37420 16589 37448
rect 16448 37408 16454 37420
rect 16577 37417 16589 37420
rect 16623 37417 16635 37451
rect 17494 37448 17500 37460
rect 17455 37420 17500 37448
rect 16577 37411 16635 37417
rect 17494 37408 17500 37420
rect 17552 37408 17558 37460
rect 17589 37451 17647 37457
rect 17589 37417 17601 37451
rect 17635 37448 17647 37451
rect 18230 37448 18236 37460
rect 17635 37420 18236 37448
rect 17635 37417 17647 37420
rect 17589 37411 17647 37417
rect 18230 37408 18236 37420
rect 18288 37408 18294 37460
rect 18693 37451 18751 37457
rect 18693 37417 18705 37451
rect 18739 37448 18751 37451
rect 19702 37448 19708 37460
rect 18739 37420 19708 37448
rect 18739 37417 18751 37420
rect 18693 37411 18751 37417
rect 19702 37408 19708 37420
rect 19760 37408 19766 37460
rect 20806 37408 20812 37460
rect 20864 37448 20870 37460
rect 23845 37451 23903 37457
rect 20864 37420 20944 37448
rect 20864 37408 20870 37420
rect 17310 37340 17316 37392
rect 17368 37380 17374 37392
rect 17405 37383 17463 37389
rect 17405 37380 17417 37383
rect 17368 37352 17417 37380
rect 17368 37340 17374 37352
rect 17405 37349 17417 37352
rect 17451 37380 17463 37383
rect 17770 37380 17776 37392
rect 17451 37352 17776 37380
rect 17451 37349 17463 37352
rect 17405 37343 17463 37349
rect 17770 37340 17776 37352
rect 17828 37340 17834 37392
rect 18322 37340 18328 37392
rect 18380 37380 18386 37392
rect 19245 37383 19303 37389
rect 19245 37380 19257 37383
rect 18380 37352 19257 37380
rect 18380 37340 18386 37352
rect 19245 37349 19257 37352
rect 19291 37349 19303 37383
rect 19245 37343 19303 37349
rect 16022 37312 16028 37324
rect 15983 37284 16028 37312
rect 16022 37272 16028 37284
rect 16080 37272 16086 37324
rect 17862 37312 17868 37324
rect 17823 37284 17868 37312
rect 17862 37272 17868 37284
rect 17920 37272 17926 37324
rect 19426 37272 19432 37324
rect 19484 37312 19490 37324
rect 19720 37312 19748 37408
rect 20257 37383 20315 37389
rect 20257 37349 20269 37383
rect 20303 37380 20315 37383
rect 20303 37352 20852 37380
rect 20303 37349 20315 37352
rect 20257 37343 20315 37349
rect 19484 37284 19656 37312
rect 19720 37284 20300 37312
rect 19484 37272 19490 37284
rect 17129 37247 17187 37253
rect 17129 37213 17141 37247
rect 17175 37244 17187 37247
rect 17218 37244 17224 37256
rect 17175 37216 17224 37244
rect 17175 37213 17187 37216
rect 17129 37207 17187 37213
rect 17218 37204 17224 37216
rect 17276 37204 17282 37256
rect 18414 37244 18420 37256
rect 18375 37216 18420 37244
rect 18414 37204 18420 37216
rect 18472 37204 18478 37256
rect 18690 37244 18696 37256
rect 18603 37216 18696 37244
rect 18690 37204 18696 37216
rect 18748 37244 18754 37256
rect 19628 37253 19656 37284
rect 19613 37247 19671 37253
rect 18748 37216 19564 37244
rect 18748 37204 18754 37216
rect 19242 37136 19248 37188
rect 19300 37176 19306 37188
rect 19429 37179 19487 37185
rect 19429 37176 19441 37179
rect 19300 37148 19441 37176
rect 19300 37136 19306 37148
rect 19429 37145 19441 37148
rect 19475 37145 19487 37179
rect 19536 37176 19564 37216
rect 19613 37213 19625 37247
rect 19659 37213 19671 37247
rect 20070 37244 20076 37256
rect 20031 37216 20076 37244
rect 19613 37207 19671 37213
rect 20070 37204 20076 37216
rect 20128 37204 20134 37256
rect 20272 37253 20300 37284
rect 20824 37253 20852 37352
rect 20916 37312 20944 37420
rect 23845 37417 23857 37451
rect 23891 37448 23903 37451
rect 23934 37448 23940 37460
rect 23891 37420 23940 37448
rect 23891 37417 23903 37420
rect 23845 37411 23903 37417
rect 23934 37408 23940 37420
rect 23992 37408 23998 37460
rect 26602 37408 26608 37460
rect 26660 37448 26666 37460
rect 26881 37451 26939 37457
rect 26881 37448 26893 37451
rect 26660 37420 26893 37448
rect 26660 37408 26666 37420
rect 26881 37417 26893 37420
rect 26927 37417 26939 37451
rect 26881 37411 26939 37417
rect 29914 37408 29920 37460
rect 29972 37448 29978 37460
rect 30837 37451 30895 37457
rect 30837 37448 30849 37451
rect 29972 37420 30849 37448
rect 29972 37408 29978 37420
rect 30837 37417 30849 37420
rect 30883 37417 30895 37451
rect 33502 37448 33508 37460
rect 33463 37420 33508 37448
rect 30837 37411 30895 37417
rect 33502 37408 33508 37420
rect 33560 37408 33566 37460
rect 34698 37408 34704 37460
rect 34756 37448 34762 37460
rect 35986 37448 35992 37460
rect 34756 37420 35992 37448
rect 34756 37408 34762 37420
rect 35986 37408 35992 37420
rect 36044 37408 36050 37460
rect 36354 37448 36360 37460
rect 36315 37420 36360 37448
rect 36354 37408 36360 37420
rect 36412 37408 36418 37460
rect 36630 37408 36636 37460
rect 36688 37448 36694 37460
rect 38194 37448 38200 37460
rect 36688 37420 37688 37448
rect 38155 37420 38200 37448
rect 36688 37408 36694 37420
rect 22370 37380 22376 37392
rect 22283 37352 22376 37380
rect 22370 37340 22376 37352
rect 22428 37380 22434 37392
rect 23658 37380 23664 37392
rect 22428 37352 23664 37380
rect 22428 37340 22434 37352
rect 23658 37340 23664 37352
rect 23716 37340 23722 37392
rect 24302 37340 24308 37392
rect 24360 37380 24366 37392
rect 24360 37352 25636 37380
rect 24360 37340 24366 37352
rect 21821 37315 21879 37321
rect 20916 37284 21036 37312
rect 20257 37247 20315 37253
rect 20257 37213 20269 37247
rect 20303 37213 20315 37247
rect 20257 37207 20315 37213
rect 20809 37247 20867 37253
rect 20809 37213 20821 37247
rect 20855 37244 20867 37247
rect 20898 37244 20904 37256
rect 20855 37216 20904 37244
rect 20855 37213 20867 37216
rect 20809 37207 20867 37213
rect 20898 37204 20904 37216
rect 20956 37204 20962 37256
rect 21008 37253 21036 37284
rect 21821 37281 21833 37315
rect 21867 37312 21879 37315
rect 22186 37312 22192 37324
rect 21867 37284 22192 37312
rect 21867 37281 21879 37284
rect 21821 37275 21879 37281
rect 22186 37272 22192 37284
rect 22244 37272 22250 37324
rect 22278 37272 22284 37324
rect 22336 37312 22342 37324
rect 23382 37312 23388 37324
rect 22336 37284 23388 37312
rect 22336 37272 22342 37284
rect 23032 37253 23060 37284
rect 23382 37272 23388 37284
rect 23440 37272 23446 37324
rect 23753 37315 23811 37321
rect 23753 37281 23765 37315
rect 23799 37312 23811 37315
rect 24026 37312 24032 37324
rect 23799 37284 24032 37312
rect 23799 37281 23811 37284
rect 23753 37275 23811 37281
rect 24026 37272 24032 37284
rect 24084 37272 24090 37324
rect 20993 37247 21051 37253
rect 20993 37213 21005 37247
rect 21039 37213 21051 37247
rect 22833 37247 22891 37253
rect 22833 37244 22845 37247
rect 20993 37207 21051 37213
rect 22480 37216 22845 37244
rect 22480 37188 22508 37216
rect 22833 37213 22845 37216
rect 22879 37213 22891 37247
rect 22833 37207 22891 37213
rect 23017 37247 23075 37253
rect 23017 37213 23029 37247
rect 23063 37213 23075 37247
rect 23017 37207 23075 37213
rect 23845 37247 23903 37253
rect 23845 37213 23857 37247
rect 23891 37244 23903 37247
rect 24486 37244 24492 37256
rect 23891 37216 24492 37244
rect 23891 37213 23903 37216
rect 23845 37207 23903 37213
rect 24486 37204 24492 37216
rect 24544 37204 24550 37256
rect 24670 37244 24676 37256
rect 24631 37216 24676 37244
rect 24670 37204 24676 37216
rect 24728 37204 24734 37256
rect 24765 37247 24823 37253
rect 24765 37213 24777 37247
rect 24811 37213 24823 37247
rect 24765 37207 24823 37213
rect 19978 37176 19984 37188
rect 19536 37148 19984 37176
rect 19429 37139 19487 37145
rect 19978 37136 19984 37148
rect 20036 37176 20042 37188
rect 22462 37176 22468 37188
rect 20036 37148 22468 37176
rect 20036 37136 20042 37148
rect 22462 37136 22468 37148
rect 22520 37136 22526 37188
rect 22925 37179 22983 37185
rect 22925 37145 22937 37179
rect 22971 37176 22983 37179
rect 24302 37176 24308 37188
rect 22971 37148 24308 37176
rect 22971 37145 22983 37148
rect 22925 37139 22983 37145
rect 24302 37136 24308 37148
rect 24360 37136 24366 37188
rect 24780 37176 24808 37207
rect 24854 37204 24860 37256
rect 24912 37244 24918 37256
rect 25056 37253 25084 37352
rect 25608 37312 25636 37352
rect 26694 37340 26700 37392
rect 26752 37380 26758 37392
rect 27062 37380 27068 37392
rect 26752 37352 27068 37380
rect 26752 37340 26758 37352
rect 27062 37340 27068 37352
rect 27120 37340 27126 37392
rect 29822 37380 29828 37392
rect 29783 37352 29828 37380
rect 29822 37340 29828 37352
rect 29880 37340 29886 37392
rect 32398 37380 32404 37392
rect 29932 37352 32404 37380
rect 25608 37284 25912 37312
rect 25041 37247 25099 37253
rect 24912 37216 24957 37244
rect 24912 37204 24918 37216
rect 25041 37213 25053 37247
rect 25087 37213 25099 37247
rect 25041 37207 25099 37213
rect 25406 37204 25412 37256
rect 25464 37244 25470 37256
rect 25777 37247 25835 37253
rect 25777 37244 25789 37247
rect 25464 37216 25789 37244
rect 25464 37204 25470 37216
rect 25777 37213 25789 37216
rect 25823 37213 25835 37247
rect 25777 37207 25835 37213
rect 25130 37176 25136 37188
rect 24780 37148 25136 37176
rect 25130 37136 25136 37148
rect 25188 37136 25194 37188
rect 25222 37136 25228 37188
rect 25280 37176 25286 37188
rect 25501 37179 25559 37185
rect 25501 37176 25513 37179
rect 25280 37148 25513 37176
rect 25280 37136 25286 37148
rect 25501 37145 25513 37148
rect 25547 37145 25559 37179
rect 25501 37139 25559 37145
rect 25685 37179 25743 37185
rect 25685 37145 25697 37179
rect 25731 37176 25743 37179
rect 25884 37176 25912 37284
rect 26418 37272 26424 37324
rect 26476 37312 26482 37324
rect 29932 37312 29960 37352
rect 32398 37340 32404 37352
rect 32456 37340 32462 37392
rect 34149 37383 34207 37389
rect 34149 37349 34161 37383
rect 34195 37380 34207 37383
rect 34606 37380 34612 37392
rect 34195 37352 34612 37380
rect 34195 37349 34207 37352
rect 34149 37343 34207 37349
rect 34606 37340 34612 37352
rect 34664 37340 34670 37392
rect 34882 37340 34888 37392
rect 34940 37380 34946 37392
rect 35345 37383 35403 37389
rect 35345 37380 35357 37383
rect 34940 37352 35357 37380
rect 34940 37340 34946 37352
rect 35345 37349 35357 37352
rect 35391 37349 35403 37383
rect 35345 37343 35403 37349
rect 37182 37340 37188 37392
rect 37240 37380 37246 37392
rect 37277 37383 37335 37389
rect 37277 37380 37289 37383
rect 37240 37352 37289 37380
rect 37240 37340 37246 37352
rect 37277 37349 37289 37352
rect 37323 37349 37335 37383
rect 37277 37343 37335 37349
rect 37369 37383 37427 37389
rect 37369 37349 37381 37383
rect 37415 37380 37427 37383
rect 37550 37380 37556 37392
rect 37415 37352 37556 37380
rect 37415 37349 37427 37352
rect 37369 37343 37427 37349
rect 26476 37284 29960 37312
rect 26476 37272 26482 37284
rect 30926 37272 30932 37324
rect 30984 37312 30990 37324
rect 30984 37284 31340 37312
rect 30984 37272 30990 37284
rect 27154 37244 27160 37256
rect 26712 37216 27160 37244
rect 26712 37185 26740 37216
rect 27154 37204 27160 37216
rect 27212 37244 27218 37256
rect 27522 37244 27528 37256
rect 27212 37216 27528 37244
rect 27212 37204 27218 37216
rect 27522 37204 27528 37216
rect 27580 37204 27586 37256
rect 27706 37204 27712 37256
rect 27764 37244 27770 37256
rect 28350 37244 28356 37256
rect 27764 37216 28356 37244
rect 27764 37204 27770 37216
rect 28350 37204 28356 37216
rect 28408 37204 28414 37256
rect 28534 37244 28540 37256
rect 28495 37216 28540 37244
rect 28534 37204 28540 37216
rect 28592 37204 28598 37256
rect 29730 37244 29736 37256
rect 29691 37216 29736 37244
rect 29730 37204 29736 37216
rect 29788 37204 29794 37256
rect 29914 37244 29920 37256
rect 29875 37216 29920 37244
rect 29914 37204 29920 37216
rect 29972 37204 29978 37256
rect 30009 37247 30067 37253
rect 30009 37213 30021 37247
rect 30055 37213 30067 37247
rect 30009 37207 30067 37213
rect 25731 37148 25912 37176
rect 26697 37179 26755 37185
rect 25731 37145 25743 37148
rect 25685 37139 25743 37145
rect 26697 37145 26709 37179
rect 26743 37145 26755 37179
rect 26697 37139 26755 37145
rect 26878 37136 26884 37188
rect 26936 37185 26942 37188
rect 26936 37179 26955 37185
rect 26943 37145 26955 37179
rect 28902 37176 28908 37188
rect 26936 37139 26955 37145
rect 28000 37148 28908 37176
rect 26936 37136 26942 37139
rect 28000 37120 28028 37148
rect 28902 37136 28908 37148
rect 28960 37136 28966 37188
rect 29638 37136 29644 37188
rect 29696 37176 29702 37188
rect 30024 37176 30052 37207
rect 30098 37204 30104 37256
rect 30156 37244 30162 37256
rect 30193 37247 30251 37253
rect 30193 37244 30205 37247
rect 30156 37216 30205 37244
rect 30156 37204 30162 37216
rect 30193 37213 30205 37216
rect 30239 37213 30251 37247
rect 30193 37207 30251 37213
rect 30650 37204 30656 37256
rect 30708 37244 30714 37256
rect 31312 37253 31340 37284
rect 32582 37272 32588 37324
rect 32640 37312 32646 37324
rect 37001 37315 37059 37321
rect 37001 37312 37013 37315
rect 32640 37284 37013 37312
rect 32640 37272 32646 37284
rect 37001 37281 37013 37284
rect 37047 37281 37059 37315
rect 37001 37275 37059 37281
rect 31021 37247 31079 37253
rect 31021 37244 31033 37247
rect 30708 37216 31033 37244
rect 30708 37204 30714 37216
rect 31021 37213 31033 37216
rect 31067 37213 31079 37247
rect 31021 37207 31079 37213
rect 31297 37247 31355 37253
rect 31297 37213 31309 37247
rect 31343 37244 31355 37247
rect 31478 37244 31484 37256
rect 31343 37216 31484 37244
rect 31343 37213 31355 37216
rect 31297 37207 31355 37213
rect 29696 37148 30052 37176
rect 29696 37136 29702 37148
rect 16942 37068 16948 37120
rect 17000 37108 17006 37120
rect 17221 37111 17279 37117
rect 17221 37108 17233 37111
rect 17000 37080 17233 37108
rect 17000 37068 17006 37080
rect 17221 37077 17233 37080
rect 17267 37077 17279 37111
rect 18506 37108 18512 37120
rect 18467 37080 18512 37108
rect 17221 37071 17279 37077
rect 18506 37068 18512 37080
rect 18564 37068 18570 37120
rect 20990 37108 20996 37120
rect 20951 37080 20996 37108
rect 20990 37068 20996 37080
rect 21048 37068 21054 37120
rect 23477 37111 23535 37117
rect 23477 37077 23489 37111
rect 23523 37108 23535 37111
rect 24210 37108 24216 37120
rect 23523 37080 24216 37108
rect 23523 37077 23535 37080
rect 23477 37071 23535 37077
rect 24210 37068 24216 37080
rect 24268 37068 24274 37120
rect 24394 37108 24400 37120
rect 24355 37080 24400 37108
rect 24394 37068 24400 37080
rect 24452 37068 24458 37120
rect 24578 37068 24584 37120
rect 24636 37108 24642 37120
rect 25599 37111 25657 37117
rect 25599 37108 25611 37111
rect 24636 37080 25611 37108
rect 24636 37068 24642 37080
rect 25599 37077 25611 37080
rect 25645 37077 25657 37111
rect 25599 37071 25657 37077
rect 27617 37111 27675 37117
rect 27617 37077 27629 37111
rect 27663 37108 27675 37111
rect 27982 37108 27988 37120
rect 27663 37080 27988 37108
rect 27663 37077 27675 37080
rect 27617 37071 27675 37077
rect 27982 37068 27988 37080
rect 28040 37068 28046 37120
rect 28445 37111 28503 37117
rect 28445 37077 28457 37111
rect 28491 37108 28503 37111
rect 28718 37108 28724 37120
rect 28491 37080 28724 37108
rect 28491 37077 28503 37080
rect 28445 37071 28503 37077
rect 28718 37068 28724 37080
rect 28776 37068 28782 37120
rect 29549 37111 29607 37117
rect 29549 37077 29561 37111
rect 29595 37108 29607 37111
rect 30742 37108 30748 37120
rect 29595 37080 30748 37108
rect 29595 37077 29607 37080
rect 29549 37071 29607 37077
rect 30742 37068 30748 37080
rect 30800 37068 30806 37120
rect 31036 37108 31064 37207
rect 31478 37204 31484 37216
rect 31536 37204 31542 37256
rect 31754 37244 31760 37256
rect 31715 37216 31760 37244
rect 31754 37204 31760 37216
rect 31812 37244 31818 37256
rect 32214 37244 32220 37256
rect 31812 37216 32220 37244
rect 31812 37204 31818 37216
rect 32214 37204 32220 37216
rect 32272 37244 32278 37256
rect 32861 37247 32919 37253
rect 32861 37244 32873 37247
rect 32272 37216 32873 37244
rect 32272 37204 32278 37216
rect 32861 37213 32873 37216
rect 32907 37213 32919 37247
rect 32861 37207 32919 37213
rect 33965 37247 34023 37253
rect 33965 37213 33977 37247
rect 34011 37213 34023 37247
rect 33965 37207 34023 37213
rect 34149 37247 34207 37253
rect 34149 37213 34161 37247
rect 34195 37244 34207 37247
rect 34238 37244 34244 37256
rect 34195 37216 34244 37244
rect 34195 37213 34207 37216
rect 34149 37207 34207 37213
rect 31205 37179 31263 37185
rect 31205 37145 31217 37179
rect 31251 37176 31263 37179
rect 32122 37176 32128 37188
rect 31251 37148 32128 37176
rect 31251 37145 31263 37148
rect 31205 37139 31263 37145
rect 32122 37136 32128 37148
rect 32180 37136 32186 37188
rect 32950 37176 32956 37188
rect 32232 37148 32956 37176
rect 32232 37108 32260 37148
rect 32950 37136 32956 37148
rect 33008 37136 33014 37188
rect 33410 37136 33416 37188
rect 33468 37176 33474 37188
rect 33980 37176 34008 37207
rect 34238 37204 34244 37216
rect 34296 37204 34302 37256
rect 34698 37244 34704 37256
rect 34659 37216 34704 37244
rect 34698 37204 34704 37216
rect 34756 37204 34762 37256
rect 34885 37247 34943 37253
rect 34885 37213 34897 37247
rect 34931 37244 34943 37247
rect 35066 37244 35072 37256
rect 34931 37216 35072 37244
rect 34931 37213 34943 37216
rect 34885 37207 34943 37213
rect 35066 37204 35072 37216
rect 35124 37244 35130 37256
rect 36357 37247 36415 37253
rect 35124 37216 36308 37244
rect 35124 37204 35130 37216
rect 35342 37176 35348 37188
rect 33468 37148 35348 37176
rect 33468 37136 33474 37148
rect 35342 37136 35348 37148
rect 35400 37136 35406 37188
rect 31036 37080 32260 37108
rect 32398 37068 32404 37120
rect 32456 37108 32462 37120
rect 33870 37108 33876 37120
rect 32456 37080 33876 37108
rect 32456 37068 32462 37080
rect 33870 37068 33876 37080
rect 33928 37068 33934 37120
rect 34790 37108 34796 37120
rect 34751 37080 34796 37108
rect 34790 37068 34796 37080
rect 34848 37068 34854 37120
rect 36280 37108 36308 37216
rect 36357 37213 36369 37247
rect 36403 37213 36415 37247
rect 36357 37207 36415 37213
rect 36541 37247 36599 37253
rect 36541 37213 36553 37247
rect 36587 37244 36599 37247
rect 37185 37247 37243 37253
rect 37185 37244 37197 37247
rect 36587 37216 37197 37244
rect 36587 37213 36599 37216
rect 36541 37207 36599 37213
rect 37185 37213 37197 37216
rect 37231 37244 37243 37247
rect 37274 37244 37280 37256
rect 37231 37216 37280 37244
rect 37231 37213 37243 37216
rect 37185 37207 37243 37213
rect 36372 37176 36400 37207
rect 37274 37204 37280 37216
rect 37332 37204 37338 37256
rect 37384 37188 37412 37343
rect 37550 37340 37556 37352
rect 37608 37340 37614 37392
rect 37660 37312 37688 37420
rect 38194 37408 38200 37420
rect 38252 37408 38258 37460
rect 38654 37408 38660 37460
rect 38712 37448 38718 37460
rect 39025 37451 39083 37457
rect 39025 37448 39037 37451
rect 38712 37420 39037 37448
rect 38712 37408 38718 37420
rect 39025 37417 39037 37420
rect 39071 37417 39083 37451
rect 52822 37448 52828 37460
rect 52783 37420 52828 37448
rect 39025 37411 39083 37417
rect 52822 37408 52828 37420
rect 52880 37408 52886 37460
rect 37660 37284 37780 37312
rect 37461 37247 37519 37253
rect 37461 37213 37473 37247
rect 37507 37213 37519 37247
rect 37642 37244 37648 37256
rect 37603 37216 37648 37244
rect 37461 37207 37519 37213
rect 37366 37176 37372 37188
rect 36372 37148 37372 37176
rect 37366 37136 37372 37148
rect 37424 37136 37430 37188
rect 37476 37176 37504 37207
rect 37642 37204 37648 37216
rect 37700 37204 37706 37256
rect 37752 37244 37780 37284
rect 38105 37247 38163 37253
rect 38105 37244 38117 37247
rect 37752 37216 38117 37244
rect 38105 37213 38117 37216
rect 38151 37213 38163 37247
rect 38105 37207 38163 37213
rect 52822 37204 52828 37256
rect 52880 37244 52886 37256
rect 53377 37247 53435 37253
rect 53377 37244 53389 37247
rect 52880 37216 53389 37244
rect 52880 37204 52886 37216
rect 53377 37213 53389 37216
rect 53423 37213 53435 37247
rect 53377 37207 53435 37213
rect 38010 37176 38016 37188
rect 37476 37148 38016 37176
rect 38010 37136 38016 37148
rect 38068 37136 38074 37188
rect 38378 37176 38384 37188
rect 38120 37148 38384 37176
rect 38120 37108 38148 37148
rect 38378 37136 38384 37148
rect 38436 37136 38442 37188
rect 36280 37080 38148 37108
rect 38286 37068 38292 37120
rect 38344 37108 38350 37120
rect 38565 37111 38623 37117
rect 38565 37108 38577 37111
rect 38344 37080 38577 37108
rect 38344 37068 38350 37080
rect 38565 37077 38577 37080
rect 38611 37077 38623 37111
rect 53558 37108 53564 37120
rect 53519 37080 53564 37108
rect 38565 37071 38623 37077
rect 53558 37068 53564 37080
rect 53616 37068 53622 37120
rect 1104 37018 54372 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 54372 37018
rect 1104 36944 54372 36966
rect 17678 36904 17684 36916
rect 17512 36876 17684 36904
rect 17512 36845 17540 36876
rect 17678 36864 17684 36876
rect 17736 36864 17742 36916
rect 18138 36864 18144 36916
rect 18196 36904 18202 36916
rect 18233 36907 18291 36913
rect 18233 36904 18245 36907
rect 18196 36876 18245 36904
rect 18196 36864 18202 36876
rect 18233 36873 18245 36876
rect 18279 36873 18291 36907
rect 18233 36867 18291 36873
rect 19705 36907 19763 36913
rect 19705 36873 19717 36907
rect 19751 36904 19763 36907
rect 19978 36904 19984 36916
rect 19751 36876 19984 36904
rect 19751 36873 19763 36876
rect 19705 36867 19763 36873
rect 19978 36864 19984 36876
rect 20036 36864 20042 36916
rect 20993 36907 21051 36913
rect 20993 36873 21005 36907
rect 21039 36904 21051 36907
rect 21634 36904 21640 36916
rect 21039 36876 21640 36904
rect 21039 36873 21051 36876
rect 20993 36867 21051 36873
rect 21634 36864 21640 36876
rect 21692 36864 21698 36916
rect 21818 36864 21824 36916
rect 21876 36904 21882 36916
rect 22005 36907 22063 36913
rect 22005 36904 22017 36907
rect 21876 36876 22017 36904
rect 21876 36864 21882 36876
rect 22005 36873 22017 36876
rect 22051 36904 22063 36907
rect 22554 36904 22560 36916
rect 22051 36876 22560 36904
rect 22051 36873 22063 36876
rect 22005 36867 22063 36873
rect 22554 36864 22560 36876
rect 22612 36864 22618 36916
rect 23753 36907 23811 36913
rect 23753 36904 23765 36907
rect 23216 36876 23765 36904
rect 17497 36839 17555 36845
rect 17497 36805 17509 36839
rect 17543 36805 17555 36839
rect 18506 36836 18512 36848
rect 17497 36799 17555 36805
rect 18156 36808 18512 36836
rect 17310 36728 17316 36780
rect 17368 36768 17374 36780
rect 17405 36771 17463 36777
rect 17405 36768 17417 36771
rect 17368 36740 17417 36768
rect 17368 36728 17374 36740
rect 17405 36737 17417 36740
rect 17451 36737 17463 36771
rect 17405 36731 17463 36737
rect 17586 36728 17592 36780
rect 17644 36768 17650 36780
rect 18156 36777 18184 36808
rect 18506 36796 18512 36808
rect 18564 36796 18570 36848
rect 20257 36839 20315 36845
rect 20257 36836 20269 36839
rect 19306 36808 20269 36836
rect 17681 36771 17739 36777
rect 17681 36768 17693 36771
rect 17644 36740 17693 36768
rect 17644 36728 17650 36740
rect 17681 36737 17693 36740
rect 17727 36737 17739 36771
rect 17681 36731 17739 36737
rect 18141 36771 18199 36777
rect 18141 36737 18153 36771
rect 18187 36737 18199 36771
rect 18141 36731 18199 36737
rect 18322 36728 18328 36780
rect 18380 36768 18386 36780
rect 18417 36771 18475 36777
rect 18417 36768 18429 36771
rect 18380 36740 18429 36768
rect 18380 36728 18386 36740
rect 18417 36737 18429 36740
rect 18463 36737 18475 36771
rect 18417 36731 18475 36737
rect 19058 36728 19064 36780
rect 19116 36768 19122 36780
rect 19306 36768 19334 36808
rect 20257 36805 20269 36808
rect 20303 36836 20315 36839
rect 22370 36836 22376 36848
rect 20303 36808 22376 36836
rect 20303 36805 20315 36808
rect 20257 36799 20315 36805
rect 22370 36796 22376 36808
rect 22428 36796 22434 36848
rect 19116 36740 19334 36768
rect 20993 36771 21051 36777
rect 19116 36728 19122 36740
rect 20993 36737 21005 36771
rect 21039 36768 21051 36771
rect 21358 36768 21364 36780
rect 21039 36740 21364 36768
rect 21039 36737 21051 36740
rect 20993 36731 21051 36737
rect 21358 36728 21364 36740
rect 21416 36728 21422 36780
rect 23014 36768 23020 36780
rect 22975 36740 23020 36768
rect 23014 36728 23020 36740
rect 23072 36728 23078 36780
rect 23216 36777 23244 36876
rect 23753 36873 23765 36876
rect 23799 36904 23811 36907
rect 24854 36904 24860 36916
rect 23799 36876 24860 36904
rect 23799 36873 23811 36876
rect 23753 36867 23811 36873
rect 24854 36864 24860 36876
rect 24912 36864 24918 36916
rect 26142 36864 26148 36916
rect 26200 36904 26206 36916
rect 28077 36907 28135 36913
rect 28077 36904 28089 36907
rect 26200 36876 28089 36904
rect 26200 36864 26206 36876
rect 28077 36873 28089 36876
rect 28123 36904 28135 36907
rect 28123 36876 28994 36904
rect 28123 36873 28135 36876
rect 28077 36867 28135 36873
rect 28966 36836 28994 36876
rect 29914 36864 29920 36916
rect 29972 36904 29978 36916
rect 30929 36907 30987 36913
rect 30929 36904 30941 36907
rect 29972 36876 30941 36904
rect 29972 36864 29978 36876
rect 30929 36873 30941 36876
rect 30975 36873 30987 36907
rect 30929 36867 30987 36873
rect 33689 36907 33747 36913
rect 33689 36873 33701 36907
rect 33735 36904 33747 36907
rect 33962 36904 33968 36916
rect 33735 36876 33968 36904
rect 33735 36873 33747 36876
rect 33689 36867 33747 36873
rect 33962 36864 33968 36876
rect 34020 36864 34026 36916
rect 35066 36904 35072 36916
rect 34440 36876 35072 36904
rect 29546 36836 29552 36848
rect 23400 36808 25728 36836
rect 28966 36808 29552 36836
rect 23201 36771 23259 36777
rect 23201 36737 23213 36771
rect 23247 36737 23259 36771
rect 23201 36731 23259 36737
rect 20162 36660 20168 36712
rect 20220 36700 20226 36712
rect 20717 36703 20775 36709
rect 20717 36700 20729 36703
rect 20220 36672 20729 36700
rect 20220 36660 20226 36672
rect 20717 36669 20729 36672
rect 20763 36669 20775 36703
rect 20717 36663 20775 36669
rect 22557 36703 22615 36709
rect 22557 36669 22569 36703
rect 22603 36700 22615 36703
rect 23400 36700 23428 36808
rect 23658 36768 23664 36780
rect 23619 36740 23664 36768
rect 23658 36728 23664 36740
rect 23716 36728 23722 36780
rect 23842 36768 23848 36780
rect 23803 36740 23848 36768
rect 23842 36728 23848 36740
rect 23900 36728 23906 36780
rect 24302 36728 24308 36780
rect 24360 36768 24366 36780
rect 24489 36771 24547 36777
rect 24489 36768 24501 36771
rect 24360 36740 24501 36768
rect 24360 36728 24366 36740
rect 24489 36737 24501 36740
rect 24535 36737 24547 36771
rect 24489 36731 24547 36737
rect 24581 36771 24639 36777
rect 24581 36737 24593 36771
rect 24627 36768 24639 36771
rect 24762 36768 24768 36780
rect 24627 36740 24768 36768
rect 24627 36737 24639 36740
rect 24581 36731 24639 36737
rect 24762 36728 24768 36740
rect 24820 36728 24826 36780
rect 25700 36777 25728 36808
rect 29546 36796 29552 36808
rect 29604 36796 29610 36848
rect 30374 36836 30380 36848
rect 30335 36808 30380 36836
rect 30374 36796 30380 36808
rect 30432 36796 30438 36848
rect 31110 36836 31116 36848
rect 30852 36808 31116 36836
rect 30852 36780 30880 36808
rect 31110 36796 31116 36808
rect 31168 36796 31174 36848
rect 33778 36796 33784 36848
rect 33836 36836 33842 36848
rect 34440 36836 34468 36876
rect 35066 36864 35072 36876
rect 35124 36864 35130 36916
rect 37274 36864 37280 36916
rect 37332 36904 37338 36916
rect 37645 36907 37703 36913
rect 37645 36904 37657 36907
rect 37332 36876 37657 36904
rect 37332 36864 37338 36876
rect 37645 36873 37657 36876
rect 37691 36904 37703 36907
rect 38194 36904 38200 36916
rect 37691 36876 38200 36904
rect 37691 36873 37703 36876
rect 37645 36867 37703 36873
rect 38194 36864 38200 36876
rect 38252 36864 38258 36916
rect 33836 36808 34468 36836
rect 33836 36796 33842 36808
rect 25685 36771 25743 36777
rect 25685 36737 25697 36771
rect 25731 36737 25743 36771
rect 25685 36731 25743 36737
rect 22603 36672 23428 36700
rect 22603 36669 22615 36672
rect 22557 36663 22615 36669
rect 23750 36660 23756 36712
rect 23808 36700 23814 36712
rect 24026 36700 24032 36712
rect 23808 36672 24032 36700
rect 23808 36660 23814 36672
rect 24026 36660 24032 36672
rect 24084 36700 24090 36712
rect 24397 36703 24455 36709
rect 24397 36700 24409 36703
rect 24084 36672 24409 36700
rect 24084 36660 24090 36672
rect 24397 36669 24409 36672
rect 24443 36669 24455 36703
rect 24397 36663 24455 36669
rect 24673 36703 24731 36709
rect 24673 36669 24685 36703
rect 24719 36700 24731 36703
rect 25222 36700 25228 36712
rect 24719 36672 25228 36700
rect 24719 36669 24731 36672
rect 24673 36663 24731 36669
rect 17589 36635 17647 36641
rect 17589 36601 17601 36635
rect 17635 36632 17647 36635
rect 18414 36632 18420 36644
rect 17635 36604 18420 36632
rect 17635 36601 17647 36604
rect 17589 36595 17647 36601
rect 18414 36592 18420 36604
rect 18472 36592 18478 36644
rect 20901 36635 20959 36641
rect 20901 36601 20913 36635
rect 20947 36632 20959 36635
rect 21082 36632 21088 36644
rect 20947 36604 21088 36632
rect 20947 36601 20959 36604
rect 20901 36595 20959 36601
rect 21082 36592 21088 36604
rect 21140 36632 21146 36644
rect 21726 36632 21732 36644
rect 21140 36604 21732 36632
rect 21140 36592 21146 36604
rect 21726 36592 21732 36604
rect 21784 36592 21790 36644
rect 23109 36635 23167 36641
rect 23109 36601 23121 36635
rect 23155 36632 23167 36635
rect 23934 36632 23940 36644
rect 23155 36604 23940 36632
rect 23155 36601 23167 36604
rect 23109 36595 23167 36601
rect 23934 36592 23940 36604
rect 23992 36632 23998 36644
rect 24688 36632 24716 36663
rect 25222 36660 25228 36672
rect 25280 36660 25286 36712
rect 25406 36700 25412 36712
rect 25367 36672 25412 36700
rect 25406 36660 25412 36672
rect 25464 36660 25470 36712
rect 25700 36700 25728 36731
rect 26878 36728 26884 36780
rect 26936 36768 26942 36780
rect 26973 36771 27031 36777
rect 26973 36768 26985 36771
rect 26936 36740 26985 36768
rect 26936 36728 26942 36740
rect 26973 36737 26985 36740
rect 27019 36737 27031 36771
rect 26973 36731 27031 36737
rect 27062 36728 27068 36780
rect 27120 36768 27126 36780
rect 27430 36768 27436 36780
rect 27120 36740 27436 36768
rect 27120 36728 27126 36740
rect 27430 36728 27436 36740
rect 27488 36728 27494 36780
rect 30834 36768 30840 36780
rect 30747 36740 30840 36768
rect 30834 36728 30840 36740
rect 30892 36728 30898 36780
rect 31018 36728 31024 36780
rect 31076 36768 31082 36780
rect 32125 36771 32183 36777
rect 32125 36768 32137 36771
rect 31076 36740 32137 36768
rect 31076 36728 31082 36740
rect 32125 36737 32137 36740
rect 32171 36737 32183 36771
rect 33410 36768 33416 36780
rect 33371 36740 33416 36768
rect 32125 36731 32183 36737
rect 33410 36728 33416 36740
rect 33468 36728 33474 36780
rect 33505 36771 33563 36777
rect 33505 36737 33517 36771
rect 33551 36768 33563 36771
rect 34238 36768 34244 36780
rect 33551 36740 34244 36768
rect 33551 36737 33563 36740
rect 33505 36731 33563 36737
rect 34238 36728 34244 36740
rect 34296 36728 34302 36780
rect 34348 36777 34376 36808
rect 34790 36796 34796 36848
rect 34848 36836 34854 36848
rect 34977 36839 35035 36845
rect 34977 36836 34989 36839
rect 34848 36808 34989 36836
rect 34848 36796 34854 36808
rect 34977 36805 34989 36808
rect 35023 36805 35035 36839
rect 34977 36799 35035 36805
rect 34333 36771 34391 36777
rect 34333 36737 34345 36771
rect 34379 36737 34391 36771
rect 35158 36768 35164 36780
rect 35119 36740 35164 36768
rect 34333 36731 34391 36737
rect 35158 36728 35164 36740
rect 35216 36768 35222 36780
rect 35526 36768 35532 36780
rect 35216 36740 35532 36768
rect 35216 36728 35222 36740
rect 35526 36728 35532 36740
rect 35584 36728 35590 36780
rect 36541 36771 36599 36777
rect 36541 36737 36553 36771
rect 36587 36768 36599 36771
rect 37292 36768 37320 36864
rect 38304 36808 39528 36836
rect 36587 36740 37320 36768
rect 36587 36737 36599 36740
rect 36541 36731 36599 36737
rect 37826 36728 37832 36780
rect 37884 36768 37890 36780
rect 38304 36777 38332 36808
rect 38289 36771 38347 36777
rect 38289 36768 38301 36771
rect 37884 36740 38301 36768
rect 37884 36728 37890 36740
rect 38289 36737 38301 36740
rect 38335 36737 38347 36771
rect 38289 36731 38347 36737
rect 38657 36771 38715 36777
rect 38657 36737 38669 36771
rect 38703 36737 38715 36771
rect 38657 36731 38715 36737
rect 26510 36700 26516 36712
rect 25700 36672 26516 36700
rect 26510 36660 26516 36672
rect 26568 36660 26574 36712
rect 27249 36703 27307 36709
rect 27249 36669 27261 36703
rect 27295 36700 27307 36703
rect 27338 36700 27344 36712
rect 27295 36672 27344 36700
rect 27295 36669 27307 36672
rect 27249 36663 27307 36669
rect 27338 36660 27344 36672
rect 27396 36660 27402 36712
rect 29178 36660 29184 36712
rect 29236 36700 29242 36712
rect 31036 36700 31064 36728
rect 29236 36672 31064 36700
rect 29236 36660 29242 36672
rect 31110 36660 31116 36712
rect 31168 36700 31174 36712
rect 32769 36703 32827 36709
rect 32769 36700 32781 36703
rect 31168 36672 32781 36700
rect 31168 36660 31174 36672
rect 32769 36669 32781 36672
rect 32815 36700 32827 36703
rect 33686 36700 33692 36712
rect 32815 36672 33692 36700
rect 32815 36669 32827 36672
rect 32769 36663 32827 36669
rect 33686 36660 33692 36672
rect 33744 36660 33750 36712
rect 33962 36660 33968 36712
rect 34020 36700 34026 36712
rect 34149 36703 34207 36709
rect 34149 36700 34161 36703
rect 34020 36672 34161 36700
rect 34020 36660 34026 36672
rect 34149 36669 34161 36672
rect 34195 36700 34207 36703
rect 34698 36700 34704 36712
rect 34195 36672 34704 36700
rect 34195 36669 34207 36672
rect 34149 36663 34207 36669
rect 34698 36660 34704 36672
rect 34756 36660 34762 36712
rect 36630 36700 36636 36712
rect 36591 36672 36636 36700
rect 36630 36660 36636 36672
rect 36688 36660 36694 36712
rect 38010 36660 38016 36712
rect 38068 36700 38074 36712
rect 38672 36700 38700 36731
rect 38746 36728 38752 36780
rect 38804 36768 38810 36780
rect 39500 36777 39528 36808
rect 39301 36771 39359 36777
rect 39301 36768 39313 36771
rect 38804 36740 39313 36768
rect 38804 36728 38810 36740
rect 39301 36737 39313 36740
rect 39347 36737 39359 36771
rect 39301 36731 39359 36737
rect 39393 36771 39451 36777
rect 39393 36737 39405 36771
rect 39439 36737 39451 36771
rect 39393 36731 39451 36737
rect 39485 36771 39543 36777
rect 39485 36737 39497 36771
rect 39531 36737 39543 36771
rect 39485 36731 39543 36737
rect 39022 36700 39028 36712
rect 38068 36672 38608 36700
rect 38672 36672 39028 36700
rect 38068 36660 38074 36672
rect 23992 36604 24716 36632
rect 25501 36635 25559 36641
rect 23992 36592 23998 36604
rect 25501 36601 25513 36635
rect 25547 36632 25559 36635
rect 26234 36632 26240 36644
rect 25547 36604 26240 36632
rect 25547 36601 25559 36604
rect 25501 36595 25559 36601
rect 26234 36592 26240 36604
rect 26292 36592 26298 36644
rect 26970 36592 26976 36644
rect 27028 36632 27034 36644
rect 29089 36635 29147 36641
rect 29089 36632 29101 36635
rect 27028 36604 29101 36632
rect 27028 36592 27034 36604
rect 29089 36601 29101 36604
rect 29135 36601 29147 36635
rect 33134 36632 33140 36644
rect 29089 36595 29147 36601
rect 32869 36604 33140 36632
rect 18598 36564 18604 36576
rect 18559 36536 18604 36564
rect 18598 36524 18604 36536
rect 18656 36524 18662 36576
rect 19153 36567 19211 36573
rect 19153 36533 19165 36567
rect 19199 36564 19211 36567
rect 19242 36564 19248 36576
rect 19199 36536 19248 36564
rect 19199 36533 19211 36536
rect 19153 36527 19211 36533
rect 19242 36524 19248 36536
rect 19300 36564 19306 36576
rect 22278 36564 22284 36576
rect 19300 36536 22284 36564
rect 19300 36524 19306 36536
rect 22278 36524 22284 36536
rect 22336 36524 22342 36576
rect 24762 36524 24768 36576
rect 24820 36564 24826 36576
rect 24857 36567 24915 36573
rect 24857 36564 24869 36567
rect 24820 36536 24869 36564
rect 24820 36524 24826 36536
rect 24857 36533 24869 36536
rect 24903 36533 24915 36567
rect 25866 36564 25872 36576
rect 25827 36536 25872 36564
rect 24857 36527 24915 36533
rect 25866 36524 25872 36536
rect 25924 36524 25930 36576
rect 26326 36564 26332 36576
rect 26287 36536 26332 36564
rect 26326 36524 26332 36536
rect 26384 36524 26390 36576
rect 27154 36524 27160 36576
rect 27212 36564 27218 36576
rect 27212 36536 27257 36564
rect 27212 36524 27218 36536
rect 30650 36524 30656 36576
rect 30708 36564 30714 36576
rect 31481 36567 31539 36573
rect 31481 36564 31493 36567
rect 30708 36536 31493 36564
rect 30708 36524 30714 36536
rect 31481 36533 31493 36536
rect 31527 36564 31539 36567
rect 31754 36564 31760 36576
rect 31527 36536 31760 36564
rect 31527 36533 31539 36536
rect 31481 36527 31539 36533
rect 31754 36524 31760 36536
rect 31812 36524 31818 36576
rect 32030 36524 32036 36576
rect 32088 36564 32094 36576
rect 32869 36564 32897 36604
rect 33134 36592 33140 36604
rect 33192 36632 33198 36644
rect 33502 36632 33508 36644
rect 33192 36604 33508 36632
rect 33192 36592 33198 36604
rect 33502 36592 33508 36604
rect 33560 36592 33566 36644
rect 33778 36592 33784 36644
rect 33836 36632 33842 36644
rect 36173 36635 36231 36641
rect 36173 36632 36185 36635
rect 33836 36604 36185 36632
rect 33836 36592 33842 36604
rect 36173 36601 36185 36604
rect 36219 36601 36231 36635
rect 38580 36632 38608 36672
rect 39022 36660 39028 36672
rect 39080 36700 39086 36712
rect 39408 36700 39436 36731
rect 39080 36672 39436 36700
rect 39080 36660 39086 36672
rect 39669 36635 39727 36641
rect 39669 36632 39681 36635
rect 38580 36604 39681 36632
rect 36173 36595 36231 36601
rect 39669 36601 39681 36604
rect 39715 36601 39727 36635
rect 39669 36595 39727 36601
rect 32088 36536 32897 36564
rect 32088 36524 32094 36536
rect 33318 36524 33324 36576
rect 33376 36564 33382 36576
rect 33962 36564 33968 36576
rect 33376 36536 33968 36564
rect 33376 36524 33382 36536
rect 33962 36524 33968 36536
rect 34020 36524 34026 36576
rect 34146 36524 34152 36576
rect 34204 36564 34210 36576
rect 34517 36567 34575 36573
rect 34517 36564 34529 36567
rect 34204 36536 34529 36564
rect 34204 36524 34210 36536
rect 34517 36533 34529 36536
rect 34563 36564 34575 36567
rect 35158 36564 35164 36576
rect 34563 36536 35164 36564
rect 34563 36533 34575 36536
rect 34517 36527 34575 36533
rect 35158 36524 35164 36536
rect 35216 36524 35222 36576
rect 35342 36564 35348 36576
rect 35303 36536 35348 36564
rect 35342 36524 35348 36536
rect 35400 36524 35406 36576
rect 1104 36474 54372 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 54372 36474
rect 1104 36400 54372 36422
rect 20625 36363 20683 36369
rect 20625 36329 20637 36363
rect 20671 36360 20683 36363
rect 21082 36360 21088 36372
rect 20671 36332 21088 36360
rect 20671 36329 20683 36332
rect 20625 36323 20683 36329
rect 21082 36320 21088 36332
rect 21140 36320 21146 36372
rect 23014 36320 23020 36372
rect 23072 36360 23078 36372
rect 23477 36363 23535 36369
rect 23477 36360 23489 36363
rect 23072 36332 23489 36360
rect 23072 36320 23078 36332
rect 23477 36329 23489 36332
rect 23523 36329 23535 36363
rect 23477 36323 23535 36329
rect 24765 36363 24823 36369
rect 24765 36329 24777 36363
rect 24811 36360 24823 36363
rect 25406 36360 25412 36372
rect 24811 36332 25412 36360
rect 24811 36329 24823 36332
rect 24765 36323 24823 36329
rect 25406 36320 25412 36332
rect 25464 36320 25470 36372
rect 28534 36320 28540 36372
rect 28592 36360 28598 36372
rect 30561 36363 30619 36369
rect 30561 36360 30573 36363
rect 28592 36332 30573 36360
rect 28592 36320 28598 36332
rect 30561 36329 30573 36332
rect 30607 36329 30619 36363
rect 33686 36360 33692 36372
rect 30561 36323 30619 36329
rect 31726 36332 33692 36360
rect 17586 36252 17592 36304
rect 17644 36292 17650 36304
rect 17865 36295 17923 36301
rect 17865 36292 17877 36295
rect 17644 36264 17877 36292
rect 17644 36252 17650 36264
rect 17865 36261 17877 36264
rect 17911 36261 17923 36295
rect 17865 36255 17923 36261
rect 17954 36252 17960 36304
rect 18012 36292 18018 36304
rect 18230 36292 18236 36304
rect 18012 36264 18236 36292
rect 18012 36252 18018 36264
rect 18230 36252 18236 36264
rect 18288 36252 18294 36304
rect 21910 36292 21916 36304
rect 20548 36264 21916 36292
rect 18138 36184 18144 36236
rect 18196 36224 18202 36236
rect 18196 36196 19564 36224
rect 18196 36184 18202 36196
rect 17310 36116 17316 36168
rect 17368 36156 17374 36168
rect 17773 36159 17831 36165
rect 17773 36156 17785 36159
rect 17368 36128 17785 36156
rect 17368 36116 17374 36128
rect 17773 36125 17785 36128
rect 17819 36125 17831 36159
rect 17773 36119 17831 36125
rect 18046 36116 18052 36168
rect 18104 36156 18110 36168
rect 18230 36156 18236 36168
rect 18104 36128 18149 36156
rect 18191 36128 18236 36156
rect 18104 36116 18110 36128
rect 18230 36116 18236 36128
rect 18288 36116 18294 36168
rect 18506 36116 18512 36168
rect 18564 36156 18570 36168
rect 19536 36165 19564 36196
rect 20162 36184 20168 36236
rect 20220 36224 20226 36236
rect 20548 36233 20576 36264
rect 21910 36252 21916 36264
rect 21968 36292 21974 36304
rect 29638 36292 29644 36304
rect 21968 36264 22324 36292
rect 29599 36264 29644 36292
rect 21968 36252 21974 36264
rect 20533 36227 20591 36233
rect 20533 36224 20545 36227
rect 20220 36196 20545 36224
rect 20220 36184 20226 36196
rect 20533 36193 20545 36196
rect 20579 36193 20591 36227
rect 21634 36224 21640 36236
rect 21547 36196 21640 36224
rect 20533 36187 20591 36193
rect 21634 36184 21640 36196
rect 21692 36224 21698 36236
rect 22189 36227 22247 36233
rect 22189 36224 22201 36227
rect 21692 36196 22201 36224
rect 21692 36184 21698 36196
rect 22189 36193 22201 36196
rect 22235 36193 22247 36227
rect 22189 36187 22247 36193
rect 19429 36159 19487 36165
rect 19429 36156 19441 36159
rect 18564 36128 19441 36156
rect 18564 36116 18570 36128
rect 19429 36125 19441 36128
rect 19475 36125 19487 36159
rect 19429 36119 19487 36125
rect 19521 36159 19579 36165
rect 19521 36125 19533 36159
rect 19567 36125 19579 36159
rect 19521 36119 19579 36125
rect 20441 36159 20499 36165
rect 20441 36125 20453 36159
rect 20487 36125 20499 36159
rect 21450 36156 21456 36168
rect 21411 36128 21456 36156
rect 20441 36119 20499 36125
rect 1854 36088 1860 36100
rect 1815 36060 1860 36088
rect 1854 36048 1860 36060
rect 1912 36048 1918 36100
rect 16390 36048 16396 36100
rect 16448 36088 16454 36100
rect 17129 36091 17187 36097
rect 17129 36088 17141 36091
rect 16448 36060 17141 36088
rect 16448 36048 16454 36060
rect 17129 36057 17141 36060
rect 17175 36088 17187 36091
rect 18690 36088 18696 36100
rect 17175 36060 18696 36088
rect 17175 36057 17187 36060
rect 17129 36051 17187 36057
rect 18690 36048 18696 36060
rect 18748 36048 18754 36100
rect 19245 36091 19303 36097
rect 19245 36057 19257 36091
rect 19291 36057 19303 36091
rect 20456 36088 20484 36119
rect 21450 36116 21456 36128
rect 21508 36116 21514 36168
rect 21726 36116 21732 36168
rect 21784 36156 21790 36168
rect 22296 36165 22324 36264
rect 29638 36252 29644 36264
rect 29696 36292 29702 36304
rect 30098 36292 30104 36304
rect 29696 36264 30104 36292
rect 29696 36252 29702 36264
rect 30098 36252 30104 36264
rect 30156 36252 30162 36304
rect 31726 36292 31754 36332
rect 33686 36320 33692 36332
rect 33744 36360 33750 36372
rect 33744 36332 34560 36360
rect 33744 36320 33750 36332
rect 33042 36292 33048 36304
rect 30484 36264 31754 36292
rect 32692 36264 33048 36292
rect 25866 36184 25872 36236
rect 25924 36224 25930 36236
rect 26605 36227 26663 36233
rect 26605 36224 26617 36227
rect 25924 36196 26617 36224
rect 25924 36184 25930 36196
rect 26605 36193 26617 36196
rect 26651 36193 26663 36227
rect 26605 36187 26663 36193
rect 26881 36227 26939 36233
rect 26881 36193 26893 36227
rect 26927 36224 26939 36227
rect 26970 36224 26976 36236
rect 26927 36196 26976 36224
rect 26927 36193 26939 36196
rect 26881 36187 26939 36193
rect 26970 36184 26976 36196
rect 27028 36184 27034 36236
rect 28718 36224 28724 36236
rect 28679 36196 28724 36224
rect 28718 36184 28724 36196
rect 28776 36184 28782 36236
rect 30484 36224 30512 36264
rect 32692 36233 32720 36264
rect 33042 36252 33048 36264
rect 33100 36252 33106 36304
rect 33778 36252 33784 36304
rect 33836 36252 33842 36304
rect 34532 36292 34560 36332
rect 34606 36320 34612 36372
rect 34664 36360 34670 36372
rect 35529 36363 35587 36369
rect 35529 36360 35541 36363
rect 34664 36332 35541 36360
rect 34664 36320 34670 36332
rect 35529 36329 35541 36332
rect 35575 36329 35587 36363
rect 38746 36360 38752 36372
rect 38707 36332 38752 36360
rect 35529 36323 35587 36329
rect 38746 36320 38752 36332
rect 38804 36320 38810 36372
rect 34882 36292 34888 36304
rect 34532 36264 34888 36292
rect 34882 36252 34888 36264
rect 34940 36252 34946 36304
rect 34977 36295 35035 36301
rect 34977 36261 34989 36295
rect 35023 36261 35035 36295
rect 39022 36292 39028 36304
rect 34977 36255 35035 36261
rect 37844 36264 39028 36292
rect 31021 36227 31079 36233
rect 31021 36224 31033 36227
rect 28828 36196 30512 36224
rect 30576 36196 31033 36224
rect 22097 36159 22155 36165
rect 22097 36156 22109 36159
rect 21784 36128 22109 36156
rect 21784 36116 21790 36128
rect 22097 36125 22109 36128
rect 22143 36125 22155 36159
rect 22097 36119 22155 36125
rect 22281 36159 22339 36165
rect 22281 36125 22293 36159
rect 22327 36125 22339 36159
rect 24578 36156 24584 36168
rect 24539 36128 24584 36156
rect 22281 36119 22339 36125
rect 24578 36116 24584 36128
rect 24636 36116 24642 36168
rect 24762 36156 24768 36168
rect 24723 36128 24768 36156
rect 24762 36116 24768 36128
rect 24820 36116 24826 36168
rect 26326 36156 26332 36168
rect 25240 36128 26332 36156
rect 21358 36088 21364 36100
rect 20456 36060 21364 36088
rect 19245 36051 19303 36057
rect 1949 36023 2007 36029
rect 1949 35989 1961 36023
rect 1995 36020 2007 36023
rect 15470 36020 15476 36032
rect 1995 35992 15476 36020
rect 1995 35989 2007 35992
rect 1949 35983 2007 35989
rect 15470 35980 15476 35992
rect 15528 35980 15534 36032
rect 16577 36023 16635 36029
rect 16577 35989 16589 36023
rect 16623 36020 16635 36023
rect 16942 36020 16948 36032
rect 16623 35992 16948 36020
rect 16623 35989 16635 35992
rect 16577 35983 16635 35989
rect 16942 35980 16948 35992
rect 17000 35980 17006 36032
rect 17586 36020 17592 36032
rect 17547 35992 17592 36020
rect 17586 35980 17592 35992
rect 17644 35980 17650 36032
rect 17954 35980 17960 36032
rect 18012 36020 18018 36032
rect 19260 36020 19288 36051
rect 21358 36048 21364 36060
rect 21416 36048 21422 36100
rect 23658 36088 23664 36100
rect 23619 36060 23664 36088
rect 23658 36048 23664 36060
rect 23716 36048 23722 36100
rect 23842 36088 23848 36100
rect 23803 36060 23848 36088
rect 23842 36048 23848 36060
rect 23900 36088 23906 36100
rect 25240 36097 25268 36128
rect 26326 36116 26332 36128
rect 26384 36156 26390 36168
rect 26384 36128 26924 36156
rect 26384 36116 26390 36128
rect 26896 36100 26924 36128
rect 27706 36116 27712 36168
rect 27764 36156 27770 36168
rect 28828 36156 28856 36196
rect 28994 36156 29000 36168
rect 27764 36128 28856 36156
rect 28955 36128 29000 36156
rect 27764 36116 27770 36128
rect 28994 36116 29000 36128
rect 29052 36116 29058 36168
rect 29546 36116 29552 36168
rect 29604 36156 29610 36168
rect 29641 36159 29699 36165
rect 29641 36156 29653 36159
rect 29604 36128 29653 36156
rect 29604 36116 29610 36128
rect 29641 36125 29653 36128
rect 29687 36156 29699 36159
rect 30466 36156 30472 36168
rect 29687 36128 30472 36156
rect 29687 36125 29699 36128
rect 29641 36119 29699 36125
rect 30466 36116 30472 36128
rect 30524 36116 30530 36168
rect 25225 36091 25283 36097
rect 25225 36088 25237 36091
rect 23900 36060 25237 36088
rect 23900 36048 23906 36060
rect 25225 36057 25237 36060
rect 25271 36057 25283 36091
rect 25225 36051 25283 36057
rect 26878 36048 26884 36100
rect 26936 36048 26942 36100
rect 30190 36048 30196 36100
rect 30248 36088 30254 36100
rect 30576 36088 30604 36196
rect 31021 36193 31033 36196
rect 31067 36193 31079 36227
rect 31021 36187 31079 36193
rect 32677 36227 32735 36233
rect 32677 36193 32689 36227
rect 32723 36193 32735 36227
rect 32677 36187 32735 36193
rect 32953 36227 33011 36233
rect 32953 36193 32965 36227
rect 32999 36224 33011 36227
rect 32999 36196 33732 36224
rect 32999 36193 33011 36196
rect 32953 36187 33011 36193
rect 30742 36156 30748 36168
rect 30703 36128 30748 36156
rect 30742 36116 30748 36128
rect 30800 36116 30806 36168
rect 30837 36159 30895 36165
rect 30837 36125 30849 36159
rect 30883 36125 30895 36159
rect 31110 36156 31116 36168
rect 31071 36128 31116 36156
rect 30837 36119 30895 36125
rect 30248 36060 30604 36088
rect 30248 36048 30254 36060
rect 30650 36048 30656 36100
rect 30708 36088 30714 36100
rect 30852 36088 30880 36119
rect 31110 36116 31116 36128
rect 31168 36116 31174 36168
rect 32585 36159 32643 36165
rect 32585 36125 32597 36159
rect 32631 36156 32643 36159
rect 32858 36156 32864 36168
rect 32631 36128 32864 36156
rect 32631 36125 32643 36128
rect 32585 36119 32643 36125
rect 32858 36116 32864 36128
rect 32916 36116 32922 36168
rect 33502 36116 33508 36168
rect 33560 36154 33566 36168
rect 33597 36159 33655 36165
rect 33597 36154 33609 36159
rect 33560 36126 33609 36154
rect 33560 36116 33566 36126
rect 33597 36125 33609 36126
rect 33643 36125 33655 36159
rect 33597 36119 33655 36125
rect 30708 36060 30880 36088
rect 30708 36048 30714 36060
rect 31938 36048 31944 36100
rect 31996 36088 32002 36100
rect 33704 36088 33732 36196
rect 33796 36165 33824 36252
rect 33870 36184 33876 36236
rect 33928 36224 33934 36236
rect 34992 36224 35020 36255
rect 33928 36196 33973 36224
rect 34256 36196 35020 36224
rect 33928 36184 33934 36196
rect 33781 36159 33839 36165
rect 33781 36125 33793 36159
rect 33827 36125 33839 36159
rect 33781 36119 33839 36125
rect 33965 36157 34023 36163
rect 33965 36123 33977 36157
rect 34011 36123 34023 36157
rect 33965 36117 34023 36123
rect 34149 36161 34207 36167
rect 34149 36127 34161 36161
rect 34195 36158 34207 36161
rect 34256 36158 34284 36196
rect 35158 36184 35164 36236
rect 35216 36224 35222 36236
rect 35713 36227 35771 36233
rect 35713 36224 35725 36227
rect 35216 36196 35725 36224
rect 35216 36184 35222 36196
rect 35713 36193 35725 36196
rect 35759 36193 35771 36227
rect 35713 36187 35771 36193
rect 34195 36130 34284 36158
rect 34195 36127 34207 36130
rect 34149 36121 34207 36127
rect 33980 36088 34008 36117
rect 34330 36116 34336 36168
rect 34388 36156 34394 36168
rect 34701 36159 34759 36165
rect 34701 36156 34713 36159
rect 34388 36128 34713 36156
rect 34388 36116 34394 36128
rect 34701 36125 34713 36128
rect 34747 36125 34759 36159
rect 34701 36119 34759 36125
rect 35437 36159 35495 36165
rect 35437 36125 35449 36159
rect 35483 36156 35495 36159
rect 35526 36156 35532 36168
rect 35483 36128 35532 36156
rect 35483 36125 35495 36128
rect 35437 36119 35495 36125
rect 35526 36116 35532 36128
rect 35584 36116 35590 36168
rect 35728 36156 35756 36187
rect 35802 36184 35808 36236
rect 35860 36224 35866 36236
rect 37844 36233 37872 36264
rect 39022 36252 39028 36264
rect 39080 36252 39086 36304
rect 36633 36227 36691 36233
rect 36633 36224 36645 36227
rect 35860 36196 36645 36224
rect 35860 36184 35866 36196
rect 36633 36193 36645 36196
rect 36679 36193 36691 36227
rect 36633 36187 36691 36193
rect 37093 36227 37151 36233
rect 37093 36193 37105 36227
rect 37139 36224 37151 36227
rect 37645 36227 37703 36233
rect 37645 36224 37657 36227
rect 37139 36196 37657 36224
rect 37139 36193 37151 36196
rect 37093 36187 37151 36193
rect 37645 36193 37657 36196
rect 37691 36193 37703 36227
rect 37645 36187 37703 36193
rect 37829 36227 37887 36233
rect 37829 36193 37841 36227
rect 37875 36193 37887 36227
rect 38286 36224 38292 36236
rect 38247 36196 38292 36224
rect 37829 36187 37887 36193
rect 38286 36184 38292 36196
rect 38344 36184 38350 36236
rect 36170 36156 36176 36168
rect 35728 36128 36176 36156
rect 36170 36116 36176 36128
rect 36228 36116 36234 36168
rect 37001 36159 37059 36165
rect 37001 36125 37013 36159
rect 37047 36156 37059 36159
rect 37366 36156 37372 36168
rect 37047 36128 37372 36156
rect 37047 36125 37059 36128
rect 37001 36119 37059 36125
rect 37366 36116 37372 36128
rect 37424 36116 37430 36168
rect 37921 36159 37979 36165
rect 37921 36125 37933 36159
rect 37967 36125 37979 36159
rect 38746 36156 38752 36168
rect 38707 36128 38752 36156
rect 37921 36119 37979 36125
rect 31996 36060 33548 36088
rect 33704 36060 34008 36088
rect 31996 36048 32002 36060
rect 18012 35992 19288 36020
rect 19521 36023 19579 36029
rect 18012 35980 18018 35992
rect 19521 35989 19533 36023
rect 19567 36020 19579 36023
rect 19978 36020 19984 36032
rect 19567 35992 19984 36020
rect 19567 35989 19579 35992
rect 19521 35983 19579 35989
rect 19978 35980 19984 35992
rect 20036 35980 20042 36032
rect 20809 36023 20867 36029
rect 20809 35989 20821 36023
rect 20855 36020 20867 36023
rect 20898 36020 20904 36032
rect 20855 35992 20904 36020
rect 20855 35989 20867 35992
rect 20809 35983 20867 35989
rect 20898 35980 20904 35992
rect 20956 35980 20962 36032
rect 21266 36020 21272 36032
rect 21227 35992 21272 36020
rect 21266 35980 21272 35992
rect 21324 35980 21330 36032
rect 23017 36023 23075 36029
rect 23017 35989 23029 36023
rect 23063 36020 23075 36023
rect 24026 36020 24032 36032
rect 23063 35992 24032 36020
rect 23063 35989 23075 35992
rect 23017 35983 23075 35989
rect 24026 35980 24032 35992
rect 24084 35980 24090 36032
rect 27433 36023 27491 36029
rect 27433 35989 27445 36023
rect 27479 36020 27491 36023
rect 29178 36020 29184 36032
rect 27479 35992 29184 36020
rect 27479 35989 27491 35992
rect 27433 35983 27491 35989
rect 29178 35980 29184 35992
rect 29236 35980 29242 36032
rect 31570 36020 31576 36032
rect 31531 35992 31576 36020
rect 31570 35980 31576 35992
rect 31628 35980 31634 36032
rect 31846 35980 31852 36032
rect 31904 36020 31910 36032
rect 33413 36023 33471 36029
rect 33413 36020 33425 36023
rect 31904 35992 33425 36020
rect 31904 35980 31910 35992
rect 33413 35989 33425 35992
rect 33459 35989 33471 36023
rect 33520 36020 33548 36060
rect 34882 36048 34888 36100
rect 34940 36088 34946 36100
rect 34977 36091 35035 36097
rect 34977 36088 34989 36091
rect 34940 36060 34989 36088
rect 34940 36048 34946 36060
rect 34977 36057 34989 36060
rect 35023 36088 35035 36091
rect 35023 36060 35848 36088
rect 35023 36057 35035 36060
rect 34977 36051 35035 36057
rect 34422 36020 34428 36032
rect 33520 35992 34428 36020
rect 33413 35983 33471 35989
rect 34422 35980 34428 35992
rect 34480 35980 34486 36032
rect 34793 36023 34851 36029
rect 34793 35989 34805 36023
rect 34839 36020 34851 36023
rect 35713 36023 35771 36029
rect 35713 36020 35725 36023
rect 34839 35992 35725 36020
rect 34839 35989 34851 35992
rect 34793 35983 34851 35989
rect 35713 35989 35725 35992
rect 35759 35989 35771 36023
rect 35820 36020 35848 36060
rect 35986 36048 35992 36100
rect 36044 36088 36050 36100
rect 37642 36088 37648 36100
rect 36044 36060 37648 36088
rect 36044 36048 36050 36060
rect 37642 36048 37648 36060
rect 37700 36048 37706 36100
rect 37826 36048 37832 36100
rect 37884 36088 37890 36100
rect 37936 36088 37964 36119
rect 38746 36116 38752 36128
rect 38804 36116 38810 36168
rect 38933 36159 38991 36165
rect 38933 36125 38945 36159
rect 38979 36125 38991 36159
rect 38933 36119 38991 36125
rect 37884 36060 37964 36088
rect 38948 36088 38976 36119
rect 39758 36088 39764 36100
rect 38948 36060 39764 36088
rect 37884 36048 37890 36060
rect 39758 36048 39764 36060
rect 39816 36088 39822 36100
rect 39816 36060 40540 36088
rect 39816 36048 39822 36060
rect 40512 36029 40540 36060
rect 39853 36023 39911 36029
rect 39853 36020 39865 36023
rect 35820 35992 39865 36020
rect 35713 35983 35771 35989
rect 39853 35989 39865 35992
rect 39899 35989 39911 36023
rect 39853 35983 39911 35989
rect 40497 36023 40555 36029
rect 40497 35989 40509 36023
rect 40543 36020 40555 36023
rect 52362 36020 52368 36032
rect 40543 35992 52368 36020
rect 40543 35989 40555 35992
rect 40497 35983 40555 35989
rect 52362 35980 52368 35992
rect 52420 35980 52426 36032
rect 1104 35930 54372 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 54372 35930
rect 1104 35856 54372 35878
rect 1673 35819 1731 35825
rect 1673 35785 1685 35819
rect 1719 35816 1731 35819
rect 1854 35816 1860 35828
rect 1719 35788 1860 35816
rect 1719 35785 1731 35788
rect 1673 35779 1731 35785
rect 1854 35776 1860 35788
rect 1912 35776 1918 35828
rect 18046 35816 18052 35828
rect 18007 35788 18052 35816
rect 18046 35776 18052 35788
rect 18104 35776 18110 35828
rect 18598 35776 18604 35828
rect 18656 35816 18662 35828
rect 19242 35816 19248 35828
rect 18656 35788 19248 35816
rect 18656 35776 18662 35788
rect 19242 35776 19248 35788
rect 19300 35776 19306 35828
rect 19978 35816 19984 35828
rect 20036 35825 20042 35828
rect 20036 35819 20055 35825
rect 19352 35788 19984 35816
rect 17497 35751 17555 35757
rect 17497 35717 17509 35751
rect 17543 35748 17555 35751
rect 17954 35748 17960 35760
rect 17543 35720 17960 35748
rect 17543 35717 17555 35720
rect 17497 35711 17555 35717
rect 17954 35708 17960 35720
rect 18012 35708 18018 35760
rect 17405 35683 17463 35689
rect 17405 35649 17417 35683
rect 17451 35649 17463 35683
rect 17405 35643 17463 35649
rect 17589 35683 17647 35689
rect 17589 35649 17601 35683
rect 17635 35680 17647 35683
rect 18509 35683 18567 35689
rect 18509 35680 18521 35683
rect 17635 35652 18521 35680
rect 17635 35649 17647 35652
rect 17589 35643 17647 35649
rect 18509 35649 18521 35652
rect 18555 35680 18567 35683
rect 18874 35680 18880 35692
rect 18555 35652 18880 35680
rect 18555 35649 18567 35652
rect 18509 35643 18567 35649
rect 17420 35612 17448 35643
rect 18874 35640 18880 35652
rect 18932 35640 18938 35692
rect 19352 35689 19380 35788
rect 19978 35776 19984 35788
rect 20043 35785 20055 35819
rect 20162 35816 20168 35828
rect 20123 35788 20168 35816
rect 20036 35779 20055 35785
rect 20036 35776 20042 35779
rect 20162 35776 20168 35788
rect 20220 35776 20226 35828
rect 20622 35776 20628 35828
rect 20680 35816 20686 35828
rect 25225 35819 25283 35825
rect 20680 35788 21128 35816
rect 20680 35776 20686 35788
rect 19797 35751 19855 35757
rect 19797 35748 19809 35751
rect 19720 35720 19809 35748
rect 19061 35683 19119 35689
rect 19061 35649 19073 35683
rect 19107 35649 19119 35683
rect 19061 35643 19119 35649
rect 19337 35683 19395 35689
rect 19337 35649 19349 35683
rect 19383 35649 19395 35683
rect 19337 35643 19395 35649
rect 18230 35612 18236 35624
rect 17420 35584 18236 35612
rect 18230 35572 18236 35584
rect 18288 35572 18294 35624
rect 18690 35572 18696 35624
rect 18748 35612 18754 35624
rect 19076 35612 19104 35643
rect 19150 35612 19156 35624
rect 18748 35584 19156 35612
rect 18748 35572 18754 35584
rect 19150 35572 19156 35584
rect 19208 35612 19214 35624
rect 19720 35612 19748 35720
rect 19797 35717 19809 35720
rect 19843 35748 19855 35751
rect 19843 35720 21036 35748
rect 19843 35717 19855 35720
rect 19797 35711 19855 35717
rect 20622 35680 20628 35692
rect 20583 35652 20628 35680
rect 20622 35640 20628 35652
rect 20680 35640 20686 35692
rect 20806 35680 20812 35692
rect 20767 35652 20812 35680
rect 20806 35640 20812 35652
rect 20864 35640 20870 35692
rect 20898 35612 20904 35624
rect 19208 35584 19748 35612
rect 20859 35584 20904 35612
rect 19208 35572 19214 35584
rect 20898 35572 20904 35584
rect 20956 35572 20962 35624
rect 21008 35612 21036 35720
rect 21100 35689 21128 35788
rect 25225 35785 25237 35819
rect 25271 35816 25283 35819
rect 25314 35816 25320 35828
rect 25271 35788 25320 35816
rect 25271 35785 25283 35788
rect 25225 35779 25283 35785
rect 25314 35776 25320 35788
rect 25372 35776 25378 35828
rect 26234 35776 26240 35828
rect 26292 35816 26298 35828
rect 26329 35819 26387 35825
rect 26329 35816 26341 35819
rect 26292 35788 26341 35816
rect 26292 35776 26298 35788
rect 26329 35785 26341 35788
rect 26375 35785 26387 35819
rect 26329 35779 26387 35785
rect 31754 35776 31760 35828
rect 31812 35816 31818 35828
rect 34330 35816 34336 35828
rect 31812 35788 32536 35816
rect 34291 35788 34336 35816
rect 31812 35776 31818 35788
rect 25777 35751 25835 35757
rect 25777 35748 25789 35751
rect 23308 35720 25789 35748
rect 21085 35683 21143 35689
rect 21085 35649 21097 35683
rect 21131 35649 21143 35683
rect 21085 35643 21143 35649
rect 21634 35640 21640 35692
rect 21692 35680 21698 35692
rect 22005 35683 22063 35689
rect 22005 35680 22017 35683
rect 21692 35652 22017 35680
rect 21692 35640 21698 35652
rect 22005 35649 22017 35652
rect 22051 35649 22063 35683
rect 22005 35643 22063 35649
rect 22738 35640 22744 35692
rect 22796 35680 22802 35692
rect 23308 35680 23336 35720
rect 25777 35717 25789 35720
rect 25823 35748 25835 35751
rect 27982 35748 27988 35760
rect 25823 35720 27988 35748
rect 25823 35717 25835 35720
rect 25777 35711 25835 35717
rect 27982 35708 27988 35720
rect 28040 35708 28046 35760
rect 30374 35748 30380 35760
rect 30335 35720 30380 35748
rect 30374 35708 30380 35720
rect 30432 35708 30438 35760
rect 30742 35708 30748 35760
rect 30800 35748 30806 35760
rect 30800 35720 32260 35748
rect 30800 35708 30806 35720
rect 24118 35680 24124 35692
rect 22796 35652 23336 35680
rect 24079 35652 24124 35680
rect 22796 35640 22802 35652
rect 24118 35640 24124 35652
rect 24176 35640 24182 35692
rect 24210 35640 24216 35692
rect 24268 35680 24274 35692
rect 24305 35683 24363 35689
rect 24305 35680 24317 35683
rect 24268 35652 24317 35680
rect 24268 35640 24274 35652
rect 24305 35649 24317 35652
rect 24351 35649 24363 35683
rect 24305 35643 24363 35649
rect 24397 35683 24455 35689
rect 24397 35649 24409 35683
rect 24443 35680 24455 35683
rect 24762 35680 24768 35692
rect 24443 35652 24768 35680
rect 24443 35649 24455 35652
rect 24397 35643 24455 35649
rect 24762 35640 24768 35652
rect 24820 35640 24826 35692
rect 26053 35683 26111 35689
rect 26053 35649 26065 35683
rect 26099 35680 26111 35683
rect 27062 35680 27068 35692
rect 26099 35652 27068 35680
rect 26099 35649 26111 35652
rect 26053 35643 26111 35649
rect 27062 35640 27068 35652
rect 27120 35640 27126 35692
rect 27157 35683 27215 35689
rect 27157 35649 27169 35683
rect 27203 35680 27215 35683
rect 27430 35680 27436 35692
rect 27203 35652 27436 35680
rect 27203 35649 27215 35652
rect 27157 35643 27215 35649
rect 27430 35640 27436 35652
rect 27488 35640 27494 35692
rect 32030 35640 32036 35692
rect 32088 35680 32094 35692
rect 32125 35683 32183 35689
rect 32125 35680 32137 35683
rect 32088 35652 32137 35680
rect 32088 35640 32094 35652
rect 32125 35649 32137 35652
rect 32171 35649 32183 35683
rect 32232 35680 32260 35720
rect 32508 35689 32536 35788
rect 34330 35776 34336 35788
rect 34388 35776 34394 35828
rect 34698 35776 34704 35828
rect 34756 35816 34762 35828
rect 34793 35819 34851 35825
rect 34793 35816 34805 35819
rect 34756 35788 34805 35816
rect 34756 35776 34762 35788
rect 34793 35785 34805 35788
rect 34839 35785 34851 35819
rect 34793 35779 34851 35785
rect 36541 35819 36599 35825
rect 36541 35785 36553 35819
rect 36587 35816 36599 35819
rect 36630 35816 36636 35828
rect 36587 35788 36636 35816
rect 36587 35785 36599 35788
rect 36541 35779 36599 35785
rect 36630 35776 36636 35788
rect 36688 35776 36694 35828
rect 37277 35819 37335 35825
rect 37277 35816 37289 35819
rect 36740 35788 37289 35816
rect 35342 35748 35348 35760
rect 34992 35720 35348 35748
rect 32304 35683 32362 35689
rect 32304 35680 32316 35683
rect 32232 35652 32316 35680
rect 32125 35643 32183 35649
rect 32304 35649 32316 35652
rect 32350 35649 32362 35683
rect 32304 35643 32362 35649
rect 32401 35683 32459 35689
rect 32401 35649 32413 35683
rect 32447 35649 32459 35683
rect 32401 35643 32459 35649
rect 32493 35683 32551 35689
rect 32493 35649 32505 35683
rect 32539 35649 32551 35683
rect 32493 35643 32551 35649
rect 33873 35683 33931 35689
rect 33873 35649 33885 35683
rect 33919 35680 33931 35683
rect 33962 35680 33968 35692
rect 33919 35652 33968 35680
rect 33919 35649 33931 35652
rect 33873 35643 33931 35649
rect 21008 35584 21404 35612
rect 19061 35547 19119 35553
rect 19061 35513 19073 35547
rect 19107 35544 19119 35547
rect 20993 35547 21051 35553
rect 19107 35516 20944 35544
rect 19107 35513 19119 35516
rect 19061 35507 19119 35513
rect 20916 35488 20944 35516
rect 20993 35513 21005 35547
rect 21039 35544 21051 35547
rect 21082 35544 21088 35556
rect 21039 35516 21088 35544
rect 21039 35513 21051 35516
rect 20993 35507 21051 35513
rect 21082 35504 21088 35516
rect 21140 35504 21146 35556
rect 21376 35544 21404 35584
rect 21450 35572 21456 35624
rect 21508 35612 21514 35624
rect 21913 35615 21971 35621
rect 21913 35612 21925 35615
rect 21508 35584 21925 35612
rect 21508 35572 21514 35584
rect 21913 35581 21925 35584
rect 21959 35581 21971 35615
rect 21913 35575 21971 35581
rect 22373 35615 22431 35621
rect 22373 35581 22385 35615
rect 22419 35612 22431 35615
rect 25685 35615 25743 35621
rect 25685 35612 25697 35615
rect 22419 35584 25697 35612
rect 22419 35581 22431 35584
rect 22373 35575 22431 35581
rect 25685 35581 25697 35584
rect 25731 35581 25743 35615
rect 25685 35575 25743 35581
rect 26176 35615 26234 35621
rect 26176 35581 26188 35615
rect 26222 35612 26234 35615
rect 26222 35584 26464 35612
rect 26222 35581 26234 35584
rect 26176 35575 26234 35581
rect 22925 35547 22983 35553
rect 21376 35516 22876 35544
rect 15930 35436 15936 35488
rect 15988 35476 15994 35488
rect 16025 35479 16083 35485
rect 16025 35476 16037 35479
rect 15988 35448 16037 35476
rect 15988 35436 15994 35448
rect 16025 35445 16037 35448
rect 16071 35476 16083 35479
rect 16390 35476 16396 35488
rect 16071 35448 16396 35476
rect 16071 35445 16083 35448
rect 16025 35439 16083 35445
rect 16390 35436 16396 35448
rect 16448 35436 16454 35488
rect 16850 35476 16856 35488
rect 16811 35448 16856 35476
rect 16850 35436 16856 35448
rect 16908 35436 16914 35488
rect 18138 35436 18144 35488
rect 18196 35476 18202 35488
rect 18233 35479 18291 35485
rect 18233 35476 18245 35479
rect 18196 35448 18245 35476
rect 18196 35436 18202 35448
rect 18233 35445 18245 35448
rect 18279 35445 18291 35479
rect 18233 35439 18291 35445
rect 19242 35436 19248 35488
rect 19300 35476 19306 35488
rect 19981 35479 20039 35485
rect 19981 35476 19993 35479
rect 19300 35448 19993 35476
rect 19300 35436 19306 35448
rect 19981 35445 19993 35448
rect 20027 35445 20039 35479
rect 19981 35439 20039 35445
rect 20898 35436 20904 35488
rect 20956 35476 20962 35488
rect 21174 35476 21180 35488
rect 20956 35448 21180 35476
rect 20956 35436 20962 35448
rect 21174 35436 21180 35448
rect 21232 35436 21238 35488
rect 21269 35479 21327 35485
rect 21269 35445 21281 35479
rect 21315 35476 21327 35479
rect 21818 35476 21824 35488
rect 21315 35448 21824 35476
rect 21315 35445 21327 35448
rect 21269 35439 21327 35445
rect 21818 35436 21824 35448
rect 21876 35436 21882 35488
rect 22848 35476 22876 35516
rect 22925 35513 22937 35547
rect 22971 35544 22983 35547
rect 24213 35547 24271 35553
rect 22971 35516 24164 35544
rect 22971 35513 22983 35516
rect 22925 35507 22983 35513
rect 23382 35476 23388 35488
rect 22848 35448 23388 35476
rect 23382 35436 23388 35448
rect 23440 35436 23446 35488
rect 23566 35436 23572 35488
rect 23624 35476 23630 35488
rect 23937 35479 23995 35485
rect 23937 35476 23949 35479
rect 23624 35448 23949 35476
rect 23624 35436 23630 35448
rect 23937 35445 23949 35448
rect 23983 35445 23995 35479
rect 24136 35476 24164 35516
rect 24213 35513 24225 35547
rect 24259 35544 24271 35547
rect 25038 35544 25044 35556
rect 24259 35516 25044 35544
rect 24259 35513 24271 35516
rect 24213 35507 24271 35513
rect 25038 35504 25044 35516
rect 25096 35504 25102 35556
rect 26436 35544 26464 35584
rect 26878 35572 26884 35624
rect 26936 35612 26942 35624
rect 26973 35615 27031 35621
rect 26973 35612 26985 35615
rect 26936 35584 26985 35612
rect 26936 35572 26942 35584
rect 26973 35581 26985 35584
rect 27019 35581 27031 35615
rect 26973 35575 27031 35581
rect 29546 35572 29552 35624
rect 29604 35612 29610 35624
rect 31389 35615 31447 35621
rect 31389 35612 31401 35615
rect 29604 35584 31401 35612
rect 29604 35572 29610 35584
rect 31389 35581 31401 35584
rect 31435 35581 31447 35615
rect 31389 35575 31447 35581
rect 32416 35556 32444 35643
rect 33962 35640 33968 35652
rect 34020 35640 34026 35692
rect 34146 35680 34152 35692
rect 34107 35652 34152 35680
rect 34146 35640 34152 35652
rect 34204 35640 34210 35692
rect 34992 35689 35020 35720
rect 35342 35708 35348 35720
rect 35400 35708 35406 35760
rect 36740 35757 36768 35788
rect 37277 35785 37289 35788
rect 37323 35785 37335 35819
rect 37277 35779 37335 35785
rect 37734 35776 37740 35828
rect 37792 35816 37798 35828
rect 38841 35819 38899 35825
rect 38841 35816 38853 35819
rect 37792 35788 38853 35816
rect 37792 35776 37798 35788
rect 38841 35785 38853 35788
rect 38887 35785 38899 35819
rect 38841 35779 38899 35785
rect 39485 35819 39543 35825
rect 39485 35785 39497 35819
rect 39531 35816 39543 35819
rect 39666 35816 39672 35828
rect 39531 35788 39672 35816
rect 39531 35785 39543 35788
rect 39485 35779 39543 35785
rect 39666 35776 39672 35788
rect 39724 35776 39730 35828
rect 37458 35757 37464 35760
rect 36725 35751 36783 35757
rect 36725 35717 36737 35751
rect 36771 35717 36783 35751
rect 36725 35711 36783 35717
rect 37445 35751 37464 35757
rect 37445 35717 37457 35751
rect 37445 35711 37464 35717
rect 37458 35708 37464 35711
rect 37516 35708 37522 35760
rect 37642 35748 37648 35760
rect 37603 35720 37648 35748
rect 37642 35708 37648 35720
rect 37700 35748 37706 35760
rect 38562 35748 38568 35760
rect 37700 35720 38568 35748
rect 37700 35708 37706 35720
rect 38562 35708 38568 35720
rect 38620 35748 38626 35760
rect 40497 35751 40555 35757
rect 40497 35748 40509 35751
rect 38620 35720 40509 35748
rect 38620 35708 38626 35720
rect 40497 35717 40509 35720
rect 40543 35717 40555 35751
rect 40497 35711 40555 35717
rect 34967 35683 35025 35689
rect 34967 35649 34979 35683
rect 35013 35649 35025 35683
rect 34967 35643 35025 35649
rect 35066 35640 35072 35692
rect 35124 35680 35130 35692
rect 35253 35683 35311 35689
rect 35124 35652 35169 35680
rect 35124 35640 35130 35652
rect 35253 35649 35265 35683
rect 35299 35649 35311 35683
rect 36446 35680 36452 35692
rect 36407 35652 36452 35680
rect 35253 35643 35311 35649
rect 34057 35615 34115 35621
rect 34057 35581 34069 35615
rect 34103 35612 34115 35615
rect 34606 35612 34612 35624
rect 34103 35584 34612 35612
rect 34103 35581 34115 35584
rect 34057 35575 34115 35581
rect 34606 35572 34612 35584
rect 34664 35572 34670 35624
rect 35158 35612 35164 35624
rect 35119 35584 35164 35612
rect 35158 35572 35164 35584
rect 35216 35572 35222 35624
rect 35268 35612 35296 35643
rect 36446 35640 36452 35652
rect 36504 35640 36510 35692
rect 37476 35680 37504 35708
rect 38105 35683 38163 35689
rect 38105 35680 38117 35683
rect 37476 35652 38117 35680
rect 38105 35649 38117 35652
rect 38151 35649 38163 35683
rect 38286 35680 38292 35692
rect 38247 35652 38292 35680
rect 38105 35643 38163 35649
rect 38286 35640 38292 35652
rect 38344 35640 38350 35692
rect 38746 35680 38752 35692
rect 38707 35652 38752 35680
rect 38746 35640 38752 35652
rect 38804 35640 38810 35692
rect 38933 35683 38991 35689
rect 38933 35649 38945 35683
rect 38979 35680 38991 35683
rect 39758 35680 39764 35692
rect 38979 35652 39764 35680
rect 38979 35649 38991 35652
rect 38933 35643 38991 35649
rect 39758 35640 39764 35652
rect 39816 35640 39822 35692
rect 35268 35584 36032 35612
rect 27062 35544 27068 35556
rect 26436 35516 27068 35544
rect 27062 35504 27068 35516
rect 27120 35544 27126 35556
rect 27341 35547 27399 35553
rect 27341 35544 27353 35547
rect 27120 35516 27353 35544
rect 27120 35504 27126 35516
rect 27341 35513 27353 35516
rect 27387 35513 27399 35547
rect 27341 35507 27399 35513
rect 28994 35504 29000 35556
rect 29052 35544 29058 35556
rect 29089 35547 29147 35553
rect 29089 35544 29101 35547
rect 29052 35516 29101 35544
rect 29052 35504 29058 35516
rect 29089 35513 29101 35516
rect 29135 35544 29147 35547
rect 30282 35544 30288 35556
rect 29135 35516 30288 35544
rect 29135 35513 29147 35516
rect 29089 35507 29147 35513
rect 30282 35504 30288 35516
rect 30340 35544 30346 35556
rect 32122 35544 32128 35556
rect 30340 35516 32128 35544
rect 30340 35504 30346 35516
rect 32122 35504 32128 35516
rect 32180 35504 32186 35556
rect 32398 35504 32404 35556
rect 32456 35504 32462 35556
rect 33965 35547 34023 35553
rect 33965 35513 33977 35547
rect 34011 35544 34023 35547
rect 35176 35544 35204 35572
rect 34011 35516 35204 35544
rect 34011 35513 34023 35516
rect 33965 35507 34023 35513
rect 24578 35476 24584 35488
rect 24136 35448 24584 35476
rect 23937 35439 23995 35445
rect 24578 35436 24584 35448
rect 24636 35436 24642 35488
rect 28077 35479 28135 35485
rect 28077 35445 28089 35479
rect 28123 35476 28135 35479
rect 29546 35476 29552 35488
rect 28123 35448 29552 35476
rect 28123 35445 28135 35448
rect 28077 35439 28135 35445
rect 29546 35436 29552 35448
rect 29604 35436 29610 35488
rect 30926 35476 30932 35488
rect 30887 35448 30932 35476
rect 30926 35436 30932 35448
rect 30984 35436 30990 35488
rect 32674 35436 32680 35488
rect 32732 35476 32738 35488
rect 32769 35479 32827 35485
rect 32769 35476 32781 35479
rect 32732 35448 32781 35476
rect 32732 35436 32738 35448
rect 32769 35445 32781 35448
rect 32815 35445 32827 35479
rect 33226 35476 33232 35488
rect 33187 35448 33232 35476
rect 32769 35439 32827 35445
rect 33226 35436 33232 35448
rect 33284 35436 33290 35488
rect 34054 35436 34060 35488
rect 34112 35476 34118 35488
rect 35805 35479 35863 35485
rect 35805 35476 35817 35479
rect 34112 35448 35817 35476
rect 34112 35436 34118 35448
rect 35805 35445 35817 35448
rect 35851 35445 35863 35479
rect 36004 35476 36032 35584
rect 36170 35572 36176 35624
rect 36228 35612 36234 35624
rect 38197 35615 38255 35621
rect 38197 35612 38209 35615
rect 36228 35584 38209 35612
rect 36228 35572 36234 35584
rect 38197 35581 38209 35584
rect 38243 35581 38255 35615
rect 38197 35575 38255 35581
rect 36725 35547 36783 35553
rect 36725 35544 36737 35547
rect 36648 35516 36737 35544
rect 36648 35476 36676 35516
rect 36725 35513 36737 35516
rect 36771 35513 36783 35547
rect 36725 35507 36783 35513
rect 36004 35448 36676 35476
rect 37461 35479 37519 35485
rect 35805 35439 35863 35445
rect 37461 35445 37473 35479
rect 37507 35476 37519 35479
rect 37734 35476 37740 35488
rect 37507 35448 37740 35476
rect 37507 35445 37519 35448
rect 37461 35439 37519 35445
rect 37734 35436 37740 35448
rect 37792 35476 37798 35488
rect 38378 35476 38384 35488
rect 37792 35448 38384 35476
rect 37792 35436 37798 35448
rect 38378 35436 38384 35448
rect 38436 35476 38442 35488
rect 40037 35479 40095 35485
rect 40037 35476 40049 35479
rect 38436 35448 40049 35476
rect 38436 35436 38442 35448
rect 40037 35445 40049 35448
rect 40083 35445 40095 35479
rect 40037 35439 40095 35445
rect 1104 35386 54372 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 54372 35386
rect 1104 35312 54372 35334
rect 16945 35275 17003 35281
rect 16945 35241 16957 35275
rect 16991 35272 17003 35275
rect 18230 35272 18236 35284
rect 16991 35244 18236 35272
rect 16991 35241 17003 35244
rect 16945 35235 17003 35241
rect 18230 35232 18236 35244
rect 18288 35232 18294 35284
rect 20622 35232 20628 35284
rect 20680 35272 20686 35284
rect 20809 35275 20867 35281
rect 20809 35272 20821 35275
rect 20680 35244 20821 35272
rect 20680 35232 20686 35244
rect 20809 35241 20821 35244
rect 20855 35241 20867 35275
rect 20809 35235 20867 35241
rect 20898 35232 20904 35284
rect 20956 35272 20962 35284
rect 20993 35275 21051 35281
rect 20993 35272 21005 35275
rect 20956 35244 21005 35272
rect 20956 35232 20962 35244
rect 20993 35241 21005 35244
rect 21039 35241 21051 35275
rect 20993 35235 21051 35241
rect 21082 35232 21088 35284
rect 21140 35272 21146 35284
rect 21266 35272 21272 35284
rect 21140 35244 21272 35272
rect 21140 35232 21146 35244
rect 21266 35232 21272 35244
rect 21324 35272 21330 35284
rect 21729 35275 21787 35281
rect 21729 35272 21741 35275
rect 21324 35244 21741 35272
rect 21324 35232 21330 35244
rect 21729 35241 21741 35244
rect 21775 35241 21787 35275
rect 21729 35235 21787 35241
rect 23382 35232 23388 35284
rect 23440 35272 23446 35284
rect 23753 35275 23811 35281
rect 23753 35272 23765 35275
rect 23440 35244 23765 35272
rect 23440 35232 23446 35244
rect 23753 35241 23765 35244
rect 23799 35272 23811 35275
rect 23842 35272 23848 35284
rect 23799 35244 23848 35272
rect 23799 35241 23811 35244
rect 23753 35235 23811 35241
rect 23842 35232 23848 35244
rect 23900 35232 23906 35284
rect 24394 35232 24400 35284
rect 24452 35272 24458 35284
rect 24489 35275 24547 35281
rect 24489 35272 24501 35275
rect 24452 35244 24501 35272
rect 24452 35232 24458 35244
rect 24489 35241 24501 35244
rect 24535 35241 24547 35275
rect 24762 35272 24768 35284
rect 24723 35244 24768 35272
rect 24489 35235 24547 35241
rect 24762 35232 24768 35244
rect 24820 35232 24826 35284
rect 26145 35275 26203 35281
rect 26145 35241 26157 35275
rect 26191 35272 26203 35275
rect 28350 35272 28356 35284
rect 26191 35244 28356 35272
rect 26191 35241 26203 35244
rect 26145 35235 26203 35241
rect 28350 35232 28356 35244
rect 28408 35272 28414 35284
rect 28813 35275 28871 35281
rect 28813 35272 28825 35275
rect 28408 35244 28825 35272
rect 28408 35232 28414 35244
rect 28813 35241 28825 35244
rect 28859 35272 28871 35275
rect 28859 35244 28994 35272
rect 28859 35241 28871 35244
rect 28813 35235 28871 35241
rect 19058 35204 19064 35216
rect 17052 35176 19064 35204
rect 16942 35096 16948 35148
rect 17000 35136 17006 35148
rect 17052 35136 17080 35176
rect 19058 35164 19064 35176
rect 19116 35164 19122 35216
rect 22925 35207 22983 35213
rect 22925 35173 22937 35207
rect 22971 35173 22983 35207
rect 22925 35167 22983 35173
rect 17000 35108 17080 35136
rect 17000 35096 17006 35108
rect 15841 35071 15899 35077
rect 15841 35037 15853 35071
rect 15887 35068 15899 35071
rect 16758 35068 16764 35080
rect 15887 35040 16764 35068
rect 15887 35037 15899 35040
rect 15841 35031 15899 35037
rect 16758 35028 16764 35040
rect 16816 35068 16822 35080
rect 17052 35077 17080 35108
rect 17402 35096 17408 35148
rect 17460 35136 17466 35148
rect 17497 35139 17555 35145
rect 17497 35136 17509 35139
rect 17460 35108 17509 35136
rect 17460 35096 17466 35108
rect 17497 35105 17509 35108
rect 17543 35136 17555 35139
rect 17862 35136 17868 35148
rect 17543 35108 17868 35136
rect 17543 35105 17555 35108
rect 17497 35099 17555 35105
rect 17862 35096 17868 35108
rect 17920 35096 17926 35148
rect 17954 35096 17960 35148
rect 18012 35136 18018 35148
rect 18012 35108 18736 35136
rect 18012 35096 18018 35108
rect 16853 35071 16911 35077
rect 16853 35068 16865 35071
rect 16816 35040 16865 35068
rect 16816 35028 16822 35040
rect 16853 35037 16865 35040
rect 16899 35037 16911 35071
rect 16853 35031 16911 35037
rect 17037 35071 17095 35077
rect 17037 35037 17049 35071
rect 17083 35037 17095 35071
rect 17037 35031 17095 35037
rect 17586 35028 17592 35080
rect 17644 35068 17650 35080
rect 17681 35071 17739 35077
rect 17681 35068 17693 35071
rect 17644 35040 17693 35068
rect 17644 35028 17650 35040
rect 17681 35037 17693 35040
rect 17727 35037 17739 35071
rect 18046 35068 18052 35080
rect 18007 35040 18052 35068
rect 17681 35031 17739 35037
rect 18046 35028 18052 35040
rect 18104 35028 18110 35080
rect 18506 35068 18512 35080
rect 18467 35040 18512 35068
rect 18506 35028 18512 35040
rect 18564 35028 18570 35080
rect 18708 35077 18736 35108
rect 19242 35096 19248 35148
rect 19300 35136 19306 35148
rect 19300 35108 19840 35136
rect 19300 35096 19306 35108
rect 18693 35071 18751 35077
rect 18693 35037 18705 35071
rect 18739 35037 18751 35071
rect 19426 35068 19432 35080
rect 19387 35040 19432 35068
rect 18693 35031 18751 35037
rect 19426 35028 19432 35040
rect 19484 35028 19490 35080
rect 19812 35077 19840 35108
rect 20714 35096 20720 35148
rect 20772 35136 20778 35148
rect 21085 35139 21143 35145
rect 21085 35136 21097 35139
rect 20772 35108 21097 35136
rect 20772 35096 20778 35108
rect 21085 35105 21097 35108
rect 21131 35105 21143 35139
rect 21821 35139 21879 35145
rect 21821 35136 21833 35139
rect 21085 35099 21143 35105
rect 21468 35108 21833 35136
rect 19797 35071 19855 35077
rect 19797 35037 19809 35071
rect 19843 35037 19855 35071
rect 19797 35031 19855 35037
rect 19889 35071 19947 35077
rect 19889 35037 19901 35071
rect 19935 35068 19947 35071
rect 19978 35068 19984 35080
rect 19935 35040 19984 35068
rect 19935 35037 19947 35040
rect 19889 35031 19947 35037
rect 19978 35028 19984 35040
rect 20036 35028 20042 35080
rect 20622 35028 20628 35080
rect 20680 35068 20686 35080
rect 20993 35071 21051 35077
rect 20993 35068 21005 35071
rect 20680 35040 21005 35068
rect 20680 35028 20686 35040
rect 20993 35037 21005 35040
rect 21039 35068 21051 35071
rect 21468 35068 21496 35108
rect 21821 35105 21833 35108
rect 21867 35136 21879 35139
rect 21910 35136 21916 35148
rect 21867 35108 21916 35136
rect 21867 35105 21879 35108
rect 21821 35099 21879 35105
rect 21910 35096 21916 35108
rect 21968 35096 21974 35148
rect 22738 35136 22744 35148
rect 22699 35108 22744 35136
rect 22738 35096 22744 35108
rect 22796 35096 22802 35148
rect 22940 35136 22968 35167
rect 24118 35164 24124 35216
rect 24176 35204 24182 35216
rect 25866 35204 25872 35216
rect 24176 35176 25872 35204
rect 24176 35164 24182 35176
rect 25866 35164 25872 35176
rect 25924 35164 25930 35216
rect 26605 35139 26663 35145
rect 22940 35108 25084 35136
rect 21039 35040 21496 35068
rect 21729 35071 21787 35077
rect 21039 35037 21051 35040
rect 20993 35031 21051 35037
rect 21729 35037 21741 35071
rect 21775 35037 21787 35071
rect 22554 35068 22560 35080
rect 22515 35040 22560 35068
rect 21729 35031 21787 35037
rect 18601 35003 18659 35009
rect 18601 34969 18613 35003
rect 18647 35000 18659 35003
rect 19334 35000 19340 35012
rect 18647 34972 19340 35000
rect 18647 34969 18659 34972
rect 18601 34963 18659 34969
rect 19334 34960 19340 34972
rect 19392 35000 19398 35012
rect 19567 35003 19625 35009
rect 19567 35000 19579 35003
rect 19392 34972 19579 35000
rect 19392 34960 19398 34972
rect 19567 34969 19579 34972
rect 19613 34969 19625 35003
rect 19567 34963 19625 34969
rect 19705 35003 19763 35009
rect 19705 34969 19717 35003
rect 19751 34969 19763 35003
rect 21266 35000 21272 35012
rect 21227 34972 21272 35000
rect 19705 34963 19763 34969
rect 15930 34892 15936 34944
rect 15988 34932 15994 34944
rect 16301 34935 16359 34941
rect 16301 34932 16313 34935
rect 15988 34904 16313 34932
rect 15988 34892 15994 34904
rect 16301 34901 16313 34904
rect 16347 34901 16359 34935
rect 16301 34895 16359 34901
rect 19150 34892 19156 34944
rect 19208 34932 19214 34944
rect 19720 34932 19748 34963
rect 21266 34960 21272 34972
rect 21324 35000 21330 35012
rect 21744 35000 21772 35031
rect 22554 35028 22560 35040
rect 22612 35028 22618 35080
rect 22922 35068 22928 35080
rect 22883 35040 22928 35068
rect 22922 35028 22928 35040
rect 22980 35028 22986 35080
rect 23842 35028 23848 35080
rect 23900 35068 23906 35080
rect 24765 35071 24823 35077
rect 24765 35068 24777 35071
rect 23900 35040 24777 35068
rect 23900 35028 23906 35040
rect 24765 35037 24777 35040
rect 24811 35037 24823 35071
rect 24765 35031 24823 35037
rect 24949 35071 25007 35077
rect 24949 35037 24961 35071
rect 24995 35037 25007 35071
rect 25056 35068 25084 35108
rect 26605 35105 26617 35139
rect 26651 35136 26663 35139
rect 26970 35136 26976 35148
rect 26651 35108 26976 35136
rect 26651 35105 26663 35108
rect 26605 35099 26663 35105
rect 26970 35096 26976 35108
rect 27028 35096 27034 35148
rect 28966 35136 28994 35244
rect 31294 35232 31300 35284
rect 31352 35272 31358 35284
rect 35802 35272 35808 35284
rect 31352 35244 35808 35272
rect 31352 35232 31358 35244
rect 35802 35232 35808 35244
rect 35860 35232 35866 35284
rect 37458 35272 37464 35284
rect 37419 35244 37464 35272
rect 37458 35232 37464 35244
rect 37516 35232 37522 35284
rect 38381 35275 38439 35281
rect 38381 35241 38393 35275
rect 38427 35272 38439 35275
rect 39758 35272 39764 35284
rect 38427 35244 39764 35272
rect 38427 35241 38439 35244
rect 38381 35235 38439 35241
rect 29086 35164 29092 35216
rect 29144 35204 29150 35216
rect 29641 35207 29699 35213
rect 29641 35204 29653 35207
rect 29144 35176 29653 35204
rect 29144 35164 29150 35176
rect 29641 35173 29653 35176
rect 29687 35173 29699 35207
rect 29641 35167 29699 35173
rect 33410 35164 33416 35216
rect 33468 35204 33474 35216
rect 33781 35207 33839 35213
rect 33781 35204 33793 35207
rect 33468 35176 33793 35204
rect 33468 35164 33474 35176
rect 33781 35173 33793 35176
rect 33827 35204 33839 35207
rect 36173 35207 36231 35213
rect 36173 35204 36185 35207
rect 33827 35176 36185 35204
rect 33827 35173 33839 35176
rect 33781 35167 33839 35173
rect 36173 35173 36185 35176
rect 36219 35204 36231 35207
rect 36538 35204 36544 35216
rect 36219 35176 36544 35204
rect 36219 35173 36231 35176
rect 36173 35167 36231 35173
rect 29178 35136 29184 35148
rect 28966 35108 29184 35136
rect 29178 35096 29184 35108
rect 29236 35136 29242 35148
rect 36078 35136 36084 35148
rect 29236 35108 29960 35136
rect 29236 35096 29242 35108
rect 26881 35071 26939 35077
rect 26881 35068 26893 35071
rect 25056 35040 26893 35068
rect 24949 35031 25007 35037
rect 26881 35037 26893 35040
rect 26927 35037 26939 35071
rect 26881 35031 26939 35037
rect 21324 34972 21772 35000
rect 24964 35000 24992 35031
rect 27154 35028 27160 35080
rect 27212 35068 27218 35080
rect 29932 35077 29960 35108
rect 33888 35108 36084 35136
rect 28261 35071 28319 35077
rect 28261 35068 28273 35071
rect 27212 35040 28273 35068
rect 27212 35028 27218 35040
rect 28261 35037 28273 35040
rect 28307 35068 28319 35071
rect 29917 35071 29975 35077
rect 28307 35040 29776 35068
rect 28307 35037 28319 35040
rect 28261 35031 28319 35037
rect 25038 35000 25044 35012
rect 24964 34972 25044 35000
rect 21324 34960 21330 34972
rect 25038 34960 25044 34972
rect 25096 34960 25102 35012
rect 29638 35000 29644 35012
rect 29599 34972 29644 35000
rect 29638 34960 29644 34972
rect 29696 34960 29702 35012
rect 29748 35000 29776 35040
rect 29917 35037 29929 35071
rect 29963 35037 29975 35071
rect 29917 35031 29975 35037
rect 31685 35071 31743 35077
rect 31685 35037 31697 35071
rect 31731 35068 31743 35071
rect 31846 35068 31852 35080
rect 31731 35040 31852 35068
rect 31731 35037 31743 35040
rect 31685 35031 31743 35037
rect 31846 35028 31852 35040
rect 31904 35028 31910 35080
rect 31941 35071 31999 35077
rect 31941 35037 31953 35071
rect 31987 35068 31999 35071
rect 32122 35068 32128 35080
rect 31987 35040 32128 35068
rect 31987 35037 31999 35040
rect 31941 35031 31999 35037
rect 32122 35028 32128 35040
rect 32180 35068 32186 35080
rect 32674 35077 32680 35080
rect 32401 35071 32459 35077
rect 32401 35068 32413 35071
rect 32180 35040 32413 35068
rect 32180 35028 32186 35040
rect 32401 35037 32413 35040
rect 32447 35037 32459 35071
rect 32668 35068 32680 35077
rect 32635 35040 32680 35068
rect 32401 35031 32459 35037
rect 32668 35031 32680 35040
rect 32674 35028 32680 35031
rect 32732 35028 32738 35080
rect 33888 35000 33916 35108
rect 36078 35096 36084 35108
rect 36136 35096 36142 35148
rect 34606 35028 34612 35080
rect 34664 35068 34670 35080
rect 34701 35071 34759 35077
rect 34701 35068 34713 35071
rect 34664 35040 34713 35068
rect 34664 35028 34670 35040
rect 34701 35037 34713 35040
rect 34747 35068 34759 35071
rect 34790 35068 34796 35080
rect 34747 35040 34796 35068
rect 34747 35037 34759 35040
rect 34701 35031 34759 35037
rect 34790 35028 34796 35040
rect 34848 35028 34854 35080
rect 35342 35028 35348 35080
rect 35400 35068 35406 35080
rect 35437 35071 35495 35077
rect 35437 35068 35449 35071
rect 35400 35040 35449 35068
rect 35400 35028 35406 35040
rect 35437 35037 35449 35040
rect 35483 35068 35495 35071
rect 35526 35068 35532 35080
rect 35483 35040 35532 35068
rect 35483 35037 35495 35040
rect 35437 35031 35495 35037
rect 35526 35028 35532 35040
rect 35584 35028 35590 35080
rect 35621 35071 35679 35077
rect 35621 35037 35633 35071
rect 35667 35068 35679 35071
rect 36188 35068 36216 35167
rect 36538 35164 36544 35176
rect 36596 35204 36602 35216
rect 36725 35207 36783 35213
rect 36725 35204 36737 35207
rect 36596 35176 36737 35204
rect 36596 35164 36602 35176
rect 36725 35173 36737 35176
rect 36771 35204 36783 35207
rect 38396 35204 38424 35235
rect 39758 35232 39764 35244
rect 39816 35272 39822 35284
rect 39853 35275 39911 35281
rect 39853 35272 39865 35275
rect 39816 35244 39865 35272
rect 39816 35232 39822 35244
rect 39853 35241 39865 35244
rect 39899 35241 39911 35275
rect 39853 35235 39911 35241
rect 36771 35176 38424 35204
rect 36771 35173 36783 35176
rect 36725 35167 36783 35173
rect 37826 35068 37832 35080
rect 35667 35040 36216 35068
rect 36464 35040 37832 35068
rect 35667 35037 35679 35040
rect 35621 35031 35679 35037
rect 36464 35012 36492 35040
rect 37826 35028 37832 35040
rect 37884 35028 37890 35080
rect 36446 35000 36452 35012
rect 29748 34972 33916 35000
rect 34900 34972 36452 35000
rect 20070 34932 20076 34944
rect 19208 34904 19748 34932
rect 20031 34904 20076 34932
rect 19208 34892 19214 34904
rect 20070 34892 20076 34904
rect 20128 34892 20134 34944
rect 22097 34935 22155 34941
rect 22097 34901 22109 34935
rect 22143 34932 22155 34935
rect 22649 34935 22707 34941
rect 22649 34932 22661 34935
rect 22143 34904 22661 34932
rect 22143 34901 22155 34904
rect 22097 34895 22155 34901
rect 22649 34901 22661 34904
rect 22695 34901 22707 34935
rect 22649 34895 22707 34901
rect 25593 34935 25651 34941
rect 25593 34901 25605 34935
rect 25639 34932 25651 34935
rect 25774 34932 25780 34944
rect 25639 34904 25780 34932
rect 25639 34901 25651 34904
rect 25593 34895 25651 34901
rect 25774 34892 25780 34904
rect 25832 34932 25838 34944
rect 27706 34932 27712 34944
rect 25832 34904 27712 34932
rect 25832 34892 25838 34904
rect 27706 34892 27712 34904
rect 27764 34892 27770 34944
rect 29546 34892 29552 34944
rect 29604 34932 29610 34944
rect 29825 34935 29883 34941
rect 29825 34932 29837 34935
rect 29604 34904 29837 34932
rect 29604 34892 29610 34904
rect 29825 34901 29837 34904
rect 29871 34901 29883 34935
rect 30558 34932 30564 34944
rect 30519 34904 30564 34932
rect 29825 34895 29883 34901
rect 30558 34892 30564 34904
rect 30616 34892 30622 34944
rect 31386 34892 31392 34944
rect 31444 34932 31450 34944
rect 31662 34932 31668 34944
rect 31444 34904 31668 34932
rect 31444 34892 31450 34904
rect 31662 34892 31668 34904
rect 31720 34932 31726 34944
rect 33226 34932 33232 34944
rect 31720 34904 33232 34932
rect 31720 34892 31726 34904
rect 33226 34892 33232 34904
rect 33284 34892 33290 34944
rect 34330 34892 34336 34944
rect 34388 34932 34394 34944
rect 34900 34941 34928 34972
rect 36446 34960 36452 34972
rect 36504 34960 36510 35012
rect 37642 35000 37648 35012
rect 37603 34972 37648 35000
rect 37642 34960 37648 34972
rect 37700 34960 37706 35012
rect 52917 35003 52975 35009
rect 52917 34969 52929 35003
rect 52963 35000 52975 35003
rect 53558 35000 53564 35012
rect 52963 34972 53564 35000
rect 52963 34969 52975 34972
rect 52917 34963 52975 34969
rect 53558 34960 53564 34972
rect 53616 34960 53622 35012
rect 34885 34935 34943 34941
rect 34885 34932 34897 34935
rect 34388 34904 34897 34932
rect 34388 34892 34394 34904
rect 34885 34901 34897 34904
rect 34931 34901 34943 34935
rect 34885 34895 34943 34901
rect 35342 34892 35348 34944
rect 35400 34932 35406 34944
rect 35437 34935 35495 34941
rect 35437 34932 35449 34935
rect 35400 34904 35449 34932
rect 35400 34892 35406 34904
rect 35437 34901 35449 34904
rect 35483 34901 35495 34935
rect 35437 34895 35495 34901
rect 36630 34892 36636 34944
rect 36688 34932 36694 34944
rect 37660 34932 37688 34960
rect 38838 34932 38844 34944
rect 36688 34904 37688 34932
rect 38799 34904 38844 34932
rect 36688 34892 36694 34904
rect 38838 34892 38844 34904
rect 38896 34892 38902 34944
rect 52454 34892 52460 34944
rect 52512 34932 52518 34944
rect 53469 34935 53527 34941
rect 53469 34932 53481 34935
rect 52512 34904 53481 34932
rect 52512 34892 52518 34904
rect 53469 34901 53481 34904
rect 53515 34901 53527 34935
rect 53469 34895 53527 34901
rect 1104 34842 54372 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 54372 34842
rect 1104 34768 54372 34790
rect 15470 34728 15476 34740
rect 15431 34700 15476 34728
rect 15470 34688 15476 34700
rect 15528 34688 15534 34740
rect 16117 34731 16175 34737
rect 16117 34697 16129 34731
rect 16163 34728 16175 34731
rect 16942 34728 16948 34740
rect 16163 34700 16948 34728
rect 16163 34697 16175 34700
rect 16117 34691 16175 34697
rect 16942 34688 16948 34700
rect 17000 34688 17006 34740
rect 17589 34731 17647 34737
rect 17589 34697 17601 34731
rect 17635 34728 17647 34731
rect 18506 34728 18512 34740
rect 17635 34700 18512 34728
rect 17635 34697 17647 34700
rect 17589 34691 17647 34697
rect 18506 34688 18512 34700
rect 18564 34688 18570 34740
rect 18874 34728 18880 34740
rect 18835 34700 18880 34728
rect 18874 34688 18880 34700
rect 18932 34688 18938 34740
rect 21269 34731 21327 34737
rect 21269 34697 21281 34731
rect 21315 34728 21327 34731
rect 22554 34728 22560 34740
rect 21315 34700 22560 34728
rect 21315 34697 21327 34700
rect 21269 34691 21327 34697
rect 22554 34688 22560 34700
rect 22612 34688 22618 34740
rect 22922 34688 22928 34740
rect 22980 34728 22986 34740
rect 25133 34731 25191 34737
rect 25133 34728 25145 34731
rect 22980 34700 25145 34728
rect 22980 34688 22986 34700
rect 25133 34697 25145 34700
rect 25179 34697 25191 34731
rect 25133 34691 25191 34697
rect 25314 34688 25320 34740
rect 25372 34688 25378 34740
rect 26418 34728 26424 34740
rect 26331 34700 26424 34728
rect 26418 34688 26424 34700
rect 26476 34728 26482 34740
rect 27154 34728 27160 34740
rect 26476 34700 27160 34728
rect 26476 34688 26482 34700
rect 27154 34688 27160 34700
rect 27212 34688 27218 34740
rect 30742 34728 30748 34740
rect 30703 34700 30748 34728
rect 30742 34688 30748 34700
rect 30800 34688 30806 34740
rect 31474 34731 31532 34737
rect 31474 34697 31486 34731
rect 31520 34728 31532 34731
rect 32398 34728 32404 34740
rect 31520 34700 32404 34728
rect 31520 34697 31532 34700
rect 31474 34691 31532 34697
rect 32398 34688 32404 34700
rect 32456 34688 32462 34740
rect 34149 34731 34207 34737
rect 34149 34728 34161 34731
rect 32508 34700 34161 34728
rect 16761 34663 16819 34669
rect 16761 34629 16773 34663
rect 16807 34660 16819 34663
rect 16850 34660 16856 34672
rect 16807 34632 16856 34660
rect 16807 34629 16819 34632
rect 16761 34623 16819 34629
rect 16850 34620 16856 34632
rect 16908 34620 16914 34672
rect 17221 34663 17279 34669
rect 17221 34629 17233 34663
rect 17267 34629 17279 34663
rect 17221 34623 17279 34629
rect 17437 34663 17495 34669
rect 17437 34629 17449 34663
rect 17483 34660 17495 34663
rect 18046 34660 18052 34672
rect 17483 34632 18052 34660
rect 17483 34629 17495 34632
rect 17437 34623 17495 34629
rect 1578 34552 1584 34604
rect 1636 34592 1642 34604
rect 1857 34595 1915 34601
rect 1857 34592 1869 34595
rect 1636 34564 1869 34592
rect 1636 34552 1642 34564
rect 1857 34561 1869 34564
rect 1903 34561 1915 34595
rect 17236 34592 17264 34623
rect 18046 34620 18052 34632
rect 18104 34620 18110 34672
rect 19058 34660 19064 34672
rect 19019 34632 19064 34660
rect 19058 34620 19064 34632
rect 19116 34620 19122 34672
rect 22278 34620 22284 34672
rect 22336 34660 22342 34672
rect 22373 34663 22431 34669
rect 22373 34660 22385 34663
rect 22336 34632 22385 34660
rect 22336 34620 22342 34632
rect 22373 34629 22385 34632
rect 22419 34629 22431 34663
rect 22373 34623 22431 34629
rect 23569 34663 23627 34669
rect 23569 34629 23581 34663
rect 23615 34660 23627 34663
rect 23658 34660 23664 34672
rect 23615 34632 23664 34660
rect 23615 34629 23627 34632
rect 23569 34623 23627 34629
rect 23658 34620 23664 34632
rect 23716 34660 23722 34672
rect 25038 34660 25044 34672
rect 23716 34632 25044 34660
rect 23716 34620 23722 34632
rect 25038 34620 25044 34632
rect 25096 34620 25102 34672
rect 25332 34660 25360 34688
rect 25412 34663 25470 34669
rect 25412 34660 25424 34663
rect 25332 34632 25424 34660
rect 25412 34629 25424 34632
rect 25458 34629 25470 34663
rect 25412 34623 25470 34629
rect 25866 34620 25872 34672
rect 25924 34660 25930 34672
rect 28629 34663 28687 34669
rect 28629 34660 28641 34663
rect 25924 34632 28641 34660
rect 25924 34620 25930 34632
rect 28629 34629 28641 34632
rect 28675 34629 28687 34663
rect 28629 34623 28687 34629
rect 30466 34620 30472 34672
rect 30524 34660 30530 34672
rect 31386 34660 31392 34672
rect 30524 34632 31392 34660
rect 30524 34620 30530 34632
rect 31386 34620 31392 34632
rect 31444 34620 31450 34672
rect 31573 34663 31631 34669
rect 31573 34629 31585 34663
rect 31619 34660 31631 34663
rect 32125 34663 32183 34669
rect 32125 34660 32137 34663
rect 31619 34632 32137 34660
rect 31619 34629 31631 34632
rect 31573 34623 31631 34629
rect 32125 34629 32137 34632
rect 32171 34629 32183 34663
rect 32125 34623 32183 34629
rect 17586 34592 17592 34604
rect 17236 34564 17592 34592
rect 1857 34555 1915 34561
rect 17586 34552 17592 34564
rect 17644 34552 17650 34604
rect 18230 34592 18236 34604
rect 18191 34564 18236 34592
rect 18230 34552 18236 34564
rect 18288 34552 18294 34604
rect 19245 34595 19303 34601
rect 19245 34592 19257 34595
rect 18340 34564 19257 34592
rect 2038 34524 2044 34536
rect 1999 34496 2044 34524
rect 2038 34484 2044 34496
rect 2096 34484 2102 34536
rect 16758 34484 16764 34536
rect 16816 34524 16822 34536
rect 18340 34524 18368 34564
rect 19245 34561 19257 34564
rect 19291 34561 19303 34595
rect 19245 34555 19303 34561
rect 19426 34552 19432 34604
rect 19484 34592 19490 34604
rect 19889 34595 19947 34601
rect 19889 34592 19901 34595
rect 19484 34564 19901 34592
rect 19484 34552 19490 34564
rect 19889 34561 19901 34564
rect 19935 34561 19947 34595
rect 19889 34555 19947 34561
rect 20622 34552 20628 34604
rect 20680 34592 20686 34604
rect 20993 34595 21051 34601
rect 20993 34592 21005 34595
rect 20680 34564 21005 34592
rect 20680 34552 20686 34564
rect 20993 34561 21005 34564
rect 21039 34561 21051 34595
rect 20993 34555 21051 34561
rect 21082 34552 21088 34604
rect 21140 34592 21146 34604
rect 22189 34595 22247 34601
rect 22189 34592 22201 34595
rect 21140 34564 21185 34592
rect 22066 34564 22201 34592
rect 21140 34552 21146 34564
rect 16816 34496 18368 34524
rect 16816 34484 16822 34496
rect 18414 34484 18420 34536
rect 18472 34524 18478 34536
rect 18472 34496 18517 34524
rect 18472 34484 18478 34496
rect 19334 34484 19340 34536
rect 19392 34524 19398 34536
rect 19794 34524 19800 34536
rect 19392 34496 19800 34524
rect 19392 34484 19398 34496
rect 19794 34484 19800 34496
rect 19852 34484 19858 34536
rect 21266 34524 21272 34536
rect 21179 34496 21272 34524
rect 21266 34484 21272 34496
rect 21324 34484 21330 34536
rect 15470 34416 15476 34468
rect 15528 34456 15534 34468
rect 16390 34456 16396 34468
rect 15528 34428 16396 34456
rect 15528 34416 15534 34428
rect 16390 34416 16396 34428
rect 16448 34456 16454 34468
rect 18432 34456 18460 34484
rect 16448 34428 18460 34456
rect 20257 34459 20315 34465
rect 16448 34416 16454 34428
rect 20257 34425 20269 34459
rect 20303 34456 20315 34459
rect 21284 34456 21312 34484
rect 22066 34468 22094 34564
rect 22189 34561 22201 34564
rect 22235 34592 22247 34595
rect 24670 34592 24676 34604
rect 22235 34564 24676 34592
rect 22235 34561 22247 34564
rect 22189 34555 22247 34561
rect 24670 34552 24676 34564
rect 24728 34552 24734 34604
rect 24854 34552 24860 34604
rect 24912 34592 24918 34604
rect 25271 34595 25329 34601
rect 25271 34592 25283 34595
rect 24912 34564 25283 34592
rect 24912 34552 24918 34564
rect 25271 34561 25283 34564
rect 25317 34561 25329 34595
rect 25498 34592 25504 34604
rect 25459 34564 25504 34592
rect 25271 34555 25329 34561
rect 25498 34552 25504 34564
rect 25556 34552 25562 34604
rect 25629 34595 25687 34601
rect 25629 34561 25641 34595
rect 25675 34561 25687 34595
rect 25774 34592 25780 34604
rect 25735 34564 25780 34592
rect 25629 34555 25687 34561
rect 20303 34428 21312 34456
rect 20303 34425 20315 34428
rect 20257 34419 20315 34425
rect 22002 34416 22008 34468
rect 22060 34428 22094 34468
rect 24121 34459 24179 34465
rect 22060 34416 22066 34428
rect 24121 34425 24133 34459
rect 24167 34456 24179 34459
rect 25644 34456 25672 34555
rect 25774 34552 25780 34564
rect 25832 34552 25838 34604
rect 26878 34552 26884 34604
rect 26936 34592 26942 34604
rect 26973 34595 27031 34601
rect 26973 34592 26985 34595
rect 26936 34564 26985 34592
rect 26936 34552 26942 34564
rect 26973 34561 26985 34564
rect 27019 34561 27031 34595
rect 26973 34555 27031 34561
rect 27157 34595 27215 34601
rect 27157 34561 27169 34595
rect 27203 34561 27215 34595
rect 28810 34592 28816 34604
rect 28771 34564 28816 34592
rect 27157 34555 27215 34561
rect 26050 34484 26056 34536
rect 26108 34524 26114 34536
rect 27172 34524 27200 34555
rect 28810 34552 28816 34564
rect 28868 34552 28874 34604
rect 29086 34592 29092 34604
rect 29047 34564 29092 34592
rect 29086 34552 29092 34564
rect 29144 34552 29150 34604
rect 29825 34595 29883 34601
rect 29825 34561 29837 34595
rect 29871 34561 29883 34595
rect 29825 34555 29883 34561
rect 28994 34524 29000 34536
rect 26108 34496 27200 34524
rect 28907 34496 29000 34524
rect 26108 34484 26114 34496
rect 28994 34484 29000 34496
rect 29052 34524 29058 34536
rect 29840 34524 29868 34555
rect 30282 34552 30288 34604
rect 30340 34592 30346 34604
rect 30650 34592 30656 34604
rect 30340 34564 30656 34592
rect 30340 34552 30346 34564
rect 30650 34552 30656 34564
rect 30708 34552 30714 34604
rect 30837 34595 30895 34601
rect 30837 34561 30849 34595
rect 30883 34561 30895 34595
rect 31294 34592 31300 34604
rect 31255 34564 31300 34592
rect 30837 34555 30895 34561
rect 29052 34496 29868 34524
rect 29052 34484 29058 34496
rect 29914 34484 29920 34536
rect 29972 34524 29978 34536
rect 30190 34524 30196 34536
rect 29972 34496 30017 34524
rect 30151 34496 30196 34524
rect 29972 34484 29978 34496
rect 30190 34484 30196 34496
rect 30248 34484 30254 34536
rect 30852 34524 30880 34555
rect 31294 34552 31300 34564
rect 31352 34552 31358 34604
rect 32398 34592 32404 34604
rect 32359 34564 32404 34592
rect 32398 34552 32404 34564
rect 32456 34552 32462 34604
rect 32508 34601 32536 34700
rect 34149 34697 34161 34700
rect 34195 34697 34207 34731
rect 36538 34728 36544 34740
rect 36499 34700 36544 34728
rect 34149 34691 34207 34697
rect 36538 34688 36544 34700
rect 36596 34688 36602 34740
rect 37553 34731 37611 34737
rect 37553 34697 37565 34731
rect 37599 34728 37611 34731
rect 38286 34728 38292 34740
rect 37599 34700 38292 34728
rect 37599 34697 37611 34700
rect 37553 34691 37611 34697
rect 38286 34688 38292 34700
rect 38344 34688 38350 34740
rect 38657 34731 38715 34737
rect 38657 34697 38669 34731
rect 38703 34728 38715 34731
rect 39209 34731 39267 34737
rect 39209 34728 39221 34731
rect 38703 34700 39221 34728
rect 38703 34697 38715 34700
rect 38657 34691 38715 34697
rect 39209 34697 39221 34700
rect 39255 34728 39267 34731
rect 39666 34728 39672 34740
rect 39255 34700 39672 34728
rect 39255 34697 39267 34700
rect 39209 34691 39267 34697
rect 33042 34620 33048 34672
rect 33100 34660 33106 34672
rect 33381 34663 33439 34669
rect 33381 34660 33393 34663
rect 33100 34632 33393 34660
rect 33100 34620 33106 34632
rect 33381 34629 33393 34632
rect 33427 34629 33439 34663
rect 33381 34623 33439 34629
rect 33597 34663 33655 34669
rect 33597 34629 33609 34663
rect 33643 34660 33655 34663
rect 34330 34660 34336 34672
rect 33643 34632 34336 34660
rect 33643 34629 33655 34632
rect 33597 34623 33655 34629
rect 32493 34595 32551 34601
rect 32493 34561 32505 34595
rect 32539 34561 32551 34595
rect 32493 34555 32551 34561
rect 32508 34524 32536 34555
rect 32582 34552 32588 34604
rect 32640 34592 32646 34604
rect 32769 34595 32827 34601
rect 32640 34564 32685 34592
rect 32640 34552 32646 34564
rect 32769 34561 32781 34595
rect 32815 34561 32827 34595
rect 32769 34555 32827 34561
rect 30852 34496 32536 34524
rect 27338 34456 27344 34468
rect 24167 34428 25455 34456
rect 24167 34425 24179 34428
rect 24121 34419 24179 34425
rect 17402 34388 17408 34400
rect 17363 34360 17408 34388
rect 17402 34348 17408 34360
rect 17460 34348 17466 34400
rect 18049 34391 18107 34397
rect 18049 34357 18061 34391
rect 18095 34388 18107 34391
rect 18138 34388 18144 34400
rect 18095 34360 18144 34388
rect 18095 34357 18107 34360
rect 18049 34351 18107 34357
rect 18138 34348 18144 34360
rect 18196 34348 18202 34400
rect 22557 34391 22615 34397
rect 22557 34357 22569 34391
rect 22603 34388 22615 34391
rect 22646 34388 22652 34400
rect 22603 34360 22652 34388
rect 22603 34357 22615 34360
rect 22557 34351 22615 34357
rect 22646 34348 22652 34360
rect 22704 34348 22710 34400
rect 24670 34388 24676 34400
rect 24631 34360 24676 34388
rect 24670 34348 24676 34360
rect 24728 34348 24734 34400
rect 25427 34388 25455 34428
rect 25644 34428 27344 34456
rect 25644 34388 25672 34428
rect 27338 34416 27344 34428
rect 27396 34416 27402 34468
rect 28905 34459 28963 34465
rect 28905 34425 28917 34459
rect 28951 34456 28963 34459
rect 29822 34456 29828 34468
rect 28951 34428 29828 34456
rect 28951 34425 28963 34428
rect 28905 34419 28963 34425
rect 29822 34416 29828 34428
rect 29880 34416 29886 34468
rect 30098 34416 30104 34468
rect 30156 34456 30162 34468
rect 32784 34456 32812 34555
rect 32858 34552 32864 34604
rect 32916 34592 32922 34604
rect 33612 34592 33640 34623
rect 34330 34620 34336 34632
rect 34388 34620 34394 34672
rect 34606 34660 34612 34672
rect 34519 34632 34612 34660
rect 34532 34601 34560 34632
rect 34606 34620 34612 34632
rect 34664 34660 34670 34672
rect 35253 34663 35311 34669
rect 35253 34660 35265 34663
rect 34664 34632 35265 34660
rect 34664 34620 34670 34632
rect 35253 34629 35265 34632
rect 35299 34629 35311 34663
rect 35253 34623 35311 34629
rect 32916 34564 33640 34592
rect 34517 34595 34575 34601
rect 32916 34552 32922 34564
rect 34517 34561 34529 34595
rect 34563 34561 34575 34595
rect 34517 34555 34575 34561
rect 34790 34552 34796 34604
rect 34848 34592 34854 34604
rect 35161 34595 35219 34601
rect 35161 34592 35173 34595
rect 34848 34564 35173 34592
rect 34848 34552 34854 34564
rect 35161 34561 35173 34564
rect 35207 34561 35219 34595
rect 35342 34592 35348 34604
rect 35303 34564 35348 34592
rect 35161 34555 35219 34561
rect 35342 34552 35348 34564
rect 35400 34552 35406 34604
rect 35802 34592 35808 34604
rect 35763 34564 35808 34592
rect 35802 34552 35808 34564
rect 35860 34552 35866 34604
rect 35986 34592 35992 34604
rect 35947 34564 35992 34592
rect 35986 34552 35992 34564
rect 36044 34552 36050 34604
rect 36446 34552 36452 34604
rect 36504 34592 36510 34604
rect 37369 34595 37427 34601
rect 37369 34592 37381 34595
rect 36504 34564 37381 34592
rect 36504 34552 36510 34564
rect 37369 34561 37381 34564
rect 37415 34561 37427 34595
rect 37369 34555 37427 34561
rect 37553 34595 37611 34601
rect 37553 34561 37565 34595
rect 37599 34592 37611 34595
rect 37642 34592 37648 34604
rect 37599 34564 37648 34592
rect 37599 34561 37611 34564
rect 37553 34555 37611 34561
rect 37642 34552 37648 34564
rect 37700 34592 37706 34604
rect 38672 34592 38700 34691
rect 39666 34688 39672 34700
rect 39724 34688 39730 34740
rect 37700 34564 38700 34592
rect 37700 34552 37706 34564
rect 34609 34527 34667 34533
rect 34609 34493 34621 34527
rect 34655 34524 34667 34527
rect 34698 34524 34704 34536
rect 34655 34496 34704 34524
rect 34655 34493 34667 34496
rect 34609 34487 34667 34493
rect 34698 34484 34704 34496
rect 34756 34484 34762 34536
rect 38838 34524 38844 34536
rect 38626 34496 38844 34524
rect 30156 34428 32812 34456
rect 30156 34416 30162 34428
rect 25427 34360 25672 34388
rect 27157 34391 27215 34397
rect 27157 34357 27169 34391
rect 27203 34388 27215 34391
rect 27430 34388 27436 34400
rect 27203 34360 27436 34388
rect 27203 34357 27215 34360
rect 27157 34351 27215 34357
rect 27430 34348 27436 34360
rect 27488 34348 27494 34400
rect 28166 34388 28172 34400
rect 28127 34360 28172 34388
rect 28166 34348 28172 34360
rect 28224 34348 28230 34400
rect 31294 34348 31300 34400
rect 31352 34388 31358 34400
rect 32398 34388 32404 34400
rect 31352 34360 32404 34388
rect 31352 34348 31358 34360
rect 32398 34348 32404 34360
rect 32456 34348 32462 34400
rect 33226 34388 33232 34400
rect 33187 34360 33232 34388
rect 33226 34348 33232 34360
rect 33284 34348 33290 34400
rect 33410 34388 33416 34400
rect 33371 34360 33416 34388
rect 33410 34348 33416 34360
rect 33468 34348 33474 34400
rect 35894 34388 35900 34400
rect 35855 34360 35900 34388
rect 35894 34348 35900 34360
rect 35952 34348 35958 34400
rect 38010 34388 38016 34400
rect 37971 34360 38016 34388
rect 38010 34348 38016 34360
rect 38068 34388 38074 34400
rect 38626 34388 38654 34496
rect 38838 34484 38844 34496
rect 38896 34484 38902 34536
rect 39666 34484 39672 34536
rect 39724 34524 39730 34536
rect 50706 34524 50712 34536
rect 39724 34496 50712 34524
rect 39724 34484 39730 34496
rect 50706 34484 50712 34496
rect 50764 34484 50770 34536
rect 38068 34360 38654 34388
rect 38068 34348 38074 34360
rect 1104 34298 54372 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 54372 34298
rect 1104 34224 54372 34246
rect 16850 34144 16856 34196
rect 16908 34184 16914 34196
rect 17405 34187 17463 34193
rect 17405 34184 17417 34187
rect 16908 34156 17417 34184
rect 16908 34144 16914 34156
rect 17405 34153 17417 34156
rect 17451 34153 17463 34187
rect 17405 34147 17463 34153
rect 17957 34187 18015 34193
rect 17957 34153 17969 34187
rect 18003 34184 18015 34187
rect 18046 34184 18052 34196
rect 18003 34156 18052 34184
rect 18003 34153 18015 34156
rect 17957 34147 18015 34153
rect 1578 34116 1584 34128
rect 1539 34088 1584 34116
rect 1578 34076 1584 34088
rect 1636 34076 1642 34128
rect 17420 34116 17448 34147
rect 18046 34144 18052 34156
rect 18104 34144 18110 34196
rect 19426 34184 19432 34196
rect 18340 34156 19432 34184
rect 18340 34116 18368 34156
rect 19426 34144 19432 34156
rect 19484 34144 19490 34196
rect 19794 34144 19800 34196
rect 19852 34184 19858 34196
rect 19889 34187 19947 34193
rect 19889 34184 19901 34187
rect 19852 34156 19901 34184
rect 19852 34144 19858 34156
rect 19889 34153 19901 34156
rect 19935 34153 19947 34187
rect 19889 34147 19947 34153
rect 19981 34187 20039 34193
rect 19981 34153 19993 34187
rect 20027 34184 20039 34187
rect 20806 34184 20812 34196
rect 20027 34156 20812 34184
rect 20027 34153 20039 34156
rect 19981 34147 20039 34153
rect 20806 34144 20812 34156
rect 20864 34144 20870 34196
rect 25498 34184 25504 34196
rect 25459 34156 25504 34184
rect 25498 34144 25504 34156
rect 25556 34144 25562 34196
rect 26050 34184 26056 34196
rect 26011 34156 26056 34184
rect 26050 34144 26056 34156
rect 26108 34144 26114 34196
rect 26234 34184 26240 34196
rect 26195 34156 26240 34184
rect 26234 34144 26240 34156
rect 26292 34144 26298 34196
rect 26878 34184 26884 34196
rect 26839 34156 26884 34184
rect 26878 34144 26884 34156
rect 26936 34144 26942 34196
rect 27801 34187 27859 34193
rect 27801 34153 27813 34187
rect 27847 34184 27859 34187
rect 29914 34184 29920 34196
rect 27847 34156 29920 34184
rect 27847 34153 27859 34156
rect 27801 34147 27859 34153
rect 29914 34144 29920 34156
rect 29972 34144 29978 34196
rect 32493 34187 32551 34193
rect 32493 34153 32505 34187
rect 32539 34184 32551 34187
rect 32582 34184 32588 34196
rect 32539 34156 32588 34184
rect 32539 34153 32551 34156
rect 32493 34147 32551 34153
rect 32582 34144 32588 34156
rect 32640 34144 32646 34196
rect 32674 34144 32680 34196
rect 32732 34184 32738 34196
rect 35342 34184 35348 34196
rect 32732 34156 32777 34184
rect 33888 34156 35348 34184
rect 32732 34144 32738 34156
rect 17420 34088 18368 34116
rect 18414 34076 18420 34128
rect 18472 34116 18478 34128
rect 19337 34119 19395 34125
rect 19337 34116 19349 34119
rect 18472 34088 19349 34116
rect 18472 34076 18478 34088
rect 19337 34085 19349 34088
rect 19383 34116 19395 34119
rect 22186 34116 22192 34128
rect 19383 34088 22192 34116
rect 19383 34085 19395 34088
rect 19337 34079 19395 34085
rect 22186 34076 22192 34088
rect 22244 34076 22250 34128
rect 23845 34119 23903 34125
rect 23845 34085 23857 34119
rect 23891 34116 23903 34119
rect 24854 34116 24860 34128
rect 23891 34088 24860 34116
rect 23891 34085 23903 34088
rect 23845 34079 23903 34085
rect 24854 34076 24860 34088
rect 24912 34076 24918 34128
rect 26418 34116 26424 34128
rect 25240 34088 26424 34116
rect 16393 34051 16451 34057
rect 16393 34017 16405 34051
rect 16439 34048 16451 34051
rect 18230 34048 18236 34060
rect 16439 34020 18236 34048
rect 16439 34017 16451 34020
rect 16393 34011 16451 34017
rect 18230 34008 18236 34020
rect 18288 34008 18294 34060
rect 20070 34048 20076 34060
rect 20031 34020 20076 34048
rect 20070 34008 20076 34020
rect 20128 34008 20134 34060
rect 22097 34051 22155 34057
rect 22097 34017 22109 34051
rect 22143 34048 22155 34051
rect 23566 34048 23572 34060
rect 22143 34020 22876 34048
rect 23527 34020 23572 34048
rect 22143 34017 22155 34020
rect 22097 34011 22155 34017
rect 18138 33980 18144 33992
rect 18099 33952 18144 33980
rect 18138 33940 18144 33952
rect 18196 33940 18202 33992
rect 19426 33940 19432 33992
rect 19484 33980 19490 33992
rect 19797 33983 19855 33989
rect 19797 33980 19809 33983
rect 19484 33952 19809 33980
rect 19484 33940 19490 33952
rect 19797 33949 19809 33952
rect 19843 33980 19855 33983
rect 20901 33983 20959 33989
rect 20901 33980 20913 33983
rect 19843 33952 20913 33980
rect 19843 33949 19855 33952
rect 19797 33943 19855 33949
rect 20901 33949 20913 33952
rect 20947 33980 20959 33983
rect 22002 33980 22008 33992
rect 20947 33952 22008 33980
rect 20947 33949 20959 33952
rect 20901 33943 20959 33949
rect 22002 33940 22008 33952
rect 22060 33940 22066 33992
rect 22186 33980 22192 33992
rect 22147 33952 22192 33980
rect 22186 33940 22192 33952
rect 22244 33940 22250 33992
rect 22646 33980 22652 33992
rect 22607 33952 22652 33980
rect 22646 33940 22652 33952
rect 22704 33940 22710 33992
rect 22848 33989 22876 34020
rect 23566 34008 23572 34020
rect 23624 34008 23630 34060
rect 24670 34008 24676 34060
rect 24728 34048 24734 34060
rect 25240 34048 25268 34088
rect 26418 34076 26424 34088
rect 26476 34076 26482 34128
rect 28810 34116 28816 34128
rect 27632 34088 28816 34116
rect 24728 34020 25268 34048
rect 24728 34008 24734 34020
rect 22833 33983 22891 33989
rect 22833 33949 22845 33983
rect 22879 33980 22891 33983
rect 23290 33980 23296 33992
rect 22879 33952 23296 33980
rect 22879 33949 22891 33952
rect 22833 33943 22891 33949
rect 23290 33940 23296 33952
rect 23348 33940 23354 33992
rect 23477 33983 23535 33989
rect 23477 33949 23489 33983
rect 23523 33980 23535 33983
rect 23750 33980 23756 33992
rect 23523 33952 23756 33980
rect 23523 33949 23535 33952
rect 23477 33943 23535 33949
rect 18322 33912 18328 33924
rect 18283 33884 18328 33912
rect 18322 33872 18328 33884
rect 18380 33872 18386 33924
rect 22741 33915 22799 33921
rect 22741 33881 22753 33915
rect 22787 33912 22799 33915
rect 23492 33912 23520 33943
rect 23750 33940 23756 33952
rect 23808 33940 23814 33992
rect 25240 33989 25268 34020
rect 25317 34051 25375 34057
rect 25317 34017 25329 34051
rect 25363 34048 25375 34051
rect 25363 34020 27108 34048
rect 25363 34017 25375 34020
rect 25317 34011 25375 34017
rect 25225 33983 25283 33989
rect 25225 33949 25237 33983
rect 25271 33949 25283 33983
rect 25225 33943 25283 33949
rect 22787 33884 23520 33912
rect 22787 33881 22799 33884
rect 22741 33875 22799 33881
rect 16758 33804 16764 33856
rect 16816 33844 16822 33856
rect 16853 33847 16911 33853
rect 16853 33844 16865 33847
rect 16816 33816 16865 33844
rect 16816 33804 16822 33816
rect 16853 33813 16865 33816
rect 16899 33813 16911 33847
rect 21450 33844 21456 33856
rect 21411 33816 21456 33844
rect 16853 33807 16911 33813
rect 21450 33804 21456 33816
rect 21508 33804 21514 33856
rect 24486 33844 24492 33856
rect 24447 33816 24492 33844
rect 24486 33804 24492 33816
rect 24544 33804 24550 33856
rect 26160 33844 26188 34020
rect 27080 33992 27108 34020
rect 26234 33940 26240 33992
rect 26292 33982 26298 33992
rect 26881 33983 26939 33989
rect 26292 33980 26326 33982
rect 26881 33980 26893 33983
rect 26292 33952 26893 33980
rect 26292 33940 26298 33952
rect 26881 33949 26893 33952
rect 26927 33949 26939 33983
rect 26881 33943 26939 33949
rect 27062 33940 27068 33992
rect 27120 33980 27126 33992
rect 27632 33989 27660 34088
rect 28810 34076 28816 34088
rect 28868 34076 28874 34128
rect 28905 34119 28963 34125
rect 28905 34085 28917 34119
rect 28951 34116 28963 34119
rect 28994 34116 29000 34128
rect 28951 34088 29000 34116
rect 28951 34085 28963 34088
rect 28905 34079 28963 34085
rect 28994 34076 29000 34088
rect 29052 34076 29058 34128
rect 29270 34076 29276 34128
rect 29328 34116 29334 34128
rect 29730 34116 29736 34128
rect 29328 34088 29736 34116
rect 29328 34076 29334 34088
rect 29730 34076 29736 34088
rect 29788 34116 29794 34128
rect 29788 34088 31248 34116
rect 29788 34076 29794 34088
rect 27893 34051 27951 34057
rect 27893 34017 27905 34051
rect 27939 34048 27951 34051
rect 28258 34048 28264 34060
rect 27939 34020 28264 34048
rect 27939 34017 27951 34020
rect 27893 34011 27951 34017
rect 28258 34008 28264 34020
rect 28316 34008 28322 34060
rect 28350 34008 28356 34060
rect 28408 34048 28414 34060
rect 28445 34051 28503 34057
rect 28445 34048 28457 34051
rect 28408 34020 28457 34048
rect 28408 34008 28414 34020
rect 28445 34017 28457 34020
rect 28491 34017 28503 34051
rect 29086 34048 29092 34060
rect 28445 34011 28503 34017
rect 28644 34020 29092 34048
rect 27157 33983 27215 33989
rect 27157 33980 27169 33983
rect 27120 33952 27169 33980
rect 27120 33940 27126 33952
rect 27157 33949 27169 33952
rect 27203 33949 27215 33983
rect 27157 33943 27215 33949
rect 27617 33983 27675 33989
rect 27617 33949 27629 33983
rect 27663 33949 27675 33983
rect 27617 33943 27675 33949
rect 27709 33983 27767 33989
rect 27709 33949 27721 33983
rect 27755 33949 27767 33983
rect 27709 33943 27767 33949
rect 26418 33912 26424 33924
rect 26379 33884 26424 33912
rect 26418 33872 26424 33884
rect 26476 33872 26482 33924
rect 27724 33912 27752 33943
rect 28166 33940 28172 33992
rect 28224 33980 28230 33992
rect 28537 33983 28595 33989
rect 28537 33980 28549 33983
rect 28224 33952 28549 33980
rect 28224 33940 28230 33952
rect 28537 33949 28549 33952
rect 28583 33980 28595 33983
rect 28644 33980 28672 34020
rect 29086 34008 29092 34020
rect 29144 34048 29150 34060
rect 29546 34048 29552 34060
rect 29144 34020 29552 34048
rect 29144 34008 29150 34020
rect 29546 34008 29552 34020
rect 29604 34008 29610 34060
rect 29822 34048 29828 34060
rect 29735 34020 29828 34048
rect 29822 34008 29828 34020
rect 29880 34048 29886 34060
rect 31220 34057 31248 34088
rect 31205 34051 31263 34057
rect 29880 34020 30972 34048
rect 29880 34008 29886 34020
rect 28583 33952 28672 33980
rect 28583 33949 28595 33952
rect 28537 33943 28595 33949
rect 28810 33940 28816 33992
rect 28868 33980 28874 33992
rect 29730 33980 29736 33992
rect 28868 33952 29736 33980
rect 28868 33940 28874 33952
rect 29730 33940 29736 33952
rect 29788 33940 29794 33992
rect 29840 33912 29868 34008
rect 30098 33940 30104 33992
rect 30156 33980 30162 33992
rect 30837 33983 30895 33989
rect 30837 33980 30849 33983
rect 30156 33952 30849 33980
rect 30156 33940 30162 33952
rect 30837 33949 30849 33952
rect 30883 33949 30895 33983
rect 30837 33943 30895 33949
rect 30116 33912 30144 33940
rect 27724 33884 29868 33912
rect 29932 33884 30144 33912
rect 30944 33912 30972 34020
rect 31205 34017 31217 34051
rect 31251 34017 31263 34051
rect 31205 34011 31263 34017
rect 31386 34008 31392 34060
rect 31444 34048 31450 34060
rect 31444 34020 32904 34048
rect 31444 34008 31450 34020
rect 31294 33940 31300 33992
rect 31352 33980 31358 33992
rect 32766 33980 32772 33992
rect 31352 33952 31397 33980
rect 32727 33952 32772 33980
rect 31352 33940 31358 33952
rect 32766 33940 32772 33952
rect 32824 33940 32830 33992
rect 32876 33989 32904 34020
rect 32861 33983 32919 33989
rect 32861 33949 32873 33983
rect 32907 33980 32919 33983
rect 33226 33980 33232 33992
rect 32907 33952 33232 33980
rect 32907 33949 32919 33952
rect 32861 33943 32919 33949
rect 33226 33940 33232 33952
rect 33284 33940 33290 33992
rect 33888 33989 33916 34156
rect 35342 34144 35348 34156
rect 35400 34144 35406 34196
rect 35897 34187 35955 34193
rect 35897 34153 35909 34187
rect 35943 34184 35955 34187
rect 36538 34184 36544 34196
rect 35943 34156 36544 34184
rect 35943 34153 35955 34156
rect 35897 34147 35955 34153
rect 36538 34144 36544 34156
rect 36596 34144 36602 34196
rect 34057 34119 34115 34125
rect 34057 34085 34069 34119
rect 34103 34116 34115 34119
rect 34698 34116 34704 34128
rect 34103 34088 34704 34116
rect 34103 34085 34115 34088
rect 34057 34079 34115 34085
rect 34698 34076 34704 34088
rect 34756 34116 34762 34128
rect 34977 34119 35035 34125
rect 34977 34116 34989 34119
rect 34756 34088 34989 34116
rect 34756 34076 34762 34088
rect 34977 34085 34989 34088
rect 35023 34085 35035 34119
rect 34977 34079 35035 34085
rect 35069 34051 35127 34057
rect 35069 34017 35081 34051
rect 35115 34048 35127 34051
rect 35894 34048 35900 34060
rect 35115 34020 35900 34048
rect 35115 34017 35127 34020
rect 35069 34011 35127 34017
rect 35894 34008 35900 34020
rect 35952 34008 35958 34060
rect 33873 33983 33931 33989
rect 33873 33949 33885 33983
rect 33919 33949 33931 33983
rect 33873 33943 33931 33949
rect 34149 33983 34207 33989
rect 34149 33949 34161 33983
rect 34195 33980 34207 33983
rect 34606 33980 34612 33992
rect 34195 33952 34612 33980
rect 34195 33949 34207 33952
rect 34149 33943 34207 33949
rect 34606 33940 34612 33952
rect 34664 33980 34670 33992
rect 34885 33983 34943 33989
rect 34885 33980 34897 33983
rect 34664 33952 34897 33980
rect 34664 33940 34670 33952
rect 34885 33949 34897 33952
rect 34931 33949 34943 33983
rect 34885 33943 34943 33949
rect 35161 33983 35219 33989
rect 35161 33949 35173 33983
rect 35207 33980 35219 33983
rect 35342 33980 35348 33992
rect 35207 33952 35348 33980
rect 35207 33949 35219 33952
rect 35161 33943 35219 33949
rect 35342 33940 35348 33952
rect 35400 33940 35406 33992
rect 35526 33940 35532 33992
rect 35584 33980 35590 33992
rect 38841 33983 38899 33989
rect 35584 33952 36124 33980
rect 35584 33940 35590 33952
rect 34701 33915 34759 33921
rect 34701 33912 34713 33915
rect 30944 33884 34713 33912
rect 26216 33847 26274 33853
rect 26216 33844 26228 33847
rect 26160 33816 26228 33844
rect 26216 33813 26228 33816
rect 26262 33813 26274 33847
rect 26216 33807 26274 33813
rect 27065 33847 27123 33853
rect 27065 33813 27077 33847
rect 27111 33844 27123 33847
rect 27154 33844 27160 33856
rect 27111 33816 27160 33844
rect 27111 33813 27123 33816
rect 27065 33807 27123 33813
rect 27154 33804 27160 33816
rect 27212 33804 27218 33856
rect 27246 33804 27252 33856
rect 27304 33844 27310 33856
rect 29932 33844 29960 33884
rect 34701 33881 34713 33884
rect 34747 33881 34759 33915
rect 34701 33875 34759 33881
rect 35881 33915 35939 33921
rect 35881 33881 35893 33915
rect 35927 33912 35939 33915
rect 35986 33912 35992 33924
rect 35927 33884 35992 33912
rect 35927 33881 35939 33884
rect 35881 33875 35939 33881
rect 35986 33872 35992 33884
rect 36044 33872 36050 33924
rect 36096 33921 36124 33952
rect 38841 33949 38853 33983
rect 38887 33980 38899 33983
rect 38930 33980 38936 33992
rect 38887 33952 38936 33980
rect 38887 33949 38899 33952
rect 38841 33943 38899 33949
rect 38930 33940 38936 33952
rect 38988 33980 38994 33992
rect 53650 33980 53656 33992
rect 38988 33952 53656 33980
rect 38988 33940 38994 33952
rect 53650 33940 53656 33952
rect 53708 33940 53714 33992
rect 36081 33915 36139 33921
rect 36081 33881 36093 33915
rect 36127 33912 36139 33915
rect 37093 33915 37151 33921
rect 37093 33912 37105 33915
rect 36127 33884 37105 33912
rect 36127 33881 36139 33884
rect 36081 33875 36139 33881
rect 37093 33881 37105 33884
rect 37139 33912 37151 33915
rect 38010 33912 38016 33924
rect 37139 33884 38016 33912
rect 37139 33881 37151 33884
rect 37093 33875 37151 33881
rect 38010 33872 38016 33884
rect 38068 33872 38074 33924
rect 27304 33816 29960 33844
rect 30101 33847 30159 33853
rect 27304 33804 27310 33816
rect 30101 33813 30113 33847
rect 30147 33844 30159 33847
rect 30374 33844 30380 33856
rect 30147 33816 30380 33844
rect 30147 33813 30159 33816
rect 30101 33807 30159 33813
rect 30374 33804 30380 33816
rect 30432 33804 30438 33856
rect 30466 33804 30472 33856
rect 30524 33844 30530 33856
rect 31570 33844 31576 33856
rect 30524 33816 31576 33844
rect 30524 33804 30530 33816
rect 31570 33804 31576 33816
rect 31628 33804 31634 33856
rect 32582 33804 32588 33856
rect 32640 33844 32646 33856
rect 32858 33844 32864 33856
rect 32640 33816 32864 33844
rect 32640 33804 32646 33816
rect 32858 33804 32864 33816
rect 32916 33804 32922 33856
rect 33689 33847 33747 33853
rect 33689 33813 33701 33847
rect 33735 33844 33747 33847
rect 34330 33844 34336 33856
rect 33735 33816 34336 33844
rect 33735 33813 33747 33816
rect 33689 33807 33747 33813
rect 34330 33804 34336 33816
rect 34388 33804 34394 33856
rect 35710 33844 35716 33856
rect 35671 33816 35716 33844
rect 35710 33804 35716 33816
rect 35768 33804 35774 33856
rect 37642 33844 37648 33856
rect 37603 33816 37648 33844
rect 37642 33804 37648 33816
rect 37700 33804 37706 33856
rect 38194 33844 38200 33856
rect 38155 33816 38200 33844
rect 38194 33804 38200 33816
rect 38252 33804 38258 33856
rect 39945 33847 40003 33853
rect 39945 33813 39957 33847
rect 39991 33844 40003 33847
rect 40402 33844 40408 33856
rect 39991 33816 40408 33844
rect 39991 33813 40003 33816
rect 39945 33807 40003 33813
rect 40402 33804 40408 33816
rect 40460 33804 40466 33856
rect 1104 33754 54372 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 54372 33754
rect 1104 33680 54372 33702
rect 18049 33643 18107 33649
rect 18049 33609 18061 33643
rect 18095 33640 18107 33643
rect 18322 33640 18328 33652
rect 18095 33612 18328 33640
rect 18095 33609 18107 33612
rect 18049 33603 18107 33609
rect 18322 33600 18328 33612
rect 18380 33600 18386 33652
rect 18966 33640 18972 33652
rect 18927 33612 18972 33640
rect 18966 33600 18972 33612
rect 19024 33600 19030 33652
rect 24670 33640 24676 33652
rect 24631 33612 24676 33640
rect 24670 33600 24676 33612
rect 24728 33600 24734 33652
rect 26421 33643 26479 33649
rect 26421 33609 26433 33643
rect 26467 33640 26479 33643
rect 26510 33640 26516 33652
rect 26467 33612 26516 33640
rect 26467 33609 26479 33612
rect 26421 33603 26479 33609
rect 26510 33600 26516 33612
rect 26568 33600 26574 33652
rect 29270 33640 29276 33652
rect 27540 33612 29276 33640
rect 17497 33575 17555 33581
rect 17497 33541 17509 33575
rect 17543 33572 17555 33575
rect 17543 33544 18184 33572
rect 17543 33541 17555 33544
rect 17497 33535 17555 33541
rect 16390 33464 16396 33516
rect 16448 33504 16454 33516
rect 18156 33513 18184 33544
rect 21910 33532 21916 33584
rect 21968 33572 21974 33584
rect 24029 33575 24087 33581
rect 24029 33572 24041 33575
rect 21968 33544 24041 33572
rect 21968 33532 21974 33544
rect 24029 33541 24041 33544
rect 24075 33572 24087 33575
rect 24486 33572 24492 33584
rect 24075 33544 24492 33572
rect 24075 33541 24087 33544
rect 24029 33535 24087 33541
rect 24486 33532 24492 33544
rect 24544 33572 24550 33584
rect 25225 33575 25283 33581
rect 25225 33572 25237 33575
rect 24544 33544 25237 33572
rect 24544 33532 24550 33544
rect 25225 33541 25237 33544
rect 25271 33572 25283 33575
rect 26234 33572 26240 33584
rect 25271 33544 26240 33572
rect 25271 33541 25283 33544
rect 25225 33535 25283 33541
rect 26234 33532 26240 33544
rect 26292 33532 26298 33584
rect 16945 33507 17003 33513
rect 16945 33504 16957 33507
rect 16448 33476 16957 33504
rect 16448 33464 16454 33476
rect 16945 33473 16957 33476
rect 16991 33504 17003 33507
rect 17957 33507 18015 33513
rect 17957 33504 17969 33507
rect 16991 33476 17969 33504
rect 16991 33473 17003 33476
rect 16945 33467 17003 33473
rect 17957 33473 17969 33476
rect 18003 33473 18015 33507
rect 17957 33467 18015 33473
rect 18141 33507 18199 33513
rect 18141 33473 18153 33507
rect 18187 33504 18199 33507
rect 18230 33504 18236 33516
rect 18187 33476 18236 33504
rect 18187 33473 18199 33476
rect 18141 33467 18199 33473
rect 18230 33464 18236 33476
rect 18288 33464 18294 33516
rect 22465 33507 22523 33513
rect 22465 33473 22477 33507
rect 22511 33504 22523 33507
rect 22554 33504 22560 33516
rect 22511 33476 22560 33504
rect 22511 33473 22523 33476
rect 22465 33467 22523 33473
rect 22554 33464 22560 33476
rect 22612 33464 22618 33516
rect 22646 33464 22652 33516
rect 22704 33504 22710 33516
rect 23290 33504 23296 33516
rect 22704 33476 22749 33504
rect 23251 33476 23296 33504
rect 22704 33464 22710 33476
rect 23290 33464 23296 33476
rect 23348 33464 23354 33516
rect 23382 33464 23388 33516
rect 23440 33504 23446 33516
rect 27157 33507 27215 33513
rect 27157 33504 27169 33507
rect 23440 33476 27169 33504
rect 23440 33464 23446 33476
rect 27157 33473 27169 33476
rect 27203 33473 27215 33507
rect 27157 33467 27215 33473
rect 27246 33464 27252 33516
rect 27304 33504 27310 33516
rect 27540 33513 27568 33612
rect 29270 33600 29276 33612
rect 29328 33600 29334 33652
rect 29365 33643 29423 33649
rect 29365 33609 29377 33643
rect 29411 33640 29423 33643
rect 29638 33640 29644 33652
rect 29411 33612 29644 33640
rect 29411 33609 29423 33612
rect 29365 33603 29423 33609
rect 29638 33600 29644 33612
rect 29696 33600 29702 33652
rect 29730 33600 29736 33652
rect 29788 33640 29794 33652
rect 31297 33643 31355 33649
rect 31297 33640 31309 33643
rect 29788 33612 31309 33640
rect 29788 33600 29794 33612
rect 31297 33609 31309 33612
rect 31343 33609 31355 33643
rect 31297 33603 31355 33609
rect 32674 33600 32680 33652
rect 32732 33640 32738 33652
rect 32854 33643 32912 33649
rect 32854 33640 32866 33643
rect 32732 33612 32866 33640
rect 32732 33600 32738 33612
rect 32854 33609 32866 33612
rect 32900 33609 32912 33643
rect 32854 33603 32912 33609
rect 33318 33600 33324 33652
rect 33376 33640 33382 33652
rect 33505 33643 33563 33649
rect 33505 33640 33517 33643
rect 33376 33612 33517 33640
rect 33376 33600 33382 33612
rect 33505 33609 33517 33612
rect 33551 33640 33563 33643
rect 34698 33640 34704 33652
rect 33551 33612 34704 33640
rect 33551 33609 33563 33612
rect 33505 33603 33563 33609
rect 34698 33600 34704 33612
rect 34756 33600 34762 33652
rect 34790 33600 34796 33652
rect 34848 33640 34854 33652
rect 35069 33643 35127 33649
rect 35069 33640 35081 33643
rect 34848 33612 35081 33640
rect 34848 33600 34854 33612
rect 35069 33609 35081 33612
rect 35115 33609 35127 33643
rect 35069 33603 35127 33609
rect 35250 33600 35256 33652
rect 35308 33640 35314 33652
rect 35526 33640 35532 33652
rect 35308 33612 35532 33640
rect 35308 33600 35314 33612
rect 35526 33600 35532 33612
rect 35584 33600 35590 33652
rect 35897 33643 35955 33649
rect 35897 33609 35909 33643
rect 35943 33640 35955 33643
rect 35986 33640 35992 33652
rect 35943 33612 35992 33640
rect 35943 33609 35955 33612
rect 35897 33603 35955 33609
rect 35986 33600 35992 33612
rect 36044 33600 36050 33652
rect 28258 33532 28264 33584
rect 28316 33572 28322 33584
rect 30466 33572 30472 33584
rect 28316 33544 30144 33572
rect 30427 33544 30472 33572
rect 28316 33532 28322 33544
rect 27525 33507 27583 33513
rect 27304 33476 27349 33504
rect 27304 33464 27310 33476
rect 27525 33473 27537 33507
rect 27571 33473 27583 33507
rect 27525 33467 27583 33473
rect 28077 33507 28135 33513
rect 28077 33473 28089 33507
rect 28123 33504 28135 33507
rect 28537 33507 28595 33513
rect 28537 33504 28549 33507
rect 28123 33476 28549 33504
rect 28123 33473 28135 33476
rect 28077 33467 28135 33473
rect 28537 33473 28549 33476
rect 28583 33504 28595 33507
rect 28583 33476 28672 33504
rect 28583 33473 28595 33476
rect 28537 33467 28595 33473
rect 20073 33439 20131 33445
rect 20073 33405 20085 33439
rect 20119 33436 20131 33439
rect 21266 33436 21272 33448
rect 20119 33408 21272 33436
rect 20119 33405 20131 33408
rect 20073 33399 20131 33405
rect 21266 33396 21272 33408
rect 21324 33436 21330 33448
rect 21821 33439 21879 33445
rect 21821 33436 21833 33439
rect 21324 33408 21833 33436
rect 21324 33396 21330 33408
rect 21821 33405 21833 33408
rect 21867 33405 21879 33439
rect 21821 33399 21879 33405
rect 23569 33439 23627 33445
rect 23569 33405 23581 33439
rect 23615 33436 23627 33439
rect 23750 33436 23756 33448
rect 23615 33408 23756 33436
rect 23615 33405 23627 33408
rect 23569 33399 23627 33405
rect 23750 33396 23756 33408
rect 23808 33396 23814 33448
rect 27430 33436 27436 33448
rect 27391 33408 27436 33436
rect 27430 33396 27436 33408
rect 27488 33396 27494 33448
rect 20717 33371 20775 33377
rect 20717 33337 20729 33371
rect 20763 33368 20775 33371
rect 21358 33368 21364 33380
rect 20763 33340 21364 33368
rect 20763 33337 20775 33340
rect 20717 33331 20775 33337
rect 21358 33328 21364 33340
rect 21416 33328 21422 33380
rect 22557 33371 22615 33377
rect 22557 33337 22569 33371
rect 22603 33368 22615 33371
rect 24486 33368 24492 33380
rect 22603 33340 24492 33368
rect 22603 33337 22615 33340
rect 22557 33331 22615 33337
rect 24486 33328 24492 33340
rect 24544 33328 24550 33380
rect 19334 33260 19340 33312
rect 19392 33300 19398 33312
rect 19429 33303 19487 33309
rect 19429 33300 19441 33303
rect 19392 33272 19441 33300
rect 19392 33260 19398 33272
rect 19429 33269 19441 33272
rect 19475 33269 19487 33303
rect 19429 33263 19487 33269
rect 20806 33260 20812 33312
rect 20864 33300 20870 33312
rect 21177 33303 21235 33309
rect 21177 33300 21189 33303
rect 20864 33272 21189 33300
rect 20864 33260 20870 33272
rect 21177 33269 21189 33272
rect 21223 33300 21235 33303
rect 21450 33300 21456 33312
rect 21223 33272 21456 33300
rect 21223 33269 21235 33272
rect 21177 33263 21235 33269
rect 21450 33260 21456 33272
rect 21508 33260 21514 33312
rect 23106 33300 23112 33312
rect 23067 33272 23112 33300
rect 23106 33260 23112 33272
rect 23164 33260 23170 33312
rect 23477 33303 23535 33309
rect 23477 33269 23489 33303
rect 23523 33300 23535 33303
rect 23566 33300 23572 33312
rect 23523 33272 23572 33300
rect 23523 33269 23535 33272
rect 23477 33263 23535 33269
rect 23566 33260 23572 33272
rect 23624 33300 23630 33312
rect 23842 33300 23848 33312
rect 23624 33272 23848 33300
rect 23624 33260 23630 33272
rect 23842 33260 23848 33272
rect 23900 33260 23906 33312
rect 25774 33300 25780 33312
rect 25735 33272 25780 33300
rect 25774 33260 25780 33272
rect 25832 33260 25838 33312
rect 26418 33260 26424 33312
rect 26476 33300 26482 33312
rect 26973 33303 27031 33309
rect 26973 33300 26985 33303
rect 26476 33272 26985 33300
rect 26476 33260 26482 33272
rect 26973 33269 26985 33272
rect 27019 33269 27031 33303
rect 28644 33300 28672 33476
rect 28718 33464 28724 33516
rect 28776 33504 28782 33516
rect 28776 33476 28821 33504
rect 28776 33464 28782 33476
rect 29086 33464 29092 33516
rect 29144 33504 29150 33516
rect 29595 33507 29653 33513
rect 29595 33504 29607 33507
rect 29144 33476 29607 33504
rect 29144 33464 29150 33476
rect 29595 33473 29607 33476
rect 29641 33473 29653 33507
rect 29595 33467 29653 33473
rect 29730 33507 29788 33513
rect 29730 33473 29742 33507
rect 29776 33473 29788 33507
rect 29730 33467 29788 33473
rect 29825 33507 29883 33513
rect 29825 33473 29837 33507
rect 29871 33504 29883 33507
rect 29914 33504 29920 33516
rect 29871 33476 29920 33504
rect 29871 33473 29883 33476
rect 29825 33467 29883 33473
rect 28905 33439 28963 33445
rect 28905 33405 28917 33439
rect 28951 33436 28963 33439
rect 29362 33436 29368 33448
rect 28951 33408 29368 33436
rect 28951 33405 28963 33408
rect 28905 33399 28963 33405
rect 29362 33396 29368 33408
rect 29420 33396 29426 33448
rect 28994 33328 29000 33380
rect 29052 33368 29058 33380
rect 29178 33368 29184 33380
rect 29052 33340 29184 33368
rect 29052 33328 29058 33340
rect 29178 33328 29184 33340
rect 29236 33368 29242 33380
rect 29748 33368 29776 33467
rect 29914 33464 29920 33476
rect 29972 33464 29978 33516
rect 30009 33507 30067 33513
rect 30009 33473 30021 33507
rect 30055 33473 30067 33507
rect 30116 33504 30144 33544
rect 30466 33532 30472 33544
rect 30524 33532 30530 33584
rect 30685 33575 30743 33581
rect 30685 33541 30697 33575
rect 30731 33572 30743 33575
rect 31386 33572 31392 33584
rect 30731 33544 31392 33572
rect 30731 33541 30743 33544
rect 30685 33535 30743 33541
rect 31386 33532 31392 33544
rect 31444 33532 31450 33584
rect 33042 33572 33048 33584
rect 32692 33544 33048 33572
rect 32692 33513 32720 33544
rect 33042 33532 33048 33544
rect 33100 33532 33106 33584
rect 34514 33532 34520 33584
rect 34572 33572 34578 33584
rect 35618 33572 35624 33584
rect 34572 33544 35624 33572
rect 34572 33532 34578 33544
rect 35618 33532 35624 33544
rect 35676 33532 35682 33584
rect 36538 33572 36544 33584
rect 35912 33544 36544 33572
rect 31297 33507 31355 33513
rect 31297 33504 31309 33507
rect 30116 33476 31309 33504
rect 30009 33467 30067 33473
rect 31297 33473 31309 33476
rect 31343 33473 31355 33507
rect 31297 33467 31355 33473
rect 31481 33507 31539 33513
rect 31481 33473 31493 33507
rect 31527 33473 31539 33507
rect 31481 33467 31539 33473
rect 32677 33507 32735 33513
rect 32677 33473 32689 33507
rect 32723 33473 32735 33507
rect 32677 33467 32735 33473
rect 32769 33507 32827 33513
rect 32769 33473 32781 33507
rect 32815 33473 32827 33507
rect 32769 33467 32827 33473
rect 32953 33507 33011 33513
rect 32953 33473 32965 33507
rect 32999 33504 33011 33507
rect 33410 33504 33416 33516
rect 32999 33476 33416 33504
rect 32999 33473 33011 33476
rect 32953 33467 33011 33473
rect 30024 33436 30052 33467
rect 29932 33408 30052 33436
rect 29932 33380 29960 33408
rect 30098 33396 30104 33448
rect 30156 33436 30162 33448
rect 31496 33436 31524 33467
rect 30156 33408 31524 33436
rect 32217 33439 32275 33445
rect 30156 33396 30162 33408
rect 32217 33405 32229 33439
rect 32263 33436 32275 33439
rect 32490 33436 32496 33448
rect 32263 33408 32496 33436
rect 32263 33405 32275 33408
rect 32217 33399 32275 33405
rect 32490 33396 32496 33408
rect 32548 33396 32554 33448
rect 32582 33396 32588 33448
rect 32640 33436 32646 33448
rect 32784 33436 32812 33467
rect 33410 33464 33416 33476
rect 33468 33464 33474 33516
rect 34425 33507 34483 33513
rect 34425 33473 34437 33507
rect 34471 33473 34483 33507
rect 35250 33504 35256 33516
rect 35211 33476 35256 33504
rect 34425 33467 34483 33473
rect 32640 33408 32812 33436
rect 32640 33396 32646 33408
rect 32858 33396 32864 33448
rect 32916 33436 32922 33448
rect 34330 33436 34336 33448
rect 32916 33408 34192 33436
rect 34291 33408 34336 33436
rect 32916 33396 32922 33408
rect 29914 33368 29920 33380
rect 29236 33340 29776 33368
rect 29827 33340 29920 33368
rect 29236 33328 29242 33340
rect 29914 33328 29920 33340
rect 29972 33368 29978 33380
rect 33318 33368 33324 33380
rect 29972 33340 33324 33368
rect 29972 33328 29978 33340
rect 29932 33300 29960 33328
rect 30668 33309 30696 33340
rect 33318 33328 33324 33340
rect 33376 33328 33382 33380
rect 34054 33368 34060 33380
rect 34015 33340 34060 33368
rect 34054 33328 34060 33340
rect 34112 33328 34118 33380
rect 34164 33368 34192 33408
rect 34330 33396 34336 33408
rect 34388 33396 34394 33448
rect 34440 33436 34468 33467
rect 35250 33464 35256 33476
rect 35308 33464 35314 33516
rect 35437 33507 35495 33513
rect 35437 33473 35449 33507
rect 35483 33504 35495 33507
rect 35912 33504 35940 33544
rect 36538 33532 36544 33544
rect 36596 33532 36602 33584
rect 38194 33572 38200 33584
rect 36648 33544 38200 33572
rect 36078 33504 36084 33516
rect 35483 33476 35940 33504
rect 36039 33476 36084 33504
rect 35483 33473 35495 33476
rect 35437 33467 35495 33473
rect 36078 33464 36084 33476
rect 36136 33464 36142 33516
rect 36170 33464 36176 33516
rect 36228 33504 36234 33516
rect 36265 33507 36323 33513
rect 36265 33504 36277 33507
rect 36228 33476 36277 33504
rect 36228 33464 36234 33476
rect 36265 33473 36277 33476
rect 36311 33504 36323 33507
rect 36648 33504 36676 33544
rect 38194 33532 38200 33544
rect 38252 33532 38258 33584
rect 37458 33504 37464 33516
rect 36311 33476 36676 33504
rect 37419 33476 37464 33504
rect 36311 33473 36323 33476
rect 36265 33467 36323 33473
rect 37458 33464 37464 33476
rect 37516 33464 37522 33516
rect 38933 33507 38991 33513
rect 38933 33473 38945 33507
rect 38979 33473 38991 33507
rect 38933 33467 38991 33473
rect 39117 33507 39175 33513
rect 39117 33473 39129 33507
rect 39163 33504 39175 33507
rect 39761 33507 39819 33513
rect 39761 33504 39773 33507
rect 39163 33476 39773 33504
rect 39163 33473 39175 33476
rect 39117 33467 39175 33473
rect 39761 33473 39773 33476
rect 39807 33504 39819 33507
rect 40405 33507 40463 33513
rect 40405 33504 40417 33507
rect 39807 33476 40417 33504
rect 39807 33473 39819 33476
rect 39761 33467 39819 33473
rect 40405 33473 40417 33476
rect 40451 33504 40463 33507
rect 40957 33507 41015 33513
rect 40957 33504 40969 33507
rect 40451 33476 40969 33504
rect 40451 33473 40463 33476
rect 40405 33467 40463 33473
rect 40957 33473 40969 33476
rect 41003 33504 41015 33507
rect 41003 33476 41414 33504
rect 41003 33473 41015 33476
rect 40957 33467 41015 33473
rect 35894 33436 35900 33448
rect 34440 33408 35900 33436
rect 35894 33396 35900 33408
rect 35952 33396 35958 33448
rect 37366 33436 37372 33448
rect 37327 33408 37372 33436
rect 37366 33396 37372 33408
rect 37424 33396 37430 33448
rect 37829 33439 37887 33445
rect 37829 33405 37841 33439
rect 37875 33436 37887 33439
rect 38746 33436 38752 33448
rect 37875 33408 38752 33436
rect 37875 33405 37887 33408
rect 37829 33399 37887 33405
rect 38746 33396 38752 33408
rect 38804 33396 38810 33448
rect 38948 33436 38976 33467
rect 39945 33439 40003 33445
rect 39945 33436 39957 33439
rect 38948 33408 39957 33436
rect 39945 33405 39957 33408
rect 39991 33405 40003 33439
rect 39945 33399 40003 33405
rect 39577 33371 39635 33377
rect 39577 33368 39589 33371
rect 34164 33340 39589 33368
rect 39577 33337 39589 33340
rect 39623 33337 39635 33371
rect 39960 33368 39988 33399
rect 40402 33368 40408 33380
rect 39960 33340 40408 33368
rect 39577 33331 39635 33337
rect 40402 33328 40408 33340
rect 40460 33328 40466 33380
rect 28644 33272 29960 33300
rect 30653 33303 30711 33309
rect 26973 33263 27031 33269
rect 30653 33269 30665 33303
rect 30699 33269 30711 33303
rect 30834 33300 30840 33312
rect 30795 33272 30840 33300
rect 30653 33263 30711 33269
rect 30834 33260 30840 33272
rect 30892 33260 30898 33312
rect 32398 33260 32404 33312
rect 32456 33300 32462 33312
rect 39025 33303 39083 33309
rect 39025 33300 39037 33303
rect 32456 33272 39037 33300
rect 32456 33260 32462 33272
rect 39025 33269 39037 33272
rect 39071 33269 39083 33303
rect 41386 33300 41414 33476
rect 53098 33300 53104 33312
rect 41386 33272 53104 33300
rect 39025 33263 39083 33269
rect 53098 33260 53104 33272
rect 53156 33260 53162 33312
rect 1104 33210 54372 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 54372 33210
rect 1104 33136 54372 33158
rect 2038 33056 2044 33108
rect 2096 33096 2102 33108
rect 2096 33068 6914 33096
rect 2096 33056 2102 33068
rect 6886 33028 6914 33068
rect 17954 33056 17960 33108
rect 18012 33096 18018 33108
rect 19245 33099 19303 33105
rect 19245 33096 19257 33099
rect 18012 33068 19257 33096
rect 18012 33056 18018 33068
rect 19245 33065 19257 33068
rect 19291 33065 19303 33099
rect 33597 33099 33655 33105
rect 19245 33059 19303 33065
rect 20640 33068 31754 33096
rect 20640 33028 20668 33068
rect 6886 33000 20668 33028
rect 26234 32988 26240 33040
rect 26292 33028 26298 33040
rect 26605 33031 26663 33037
rect 26605 33028 26617 33031
rect 26292 33000 26617 33028
rect 26292 32988 26298 33000
rect 26605 32997 26617 33000
rect 26651 32997 26663 33031
rect 26605 32991 26663 32997
rect 28258 32988 28264 33040
rect 28316 33028 28322 33040
rect 28905 33031 28963 33037
rect 28905 33028 28917 33031
rect 28316 33000 28917 33028
rect 28316 32988 28322 33000
rect 28905 32997 28917 33000
rect 28951 32997 28963 33031
rect 28905 32991 28963 32997
rect 29086 32988 29092 33040
rect 29144 33028 29150 33040
rect 30742 33028 30748 33040
rect 29144 33000 30748 33028
rect 29144 32988 29150 33000
rect 30742 32988 30748 33000
rect 30800 32988 30806 33040
rect 31726 33028 31754 33068
rect 33597 33065 33609 33099
rect 33643 33096 33655 33099
rect 33686 33096 33692 33108
rect 33643 33068 33692 33096
rect 33643 33065 33655 33068
rect 33597 33059 33655 33065
rect 33686 33056 33692 33068
rect 33744 33056 33750 33108
rect 35342 33096 35348 33108
rect 35303 33068 35348 33096
rect 35342 33056 35348 33068
rect 35400 33056 35406 33108
rect 36078 33056 36084 33108
rect 36136 33096 36142 33108
rect 37921 33099 37979 33105
rect 37921 33096 37933 33099
rect 36136 33068 37933 33096
rect 36136 33056 36142 33068
rect 37921 33065 37933 33068
rect 37967 33096 37979 33099
rect 38286 33096 38292 33108
rect 37967 33068 38292 33096
rect 37967 33065 37979 33068
rect 37921 33059 37979 33065
rect 38286 33056 38292 33068
rect 38344 33096 38350 33108
rect 38930 33096 38936 33108
rect 38344 33068 38936 33096
rect 38344 33056 38350 33068
rect 38930 33056 38936 33068
rect 38988 33056 38994 33108
rect 31726 33000 35848 33028
rect 18325 32963 18383 32969
rect 18325 32929 18337 32963
rect 18371 32960 18383 32963
rect 18414 32960 18420 32972
rect 18371 32932 18420 32960
rect 18371 32929 18383 32932
rect 18325 32923 18383 32929
rect 18414 32920 18420 32932
rect 18472 32920 18478 32972
rect 18966 32920 18972 32972
rect 19024 32960 19030 32972
rect 20809 32963 20867 32969
rect 20809 32960 20821 32963
rect 19024 32932 20821 32960
rect 19024 32920 19030 32932
rect 20809 32929 20821 32932
rect 20855 32929 20867 32963
rect 20809 32923 20867 32929
rect 22925 32963 22983 32969
rect 22925 32929 22937 32963
rect 22971 32960 22983 32963
rect 23290 32960 23296 32972
rect 22971 32932 23296 32960
rect 22971 32929 22983 32932
rect 22925 32923 22983 32929
rect 17954 32852 17960 32904
rect 18012 32892 18018 32904
rect 18049 32895 18107 32901
rect 18049 32892 18061 32895
rect 18012 32864 18061 32892
rect 18012 32852 18018 32864
rect 18049 32861 18061 32864
rect 18095 32861 18107 32895
rect 18049 32855 18107 32861
rect 18141 32895 18199 32901
rect 18141 32861 18153 32895
rect 18187 32892 18199 32895
rect 18506 32892 18512 32904
rect 18187 32864 18512 32892
rect 18187 32861 18199 32864
rect 18141 32855 18199 32861
rect 18506 32852 18512 32864
rect 18564 32852 18570 32904
rect 18598 32852 18604 32904
rect 18656 32892 18662 32904
rect 19245 32895 19303 32901
rect 19245 32892 19257 32895
rect 18656 32864 19257 32892
rect 18656 32852 18662 32864
rect 19245 32861 19257 32864
rect 19291 32861 19303 32895
rect 19245 32855 19303 32861
rect 19337 32895 19395 32901
rect 19337 32861 19349 32895
rect 19383 32861 19395 32895
rect 20070 32892 20076 32904
rect 20031 32864 20076 32892
rect 19337 32855 19395 32861
rect 19352 32824 19380 32855
rect 20070 32852 20076 32864
rect 20128 32852 20134 32904
rect 20254 32892 20260 32904
rect 20215 32864 20260 32892
rect 20254 32852 20260 32864
rect 20312 32852 20318 32904
rect 18156 32796 19380 32824
rect 20824 32824 20852 32923
rect 23290 32920 23296 32932
rect 23348 32920 23354 32972
rect 24486 32960 24492 32972
rect 24447 32932 24492 32960
rect 24486 32920 24492 32932
rect 24544 32920 24550 32972
rect 26418 32960 26424 32972
rect 25700 32932 26424 32960
rect 21450 32852 21456 32904
rect 21508 32892 21514 32904
rect 22002 32892 22008 32904
rect 21508 32864 22008 32892
rect 21508 32852 21514 32864
rect 22002 32852 22008 32864
rect 22060 32892 22066 32904
rect 22097 32895 22155 32901
rect 22097 32892 22109 32895
rect 22060 32864 22109 32892
rect 22060 32852 22066 32864
rect 22097 32861 22109 32864
rect 22143 32861 22155 32895
rect 22097 32855 22155 32861
rect 22554 32852 22560 32904
rect 22612 32892 22618 32904
rect 23109 32895 23167 32901
rect 23109 32892 23121 32895
rect 22612 32864 23121 32892
rect 22612 32852 22618 32864
rect 23109 32861 23121 32864
rect 23155 32861 23167 32895
rect 23109 32855 23167 32861
rect 23198 32852 23204 32904
rect 23256 32892 23262 32904
rect 24581 32895 24639 32901
rect 24581 32892 24593 32895
rect 23256 32864 24593 32892
rect 23256 32852 23262 32864
rect 24581 32861 24593 32864
rect 24627 32861 24639 32895
rect 24581 32855 24639 32861
rect 25409 32895 25467 32901
rect 25409 32861 25421 32895
rect 25455 32861 25467 32895
rect 25590 32892 25596 32904
rect 25551 32864 25596 32892
rect 25409 32855 25467 32861
rect 21910 32824 21916 32836
rect 20824 32796 21916 32824
rect 18156 32768 18184 32796
rect 21910 32784 21916 32796
rect 21968 32784 21974 32836
rect 25424 32824 25452 32855
rect 25590 32852 25596 32864
rect 25648 32852 25654 32904
rect 25700 32901 25728 32932
rect 26418 32920 26424 32932
rect 26476 32920 26482 32972
rect 29546 32960 29552 32972
rect 29012 32932 29552 32960
rect 25685 32895 25743 32901
rect 25685 32861 25697 32895
rect 25731 32861 25743 32895
rect 25685 32855 25743 32861
rect 25774 32852 25780 32904
rect 25832 32892 25838 32904
rect 26510 32892 26516 32904
rect 25832 32864 25877 32892
rect 25976 32864 26516 32892
rect 25832 32852 25838 32864
rect 25976 32824 26004 32864
rect 26510 32852 26516 32864
rect 26568 32852 26574 32904
rect 26970 32852 26976 32904
rect 27028 32892 27034 32904
rect 27985 32895 28043 32901
rect 27985 32892 27997 32895
rect 27028 32864 27997 32892
rect 27028 32852 27034 32864
rect 27985 32861 27997 32864
rect 28031 32861 28043 32895
rect 27985 32855 28043 32861
rect 28718 32852 28724 32904
rect 28776 32892 28782 32904
rect 29012 32901 29040 32932
rect 29546 32920 29552 32932
rect 29604 32960 29610 32972
rect 29641 32963 29699 32969
rect 29641 32960 29653 32963
rect 29604 32932 29653 32960
rect 29604 32920 29610 32932
rect 29641 32929 29653 32932
rect 29687 32960 29699 32963
rect 29914 32960 29920 32972
rect 29687 32932 29920 32960
rect 29687 32929 29699 32932
rect 29641 32923 29699 32929
rect 29914 32920 29920 32932
rect 29972 32920 29978 32972
rect 31386 32960 31392 32972
rect 31128 32932 31392 32960
rect 28813 32895 28871 32901
rect 28813 32892 28825 32895
rect 28776 32864 28825 32892
rect 28776 32852 28782 32864
rect 28813 32861 28825 32864
rect 28859 32861 28871 32895
rect 28813 32855 28871 32861
rect 28997 32895 29055 32901
rect 28997 32861 29009 32895
rect 29043 32861 29055 32895
rect 28997 32855 29055 32861
rect 30285 32895 30343 32901
rect 30285 32861 30297 32895
rect 30331 32892 30343 32895
rect 30834 32892 30840 32904
rect 30331 32864 30840 32892
rect 30331 32861 30343 32864
rect 30285 32855 30343 32861
rect 30834 32852 30840 32864
rect 30892 32852 30898 32904
rect 31128 32901 31156 32932
rect 31386 32920 31392 32932
rect 31444 32920 31450 32972
rect 31662 32920 31668 32972
rect 31720 32960 31726 32972
rect 31720 32932 32444 32960
rect 31720 32920 31726 32932
rect 31113 32895 31171 32901
rect 31113 32861 31125 32895
rect 31159 32861 31171 32895
rect 31113 32855 31171 32861
rect 31202 32852 31208 32904
rect 31260 32892 31266 32904
rect 31297 32895 31355 32901
rect 31297 32892 31309 32895
rect 31260 32864 31309 32892
rect 31260 32852 31266 32864
rect 31297 32861 31309 32864
rect 31343 32892 31355 32895
rect 31570 32892 31576 32904
rect 31343 32864 31576 32892
rect 31343 32861 31355 32864
rect 31297 32855 31355 32861
rect 31570 32852 31576 32864
rect 31628 32892 31634 32904
rect 32416 32901 32444 32932
rect 32490 32920 32496 32972
rect 32548 32960 32554 32972
rect 34238 32960 34244 32972
rect 32548 32932 34244 32960
rect 32548 32920 32554 32932
rect 34238 32920 34244 32932
rect 34296 32920 34302 32972
rect 35820 32960 35848 33000
rect 38010 32988 38016 33040
rect 38068 33028 38074 33040
rect 38381 33031 38439 33037
rect 38381 33028 38393 33031
rect 38068 33000 38393 33028
rect 38068 32988 38074 33000
rect 38381 32997 38393 33000
rect 38427 32997 38439 33031
rect 38381 32991 38439 32997
rect 37642 32960 37648 32972
rect 35820 32932 37648 32960
rect 32309 32895 32367 32901
rect 31628 32864 31754 32892
rect 31628 32852 31634 32864
rect 25424 32796 26004 32824
rect 26053 32827 26111 32833
rect 26053 32793 26065 32827
rect 26099 32824 26111 32827
rect 27718 32827 27776 32833
rect 27718 32824 27730 32827
rect 26099 32796 27730 32824
rect 26099 32793 26111 32796
rect 26053 32787 26111 32793
rect 27718 32793 27730 32796
rect 27764 32793 27776 32827
rect 27718 32787 27776 32793
rect 29638 32784 29644 32836
rect 29696 32824 29702 32836
rect 30101 32827 30159 32833
rect 30101 32824 30113 32827
rect 29696 32796 30113 32824
rect 29696 32784 29702 32796
rect 30101 32793 30113 32796
rect 30147 32793 30159 32827
rect 30101 32787 30159 32793
rect 16850 32756 16856 32768
rect 16811 32728 16856 32756
rect 16850 32716 16856 32728
rect 16908 32716 16914 32768
rect 18138 32716 18144 32768
rect 18196 32716 18202 32768
rect 18322 32756 18328 32768
rect 18283 32728 18328 32756
rect 18322 32716 18328 32728
rect 18380 32716 18386 32768
rect 19242 32716 19248 32768
rect 19300 32756 19306 32768
rect 19426 32756 19432 32768
rect 19300 32728 19432 32756
rect 19300 32716 19306 32728
rect 19426 32716 19432 32728
rect 19484 32756 19490 32768
rect 19613 32759 19671 32765
rect 19613 32756 19625 32759
rect 19484 32728 19625 32756
rect 19484 32716 19490 32728
rect 19613 32725 19625 32728
rect 19659 32725 19671 32759
rect 19613 32719 19671 32725
rect 20165 32759 20223 32765
rect 20165 32725 20177 32759
rect 20211 32756 20223 32759
rect 20714 32756 20720 32768
rect 20211 32728 20720 32756
rect 20211 32725 20223 32728
rect 20165 32719 20223 32725
rect 20714 32716 20720 32728
rect 20772 32716 20778 32768
rect 21358 32756 21364 32768
rect 21319 32728 21364 32756
rect 21358 32716 21364 32728
rect 21416 32716 21422 32768
rect 22281 32759 22339 32765
rect 22281 32725 22293 32759
rect 22327 32756 22339 32759
rect 22646 32756 22652 32768
rect 22327 32728 22652 32756
rect 22327 32725 22339 32728
rect 22281 32719 22339 32725
rect 22646 32716 22652 32728
rect 22704 32756 22710 32768
rect 23014 32756 23020 32768
rect 22704 32728 23020 32756
rect 22704 32716 22710 32728
rect 23014 32716 23020 32728
rect 23072 32716 23078 32768
rect 23290 32756 23296 32768
rect 23251 32728 23296 32756
rect 23290 32716 23296 32728
rect 23348 32716 23354 32768
rect 23845 32759 23903 32765
rect 23845 32725 23857 32759
rect 23891 32756 23903 32759
rect 23934 32756 23940 32768
rect 23891 32728 23940 32756
rect 23891 32725 23903 32728
rect 23845 32719 23903 32725
rect 23934 32716 23940 32728
rect 23992 32716 23998 32768
rect 24949 32759 25007 32765
rect 24949 32725 24961 32759
rect 24995 32756 25007 32759
rect 25498 32756 25504 32768
rect 24995 32728 25504 32756
rect 24995 32725 25007 32728
rect 24949 32719 25007 32725
rect 25498 32716 25504 32728
rect 25556 32716 25562 32768
rect 25774 32716 25780 32768
rect 25832 32756 25838 32768
rect 30282 32756 30288 32768
rect 25832 32728 30288 32756
rect 25832 32716 25838 32728
rect 30282 32716 30288 32728
rect 30340 32716 30346 32768
rect 30374 32716 30380 32768
rect 30432 32756 30438 32768
rect 30469 32759 30527 32765
rect 30469 32756 30481 32759
rect 30432 32728 30481 32756
rect 30432 32716 30438 32728
rect 30469 32725 30481 32728
rect 30515 32725 30527 32759
rect 30926 32756 30932 32768
rect 30887 32728 30932 32756
rect 30469 32719 30527 32725
rect 30926 32716 30932 32728
rect 30984 32716 30990 32768
rect 31726 32756 31754 32864
rect 32309 32861 32321 32895
rect 32355 32861 32367 32895
rect 32309 32855 32367 32861
rect 32401 32895 32459 32901
rect 32401 32861 32413 32895
rect 32447 32861 32459 32895
rect 32401 32855 32459 32861
rect 33045 32895 33103 32901
rect 33045 32861 33057 32895
rect 33091 32892 33103 32895
rect 33502 32892 33508 32904
rect 33091 32864 33508 32892
rect 33091 32861 33103 32864
rect 33045 32855 33103 32861
rect 31938 32784 31944 32836
rect 31996 32824 32002 32836
rect 32125 32827 32183 32833
rect 32125 32824 32137 32827
rect 31996 32796 32137 32824
rect 31996 32784 32002 32796
rect 32125 32793 32137 32796
rect 32171 32793 32183 32827
rect 32324 32824 32352 32855
rect 32858 32824 32864 32836
rect 32324 32796 32864 32824
rect 32125 32787 32183 32793
rect 32858 32784 32864 32796
rect 32916 32784 32922 32836
rect 33060 32756 33088 32855
rect 33502 32852 33508 32864
rect 33560 32892 33566 32904
rect 34149 32895 34207 32901
rect 34149 32892 34161 32895
rect 33560 32864 34161 32892
rect 33560 32852 33566 32864
rect 34149 32861 34161 32864
rect 34195 32892 34207 32895
rect 35066 32892 35072 32904
rect 34195 32864 35072 32892
rect 34195 32861 34207 32864
rect 34149 32855 34207 32861
rect 35066 32852 35072 32864
rect 35124 32852 35130 32904
rect 35345 32895 35403 32901
rect 35345 32861 35357 32895
rect 35391 32892 35403 32895
rect 35710 32892 35716 32904
rect 35391 32864 35716 32892
rect 35391 32861 35403 32864
rect 35345 32855 35403 32861
rect 35710 32852 35716 32864
rect 35768 32852 35774 32904
rect 35820 32901 35848 32932
rect 36832 32901 36860 32932
rect 37642 32920 37648 32932
rect 37700 32960 37706 32972
rect 39853 32963 39911 32969
rect 39853 32960 39865 32963
rect 37700 32932 39865 32960
rect 37700 32920 37706 32932
rect 39853 32929 39865 32932
rect 39899 32929 39911 32963
rect 39853 32923 39911 32929
rect 35805 32895 35863 32901
rect 35805 32861 35817 32895
rect 35851 32861 35863 32895
rect 36633 32895 36691 32901
rect 36633 32892 36645 32895
rect 35805 32855 35863 32861
rect 36004 32864 36645 32892
rect 35526 32784 35532 32836
rect 35584 32824 35590 32836
rect 36004 32833 36032 32864
rect 36633 32861 36645 32864
rect 36679 32861 36691 32895
rect 36633 32855 36691 32861
rect 36817 32895 36875 32901
rect 36817 32861 36829 32895
rect 36863 32861 36875 32895
rect 36817 32855 36875 32861
rect 35989 32827 36047 32833
rect 35989 32824 36001 32827
rect 35584 32796 36001 32824
rect 35584 32784 35590 32796
rect 35989 32793 36001 32796
rect 36035 32793 36047 32827
rect 35989 32787 36047 32793
rect 38010 32784 38016 32836
rect 38068 32824 38074 32836
rect 38654 32824 38660 32836
rect 38068 32796 38660 32824
rect 38068 32784 38074 32796
rect 38654 32784 38660 32796
rect 38712 32784 38718 32836
rect 31726 32728 33088 32756
rect 35161 32759 35219 32765
rect 35161 32725 35173 32759
rect 35207 32756 35219 32759
rect 35710 32756 35716 32768
rect 35207 32728 35716 32756
rect 35207 32725 35219 32728
rect 35161 32719 35219 32725
rect 35710 32716 35716 32728
rect 35768 32716 35774 32768
rect 36173 32759 36231 32765
rect 36173 32725 36185 32759
rect 36219 32756 36231 32759
rect 36630 32756 36636 32768
rect 36219 32728 36636 32756
rect 36219 32725 36231 32728
rect 36173 32719 36231 32725
rect 36630 32716 36636 32728
rect 36688 32716 36694 32768
rect 36722 32716 36728 32768
rect 36780 32756 36786 32768
rect 37369 32759 37427 32765
rect 36780 32728 36825 32756
rect 36780 32716 36786 32728
rect 37369 32725 37381 32759
rect 37415 32756 37427 32759
rect 38194 32756 38200 32768
rect 37415 32728 38200 32756
rect 37415 32725 37427 32728
rect 37369 32719 37427 32725
rect 38194 32716 38200 32728
rect 38252 32716 38258 32768
rect 40402 32756 40408 32768
rect 40363 32728 40408 32756
rect 40402 32716 40408 32728
rect 40460 32716 40466 32768
rect 1104 32666 54372 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 54372 32666
rect 1104 32592 54372 32614
rect 18046 32552 18052 32564
rect 17420 32524 18052 32552
rect 1673 32419 1731 32425
rect 1673 32385 1685 32419
rect 1719 32416 1731 32419
rect 2225 32419 2283 32425
rect 2225 32416 2237 32419
rect 1719 32388 2237 32416
rect 1719 32385 1731 32388
rect 1673 32379 1731 32385
rect 2225 32385 2237 32388
rect 2271 32416 2283 32419
rect 16022 32416 16028 32428
rect 2271 32388 16028 32416
rect 2271 32385 2283 32388
rect 2225 32379 2283 32385
rect 16022 32376 16028 32388
rect 16080 32376 16086 32428
rect 17420 32425 17448 32524
rect 18046 32512 18052 32524
rect 18104 32512 18110 32564
rect 18141 32555 18199 32561
rect 18141 32521 18153 32555
rect 18187 32552 18199 32555
rect 18598 32552 18604 32564
rect 18187 32524 18604 32552
rect 18187 32521 18199 32524
rect 18141 32515 18199 32521
rect 17678 32444 17684 32496
rect 17736 32484 17742 32496
rect 18156 32484 18184 32515
rect 18598 32512 18604 32524
rect 18656 32512 18662 32564
rect 19337 32555 19395 32561
rect 19337 32521 19349 32555
rect 19383 32552 19395 32555
rect 20254 32552 20260 32564
rect 19383 32524 20260 32552
rect 19383 32521 19395 32524
rect 19337 32515 19395 32521
rect 20254 32512 20260 32524
rect 20312 32512 20318 32564
rect 25590 32552 25596 32564
rect 25551 32524 25596 32552
rect 25590 32512 25596 32524
rect 25648 32512 25654 32564
rect 27338 32512 27344 32564
rect 27396 32552 27402 32564
rect 28442 32552 28448 32564
rect 27396 32524 28448 32552
rect 27396 32512 27402 32524
rect 28442 32512 28448 32524
rect 28500 32512 28506 32564
rect 28718 32512 28724 32564
rect 28776 32552 28782 32564
rect 28997 32555 29055 32561
rect 28997 32552 29009 32555
rect 28776 32524 29009 32552
rect 28776 32512 28782 32524
rect 28997 32521 29009 32524
rect 29043 32521 29055 32555
rect 29638 32552 29644 32564
rect 29599 32524 29644 32552
rect 28997 32515 29055 32521
rect 29638 32512 29644 32524
rect 29696 32512 29702 32564
rect 31478 32512 31484 32564
rect 31536 32552 31542 32564
rect 32861 32555 32919 32561
rect 32861 32552 32873 32555
rect 31536 32524 32873 32552
rect 31536 32512 31542 32524
rect 32861 32521 32873 32524
rect 32907 32521 32919 32555
rect 32861 32515 32919 32521
rect 33134 32512 33140 32564
rect 33192 32552 33198 32564
rect 33318 32552 33324 32564
rect 33192 32524 33324 32552
rect 33192 32512 33198 32524
rect 33318 32512 33324 32524
rect 33376 32512 33382 32564
rect 33689 32555 33747 32561
rect 33689 32521 33701 32555
rect 33735 32552 33747 32555
rect 34146 32552 34152 32564
rect 33735 32524 34152 32552
rect 33735 32521 33747 32524
rect 33689 32515 33747 32521
rect 18966 32484 18972 32496
rect 17736 32456 18184 32484
rect 18927 32456 18972 32484
rect 17736 32444 17742 32456
rect 18966 32444 18972 32456
rect 19024 32444 19030 32496
rect 19242 32493 19248 32496
rect 19185 32487 19248 32493
rect 19185 32453 19197 32487
rect 19231 32453 19248 32487
rect 19185 32447 19248 32453
rect 19242 32444 19248 32447
rect 19300 32444 19306 32496
rect 20073 32487 20131 32493
rect 20073 32484 20085 32487
rect 19444 32456 20085 32484
rect 17405 32419 17463 32425
rect 17405 32385 17417 32419
rect 17451 32385 17463 32419
rect 17405 32379 17463 32385
rect 17604 32388 18000 32416
rect 16945 32351 17003 32357
rect 16945 32317 16957 32351
rect 16991 32348 17003 32351
rect 17604 32348 17632 32388
rect 16991 32320 17632 32348
rect 16991 32317 17003 32320
rect 16945 32311 17003 32317
rect 17678 32308 17684 32360
rect 17736 32348 17742 32360
rect 17972 32348 18000 32388
rect 18046 32376 18052 32428
rect 18104 32416 18110 32428
rect 18325 32419 18383 32425
rect 18325 32416 18337 32419
rect 18104 32388 18337 32416
rect 18104 32376 18110 32388
rect 18325 32385 18337 32388
rect 18371 32385 18383 32419
rect 18325 32379 18383 32385
rect 18414 32376 18420 32428
rect 18472 32416 18478 32428
rect 18984 32416 19012 32444
rect 19444 32416 19472 32456
rect 20073 32453 20085 32456
rect 20119 32453 20131 32487
rect 20073 32447 20131 32453
rect 22002 32444 22008 32496
rect 22060 32484 22066 32496
rect 22060 32456 22140 32484
rect 22060 32444 22066 32456
rect 18472 32388 18517 32416
rect 18984 32388 19472 32416
rect 18472 32376 18478 32388
rect 18984 32348 19012 32388
rect 19518 32376 19524 32428
rect 19576 32416 19582 32428
rect 19797 32419 19855 32425
rect 19797 32416 19809 32419
rect 19576 32388 19809 32416
rect 19576 32376 19582 32388
rect 19797 32385 19809 32388
rect 19843 32385 19855 32419
rect 19797 32379 19855 32385
rect 19889 32419 19947 32425
rect 19889 32385 19901 32419
rect 19935 32385 19947 32419
rect 20806 32416 20812 32428
rect 20767 32388 20812 32416
rect 19889 32379 19947 32385
rect 19904 32348 19932 32379
rect 20806 32376 20812 32388
rect 20864 32376 20870 32428
rect 21910 32416 21916 32428
rect 21871 32388 21916 32416
rect 21910 32376 21916 32388
rect 21968 32376 21974 32428
rect 22112 32425 22140 32456
rect 23750 32444 23756 32496
rect 23808 32484 23814 32496
rect 23808 32456 24532 32484
rect 23808 32444 23814 32456
rect 22097 32419 22155 32425
rect 22097 32385 22109 32419
rect 22143 32385 22155 32419
rect 22554 32416 22560 32428
rect 22467 32388 22560 32416
rect 22097 32379 22155 32385
rect 22554 32376 22560 32388
rect 22612 32376 22618 32428
rect 22741 32419 22799 32425
rect 22741 32385 22753 32419
rect 22787 32416 22799 32419
rect 23106 32416 23112 32428
rect 22787 32388 23112 32416
rect 22787 32385 22799 32388
rect 22741 32379 22799 32385
rect 23106 32376 23112 32388
rect 23164 32376 23170 32428
rect 23198 32376 23204 32428
rect 23256 32416 23262 32428
rect 23569 32419 23627 32425
rect 23256 32388 23301 32416
rect 23256 32376 23262 32388
rect 23569 32385 23581 32419
rect 23615 32416 23627 32419
rect 23658 32416 23664 32428
rect 23615 32388 23664 32416
rect 23615 32385 23627 32388
rect 23569 32379 23627 32385
rect 23658 32376 23664 32388
rect 23716 32416 23722 32428
rect 24213 32419 24271 32425
rect 24213 32416 24225 32419
rect 23716 32388 24225 32416
rect 23716 32376 23722 32388
rect 24213 32385 24225 32388
rect 24259 32385 24271 32419
rect 24394 32416 24400 32428
rect 24355 32388 24400 32416
rect 24213 32379 24271 32385
rect 24394 32376 24400 32388
rect 24452 32376 24458 32428
rect 24504 32425 24532 32456
rect 25314 32444 25320 32496
rect 25372 32484 25378 32496
rect 26973 32487 27031 32493
rect 26973 32484 26985 32487
rect 25372 32456 26985 32484
rect 25372 32444 25378 32456
rect 24489 32419 24547 32425
rect 24489 32385 24501 32419
rect 24535 32385 24547 32419
rect 25498 32416 25504 32428
rect 25459 32388 25504 32416
rect 24489 32379 24547 32385
rect 25498 32376 25504 32388
rect 25556 32376 25562 32428
rect 25700 32425 25728 32456
rect 26973 32453 26985 32456
rect 27019 32484 27031 32487
rect 30098 32484 30104 32496
rect 27019 32456 30104 32484
rect 27019 32453 27031 32456
rect 26973 32447 27031 32453
rect 30098 32444 30104 32456
rect 30156 32444 30162 32496
rect 30581 32487 30639 32493
rect 30581 32453 30593 32487
rect 30627 32484 30639 32487
rect 30834 32484 30840 32496
rect 30627 32456 30840 32484
rect 30627 32453 30639 32456
rect 30581 32447 30639 32453
rect 30834 32444 30840 32456
rect 30892 32484 30898 32496
rect 33594 32484 33600 32496
rect 30892 32456 33600 32484
rect 30892 32444 30898 32456
rect 33594 32444 33600 32456
rect 33652 32484 33658 32496
rect 33704 32484 33732 32515
rect 34146 32512 34152 32524
rect 34204 32512 34210 32564
rect 35802 32552 35808 32564
rect 35763 32524 35808 32552
rect 35802 32512 35808 32524
rect 35860 32512 35866 32564
rect 37277 32555 37335 32561
rect 37277 32521 37289 32555
rect 37323 32552 37335 32555
rect 37458 32552 37464 32564
rect 37323 32524 37464 32552
rect 37323 32521 37335 32524
rect 37277 32515 37335 32521
rect 37458 32512 37464 32524
rect 37516 32512 37522 32564
rect 38194 32552 38200 32564
rect 38155 32524 38200 32552
rect 38194 32512 38200 32524
rect 38252 32512 38258 32564
rect 38654 32552 38660 32564
rect 38615 32524 38660 32552
rect 38654 32512 38660 32524
rect 38712 32512 38718 32564
rect 33652 32456 33732 32484
rect 33652 32444 33658 32456
rect 35066 32444 35072 32496
rect 35124 32484 35130 32496
rect 36170 32484 36176 32496
rect 35124 32456 36176 32484
rect 35124 32444 35130 32456
rect 25685 32419 25743 32425
rect 25685 32385 25697 32419
rect 25731 32385 25743 32419
rect 29546 32416 29552 32428
rect 29507 32388 29552 32416
rect 25685 32379 25743 32385
rect 29546 32376 29552 32388
rect 29604 32376 29610 32428
rect 29730 32416 29736 32428
rect 29691 32388 29736 32416
rect 29730 32376 29736 32388
rect 29788 32376 29794 32428
rect 30193 32419 30251 32425
rect 30193 32385 30205 32419
rect 30239 32385 30251 32419
rect 30193 32379 30251 32385
rect 30286 32419 30344 32425
rect 30286 32385 30298 32419
rect 30332 32385 30344 32419
rect 30286 32379 30344 32385
rect 30469 32419 30527 32425
rect 30469 32385 30481 32419
rect 30515 32414 30527 32419
rect 30699 32419 30757 32425
rect 30515 32386 30604 32414
rect 30515 32385 30527 32386
rect 30469 32379 30527 32385
rect 20714 32348 20720 32360
rect 17736 32320 17781 32348
rect 17972 32320 19012 32348
rect 19168 32320 19932 32348
rect 20675 32320 20720 32348
rect 17736 32308 17742 32320
rect 17589 32283 17647 32289
rect 17589 32249 17601 32283
rect 17635 32280 17647 32283
rect 19168 32280 19196 32320
rect 20714 32308 20720 32320
rect 20772 32308 20778 32360
rect 22005 32351 22063 32357
rect 22005 32317 22017 32351
rect 22051 32348 22063 32351
rect 22572 32348 22600 32376
rect 22051 32320 22600 32348
rect 22051 32317 22063 32320
rect 22005 32311 22063 32317
rect 28902 32308 28908 32360
rect 28960 32348 28966 32360
rect 30208 32348 30236 32379
rect 28960 32320 30236 32348
rect 28960 32308 28966 32320
rect 20070 32280 20076 32292
rect 17635 32252 19196 32280
rect 20031 32252 20076 32280
rect 17635 32249 17647 32252
rect 17589 32243 17647 32249
rect 1486 32212 1492 32224
rect 1447 32184 1492 32212
rect 1486 32172 1492 32184
rect 1544 32172 1550 32224
rect 17497 32215 17555 32221
rect 17497 32181 17509 32215
rect 17543 32212 17555 32215
rect 17954 32212 17960 32224
rect 17543 32184 17960 32212
rect 17543 32181 17555 32184
rect 17497 32175 17555 32181
rect 17954 32172 17960 32184
rect 18012 32212 18018 32224
rect 18690 32212 18696 32224
rect 18012 32184 18696 32212
rect 18012 32172 18018 32184
rect 18690 32172 18696 32184
rect 18748 32172 18754 32224
rect 19168 32221 19196 32252
rect 20070 32240 20076 32252
rect 20128 32240 20134 32292
rect 21177 32283 21235 32289
rect 21177 32249 21189 32283
rect 21223 32280 21235 32283
rect 23382 32280 23388 32292
rect 21223 32252 23388 32280
rect 21223 32249 21235 32252
rect 21177 32243 21235 32249
rect 23382 32240 23388 32252
rect 23440 32240 23446 32292
rect 28442 32240 28448 32292
rect 28500 32280 28506 32292
rect 30300 32280 30328 32379
rect 30374 32308 30380 32360
rect 30432 32348 30438 32360
rect 30576 32348 30604 32386
rect 30699 32385 30711 32419
rect 30745 32385 30757 32419
rect 30699 32379 30757 32385
rect 30432 32320 30604 32348
rect 30432 32308 30438 32320
rect 28500 32252 30328 32280
rect 28500 32240 28506 32252
rect 30466 32240 30472 32292
rect 30524 32280 30530 32292
rect 30700 32280 30728 32379
rect 31202 32376 31208 32428
rect 31260 32416 31266 32428
rect 31297 32419 31355 32425
rect 31297 32416 31309 32419
rect 31260 32388 31309 32416
rect 31260 32376 31266 32388
rect 31297 32385 31309 32388
rect 31343 32385 31355 32419
rect 31297 32379 31355 32385
rect 31662 32376 31668 32428
rect 31720 32416 31726 32428
rect 31720 32388 32168 32416
rect 31720 32376 31726 32388
rect 31573 32351 31631 32357
rect 31573 32317 31585 32351
rect 31619 32348 31631 32351
rect 31938 32348 31944 32360
rect 31619 32320 31944 32348
rect 31619 32317 31631 32320
rect 31573 32311 31631 32317
rect 31938 32308 31944 32320
rect 31996 32308 32002 32360
rect 32140 32357 32168 32388
rect 32214 32376 32220 32428
rect 32272 32416 32278 32428
rect 32309 32419 32367 32425
rect 32309 32416 32321 32419
rect 32272 32388 32321 32416
rect 32272 32376 32278 32388
rect 32309 32385 32321 32388
rect 32355 32385 32367 32419
rect 32309 32379 32367 32385
rect 32401 32419 32459 32425
rect 32401 32385 32413 32419
rect 32447 32416 32459 32419
rect 32674 32416 32680 32428
rect 32447 32388 32680 32416
rect 32447 32385 32459 32388
rect 32401 32379 32459 32385
rect 32674 32376 32680 32388
rect 32732 32376 32738 32428
rect 32858 32416 32864 32428
rect 32819 32388 32864 32416
rect 32858 32376 32864 32388
rect 32916 32376 32922 32428
rect 32950 32376 32956 32428
rect 33008 32416 33014 32428
rect 35636 32425 35664 32456
rect 36170 32444 36176 32456
rect 36228 32444 36234 32496
rect 33137 32419 33195 32425
rect 33137 32416 33149 32419
rect 33008 32388 33149 32416
rect 33008 32376 33014 32388
rect 33137 32385 33149 32388
rect 33183 32385 33195 32419
rect 33137 32379 33195 32385
rect 35621 32419 35679 32425
rect 35621 32385 35633 32419
rect 35667 32385 35679 32419
rect 35621 32379 35679 32385
rect 35710 32376 35716 32428
rect 35768 32416 35774 32428
rect 35805 32419 35863 32425
rect 35805 32416 35817 32419
rect 35768 32388 35817 32416
rect 35768 32376 35774 32388
rect 35805 32385 35817 32388
rect 35851 32416 35863 32419
rect 36078 32416 36084 32428
rect 35851 32388 36084 32416
rect 35851 32385 35863 32388
rect 35805 32379 35863 32385
rect 36078 32376 36084 32388
rect 36136 32376 36142 32428
rect 36262 32416 36268 32428
rect 36223 32388 36268 32416
rect 36262 32376 36268 32388
rect 36320 32376 36326 32428
rect 36630 32376 36636 32428
rect 36688 32416 36694 32428
rect 37461 32419 37519 32425
rect 37461 32416 37473 32419
rect 36688 32388 37473 32416
rect 36688 32376 36694 32388
rect 37461 32385 37473 32388
rect 37507 32385 37519 32419
rect 37461 32379 37519 32385
rect 52917 32419 52975 32425
rect 52917 32385 52929 32419
rect 52963 32416 52975 32419
rect 53558 32416 53564 32428
rect 52963 32388 53564 32416
rect 52963 32385 52975 32388
rect 52917 32379 52975 32385
rect 53558 32376 53564 32388
rect 53616 32376 53622 32428
rect 32125 32351 32183 32357
rect 32125 32317 32137 32351
rect 32171 32348 32183 32351
rect 32171 32320 34284 32348
rect 32171 32317 32183 32320
rect 32125 32311 32183 32317
rect 30524 32252 30728 32280
rect 30837 32283 30895 32289
rect 30524 32240 30530 32252
rect 30837 32249 30849 32283
rect 30883 32280 30895 32283
rect 32490 32280 32496 32292
rect 30883 32252 32496 32280
rect 30883 32249 30895 32252
rect 30837 32243 30895 32249
rect 32490 32240 32496 32252
rect 32548 32240 32554 32292
rect 32953 32283 33011 32289
rect 32953 32249 32965 32283
rect 32999 32280 33011 32283
rect 33042 32280 33048 32292
rect 32999 32252 33048 32280
rect 32999 32249 33011 32252
rect 32953 32243 33011 32249
rect 33042 32240 33048 32252
rect 33100 32240 33106 32292
rect 19153 32215 19211 32221
rect 19153 32181 19165 32215
rect 19199 32181 19211 32215
rect 22646 32212 22652 32224
rect 22607 32184 22652 32212
rect 19153 32175 19211 32181
rect 22646 32172 22652 32184
rect 22704 32172 22710 32224
rect 23290 32212 23296 32224
rect 23251 32184 23296 32212
rect 23290 32172 23296 32184
rect 23348 32172 23354 32224
rect 23750 32212 23756 32224
rect 23711 32184 23756 32212
rect 23750 32172 23756 32184
rect 23808 32172 23814 32224
rect 23842 32172 23848 32224
rect 23900 32212 23906 32224
rect 24213 32215 24271 32221
rect 24213 32212 24225 32215
rect 23900 32184 24225 32212
rect 23900 32172 23906 32184
rect 24213 32181 24225 32184
rect 24259 32181 24271 32215
rect 24670 32212 24676 32224
rect 24631 32184 24676 32212
rect 24213 32175 24271 32181
rect 24670 32172 24676 32184
rect 24728 32172 24734 32224
rect 25590 32172 25596 32224
rect 25648 32212 25654 32224
rect 26145 32215 26203 32221
rect 26145 32212 26157 32215
rect 25648 32184 26157 32212
rect 25648 32172 25654 32184
rect 26145 32181 26157 32184
rect 26191 32212 26203 32215
rect 27706 32212 27712 32224
rect 26191 32184 27712 32212
rect 26191 32181 26203 32184
rect 26145 32175 26203 32181
rect 27706 32172 27712 32184
rect 27764 32172 27770 32224
rect 29730 32172 29736 32224
rect 29788 32212 29794 32224
rect 30926 32212 30932 32224
rect 29788 32184 30932 32212
rect 29788 32172 29794 32184
rect 30926 32172 30932 32184
rect 30984 32172 30990 32224
rect 31386 32212 31392 32224
rect 31347 32184 31392 32212
rect 31386 32172 31392 32184
rect 31444 32172 31450 32224
rect 31478 32172 31484 32224
rect 31536 32212 31542 32224
rect 31536 32184 31581 32212
rect 31536 32172 31542 32184
rect 31662 32172 31668 32224
rect 31720 32212 31726 32224
rect 34256 32221 34284 32320
rect 36722 32308 36728 32360
rect 36780 32348 36786 32360
rect 37642 32348 37648 32360
rect 36780 32320 37648 32348
rect 36780 32308 36786 32320
rect 37642 32308 37648 32320
rect 37700 32308 37706 32360
rect 53374 32280 53380 32292
rect 53335 32252 53380 32280
rect 53374 32240 53380 32252
rect 53432 32240 53438 32292
rect 32217 32215 32275 32221
rect 32217 32212 32229 32215
rect 31720 32184 32229 32212
rect 31720 32172 31726 32184
rect 32217 32181 32229 32184
rect 32263 32181 32275 32215
rect 32217 32175 32275 32181
rect 34241 32215 34299 32221
rect 34241 32181 34253 32215
rect 34287 32212 34299 32215
rect 34330 32212 34336 32224
rect 34287 32184 34336 32212
rect 34287 32181 34299 32184
rect 34241 32175 34299 32181
rect 34330 32172 34336 32184
rect 34388 32172 34394 32224
rect 34698 32212 34704 32224
rect 34659 32184 34704 32212
rect 34698 32172 34704 32184
rect 34756 32172 34762 32224
rect 36354 32212 36360 32224
rect 36315 32184 36360 32212
rect 36354 32172 36360 32184
rect 36412 32172 36418 32224
rect 1104 32122 54372 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 54372 32122
rect 1104 32048 54372 32070
rect 15378 31968 15384 32020
rect 15436 32008 15442 32020
rect 15473 32011 15531 32017
rect 15473 32008 15485 32011
rect 15436 31980 15485 32008
rect 15436 31968 15442 31980
rect 15473 31977 15485 31980
rect 15519 32008 15531 32011
rect 16025 32011 16083 32017
rect 16025 32008 16037 32011
rect 15519 31980 16037 32008
rect 15519 31977 15531 31980
rect 15473 31971 15531 31977
rect 16025 31977 16037 31980
rect 16071 31977 16083 32011
rect 18138 32008 18144 32020
rect 18099 31980 18144 32008
rect 16025 31971 16083 31977
rect 16040 31940 16068 31971
rect 18138 31968 18144 31980
rect 18196 31968 18202 32020
rect 18506 32008 18512 32020
rect 18467 31980 18512 32008
rect 18506 31968 18512 31980
rect 18564 31968 18570 32020
rect 23477 32011 23535 32017
rect 23477 31977 23489 32011
rect 23523 32008 23535 32011
rect 24489 32011 24547 32017
rect 24489 32008 24501 32011
rect 23523 31980 24501 32008
rect 23523 31977 23535 31980
rect 23477 31971 23535 31977
rect 24489 31977 24501 31980
rect 24535 31977 24547 32011
rect 24489 31971 24547 31977
rect 26142 31968 26148 32020
rect 26200 32008 26206 32020
rect 26421 32011 26479 32017
rect 26421 32008 26433 32011
rect 26200 31980 26433 32008
rect 26200 31968 26206 31980
rect 26421 31977 26433 31980
rect 26467 32008 26479 32011
rect 31386 32008 31392 32020
rect 26467 31980 31392 32008
rect 26467 31977 26479 31980
rect 26421 31971 26479 31977
rect 31386 31968 31392 31980
rect 31444 31968 31450 32020
rect 31662 32008 31668 32020
rect 31623 31980 31668 32008
rect 31662 31968 31668 31980
rect 31720 31968 31726 32020
rect 34054 32008 34060 32020
rect 31772 31980 34060 32008
rect 16390 31940 16396 31952
rect 16040 31912 16396 31940
rect 16390 31900 16396 31912
rect 16448 31940 16454 31952
rect 16448 31912 17632 31940
rect 16448 31900 16454 31912
rect 2222 31832 2228 31884
rect 2280 31872 2286 31884
rect 16022 31872 16028 31884
rect 2280 31844 16028 31872
rect 2280 31832 2286 31844
rect 16022 31832 16028 31844
rect 16080 31872 16086 31884
rect 17604 31881 17632 31912
rect 18414 31900 18420 31952
rect 18472 31940 18478 31952
rect 19245 31943 19303 31949
rect 19245 31940 19257 31943
rect 18472 31912 19257 31940
rect 18472 31900 18478 31912
rect 19245 31909 19257 31912
rect 19291 31909 19303 31943
rect 19245 31903 19303 31909
rect 25593 31943 25651 31949
rect 25593 31909 25605 31943
rect 25639 31940 25651 31943
rect 27246 31940 27252 31952
rect 25639 31912 27252 31940
rect 25639 31909 25651 31912
rect 25593 31903 25651 31909
rect 27246 31900 27252 31912
rect 27304 31900 27310 31952
rect 28994 31900 29000 31952
rect 29052 31940 29058 31952
rect 29733 31943 29791 31949
rect 29052 31912 29097 31940
rect 29052 31900 29058 31912
rect 29733 31909 29745 31943
rect 29779 31940 29791 31943
rect 29914 31940 29920 31952
rect 29779 31912 29920 31940
rect 29779 31909 29791 31912
rect 29733 31903 29791 31909
rect 29914 31900 29920 31912
rect 29972 31900 29978 31952
rect 31772 31940 31800 31980
rect 34054 31968 34060 31980
rect 34112 31968 34118 32020
rect 30392 31912 31800 31940
rect 33045 31943 33103 31949
rect 17589 31875 17647 31881
rect 16080 31844 16804 31872
rect 16080 31832 16086 31844
rect 16390 31764 16396 31816
rect 16448 31804 16454 31816
rect 16776 31813 16804 31844
rect 17589 31841 17601 31875
rect 17635 31872 17647 31875
rect 21358 31872 21364 31884
rect 17635 31844 21364 31872
rect 17635 31841 17647 31844
rect 17589 31835 17647 31841
rect 21358 31832 21364 31844
rect 21416 31872 21422 31884
rect 21637 31875 21695 31881
rect 21416 31844 21496 31872
rect 21416 31832 21422 31844
rect 16577 31807 16635 31813
rect 16577 31804 16589 31807
rect 16448 31776 16589 31804
rect 16448 31764 16454 31776
rect 16577 31773 16589 31776
rect 16623 31773 16635 31807
rect 16577 31767 16635 31773
rect 16761 31807 16819 31813
rect 16761 31773 16773 31807
rect 16807 31804 16819 31807
rect 16850 31804 16856 31816
rect 16807 31776 16856 31804
rect 16807 31773 16819 31776
rect 16761 31767 16819 31773
rect 16850 31764 16856 31776
rect 16908 31804 16914 31816
rect 17405 31807 17463 31813
rect 17405 31804 17417 31807
rect 16908 31776 17417 31804
rect 16908 31764 16914 31776
rect 17405 31773 17417 31776
rect 17451 31773 17463 31807
rect 18046 31804 18052 31816
rect 18007 31776 18052 31804
rect 17405 31767 17463 31773
rect 18046 31764 18052 31776
rect 18104 31764 18110 31816
rect 19334 31804 19340 31816
rect 19247 31776 19340 31804
rect 19334 31764 19340 31776
rect 19392 31804 19398 31816
rect 19613 31807 19671 31813
rect 19613 31804 19625 31807
rect 19392 31776 19625 31804
rect 19392 31764 19398 31776
rect 19613 31773 19625 31776
rect 19659 31773 19671 31807
rect 19613 31767 19671 31773
rect 20254 31764 20260 31816
rect 20312 31804 20318 31816
rect 20441 31807 20499 31813
rect 20441 31804 20453 31807
rect 20312 31776 20453 31804
rect 20312 31764 20318 31776
rect 20441 31773 20453 31776
rect 20487 31773 20499 31807
rect 20714 31804 20720 31816
rect 20675 31776 20720 31804
rect 20441 31767 20499 31773
rect 20714 31764 20720 31776
rect 20772 31804 20778 31816
rect 20990 31804 20996 31816
rect 20772 31776 20996 31804
rect 20772 31764 20778 31776
rect 20990 31764 20996 31776
rect 21048 31764 21054 31816
rect 21468 31813 21496 31844
rect 21637 31841 21649 31875
rect 21683 31872 21695 31875
rect 21683 31844 22324 31872
rect 21683 31841 21695 31844
rect 21637 31835 21695 31841
rect 21453 31807 21511 31813
rect 21453 31773 21465 31807
rect 21499 31773 21511 31807
rect 22186 31804 22192 31816
rect 22147 31776 22192 31804
rect 21453 31767 21511 31773
rect 22186 31764 22192 31776
rect 22244 31764 22250 31816
rect 22296 31813 22324 31844
rect 24026 31832 24032 31884
rect 24084 31872 24090 31884
rect 24673 31875 24731 31881
rect 24673 31872 24685 31875
rect 24084 31844 24685 31872
rect 24084 31832 24090 31844
rect 24673 31841 24685 31844
rect 24719 31872 24731 31875
rect 24719 31844 27016 31872
rect 24719 31841 24731 31844
rect 24673 31835 24731 31841
rect 22281 31807 22339 31813
rect 22281 31773 22293 31807
rect 22327 31773 22339 31807
rect 22281 31767 22339 31773
rect 22646 31764 22652 31816
rect 22704 31804 22710 31816
rect 23201 31807 23259 31813
rect 23201 31804 23213 31807
rect 22704 31776 23213 31804
rect 22704 31764 22710 31776
rect 23201 31773 23213 31776
rect 23247 31773 23259 31807
rect 23477 31807 23535 31813
rect 23477 31804 23489 31807
rect 23201 31767 23259 31773
rect 23308 31776 23489 31804
rect 17954 31696 17960 31748
rect 18012 31736 18018 31748
rect 19352 31736 19380 31764
rect 18012 31708 19380 31736
rect 19429 31739 19487 31745
rect 18012 31696 18018 31708
rect 19429 31705 19441 31739
rect 19475 31736 19487 31739
rect 20530 31736 20536 31748
rect 19475 31708 20536 31736
rect 19475 31705 19487 31708
rect 19429 31699 19487 31705
rect 16669 31671 16727 31677
rect 16669 31637 16681 31671
rect 16715 31668 16727 31671
rect 16942 31668 16948 31680
rect 16715 31640 16948 31668
rect 16715 31637 16727 31640
rect 16669 31631 16727 31637
rect 16942 31628 16948 31640
rect 17000 31628 17006 31680
rect 17218 31668 17224 31680
rect 17179 31640 17224 31668
rect 17218 31628 17224 31640
rect 17276 31628 17282 31680
rect 17586 31628 17592 31680
rect 17644 31668 17650 31680
rect 19444 31668 19472 31699
rect 20530 31696 20536 31708
rect 20588 31696 20594 31748
rect 20625 31739 20683 31745
rect 20625 31705 20637 31739
rect 20671 31736 20683 31739
rect 20806 31736 20812 31748
rect 20671 31708 20812 31736
rect 20671 31705 20683 31708
rect 20625 31699 20683 31705
rect 20806 31696 20812 31708
rect 20864 31696 20870 31748
rect 21266 31736 21272 31748
rect 21227 31708 21272 31736
rect 21266 31696 21272 31708
rect 21324 31696 21330 31748
rect 22465 31739 22523 31745
rect 22465 31705 22477 31739
rect 22511 31736 22523 31739
rect 23106 31736 23112 31748
rect 22511 31708 23112 31736
rect 22511 31705 22523 31708
rect 22465 31699 22523 31705
rect 23106 31696 23112 31708
rect 23164 31736 23170 31748
rect 23308 31736 23336 31776
rect 23477 31773 23489 31776
rect 23523 31773 23535 31807
rect 23477 31767 23535 31773
rect 23566 31764 23572 31816
rect 23624 31804 23630 31816
rect 24397 31807 24455 31813
rect 24397 31804 24409 31807
rect 23624 31776 24409 31804
rect 23624 31764 23630 31776
rect 24397 31773 24409 31776
rect 24443 31773 24455 31807
rect 25777 31807 25835 31813
rect 25777 31804 25789 31807
rect 24397 31767 24455 31773
rect 24964 31776 25789 31804
rect 23164 31708 23336 31736
rect 23164 31696 23170 31708
rect 17644 31640 19472 31668
rect 20257 31671 20315 31677
rect 17644 31628 17650 31640
rect 20257 31637 20269 31671
rect 20303 31668 20315 31671
rect 20438 31668 20444 31680
rect 20303 31640 20444 31668
rect 20303 31637 20315 31640
rect 20257 31631 20315 31637
rect 20438 31628 20444 31640
rect 20496 31628 20502 31680
rect 22554 31628 22560 31680
rect 22612 31668 22618 31680
rect 23198 31668 23204 31680
rect 22612 31640 23204 31668
rect 22612 31628 22618 31640
rect 23198 31628 23204 31640
rect 23256 31668 23262 31680
rect 24964 31677 24992 31776
rect 25777 31773 25789 31776
rect 25823 31773 25835 31807
rect 25777 31767 25835 31773
rect 25866 31764 25872 31816
rect 25924 31804 25930 31816
rect 25924 31776 25969 31804
rect 25924 31764 25930 31776
rect 26142 31764 26148 31816
rect 26200 31804 26206 31816
rect 26988 31813 27016 31844
rect 30392 31813 30420 31912
rect 33045 31909 33057 31943
rect 33091 31909 33103 31943
rect 33045 31903 33103 31909
rect 30653 31875 30711 31881
rect 30653 31841 30665 31875
rect 30699 31872 30711 31875
rect 31205 31875 31263 31881
rect 31205 31872 31217 31875
rect 30699 31844 31217 31872
rect 30699 31841 30711 31844
rect 30653 31835 30711 31841
rect 31205 31841 31217 31844
rect 31251 31841 31263 31875
rect 31205 31835 31263 31841
rect 32585 31875 32643 31881
rect 32585 31841 32597 31875
rect 32631 31872 32643 31875
rect 32674 31872 32680 31884
rect 32631 31844 32680 31872
rect 32631 31841 32643 31844
rect 32585 31835 32643 31841
rect 32674 31832 32680 31844
rect 32732 31872 32738 31884
rect 33060 31872 33088 31903
rect 33134 31900 33140 31952
rect 33192 31940 33198 31952
rect 33689 31943 33747 31949
rect 33689 31940 33701 31943
rect 33192 31912 33701 31940
rect 33192 31900 33198 31912
rect 33689 31909 33701 31912
rect 33735 31909 33747 31943
rect 33689 31903 33747 31909
rect 34330 31900 34336 31952
rect 34388 31940 34394 31952
rect 34701 31943 34759 31949
rect 34701 31940 34713 31943
rect 34388 31912 34713 31940
rect 34388 31900 34394 31912
rect 34701 31909 34713 31912
rect 34747 31909 34759 31943
rect 34701 31903 34759 31909
rect 36081 31943 36139 31949
rect 36081 31909 36093 31943
rect 36127 31940 36139 31943
rect 36262 31940 36268 31952
rect 36127 31912 36268 31940
rect 36127 31909 36139 31912
rect 36081 31903 36139 31909
rect 36262 31900 36268 31912
rect 36320 31900 36326 31952
rect 36817 31943 36875 31949
rect 36817 31909 36829 31943
rect 36863 31940 36875 31943
rect 37090 31940 37096 31952
rect 36863 31912 37096 31940
rect 36863 31909 36875 31912
rect 36817 31903 36875 31909
rect 37090 31900 37096 31912
rect 37148 31900 37154 31952
rect 37458 31900 37464 31952
rect 37516 31940 37522 31952
rect 37516 31912 37596 31940
rect 37516 31900 37522 31912
rect 32732 31844 33088 31872
rect 32732 31832 32738 31844
rect 33778 31832 33784 31884
rect 33836 31872 33842 31884
rect 36630 31872 36636 31884
rect 33836 31844 34192 31872
rect 36591 31844 36636 31872
rect 33836 31832 33842 31844
rect 26973 31807 27031 31813
rect 26200 31764 26234 31804
rect 26973 31773 26985 31807
rect 27019 31804 27031 31807
rect 30377 31807 30435 31813
rect 27019 31776 30329 31804
rect 27019 31773 27031 31776
rect 26973 31767 27031 31773
rect 25590 31736 25596 31748
rect 25551 31708 25596 31736
rect 25590 31696 25596 31708
rect 25648 31696 25654 31748
rect 23293 31671 23351 31677
rect 23293 31668 23305 31671
rect 23256 31640 23305 31668
rect 23256 31628 23262 31640
rect 23293 31637 23305 31640
rect 23339 31637 23351 31671
rect 23293 31631 23351 31637
rect 24949 31671 25007 31677
rect 24949 31637 24961 31671
rect 24995 31637 25007 31671
rect 24949 31631 25007 31637
rect 25498 31628 25504 31680
rect 25556 31668 25562 31680
rect 26206 31668 26234 31764
rect 27706 31696 27712 31748
rect 27764 31736 27770 31748
rect 28902 31736 28908 31748
rect 27764 31708 28908 31736
rect 27764 31696 27770 31708
rect 28902 31696 28908 31708
rect 28960 31696 28966 31748
rect 25556 31640 26234 31668
rect 25556 31628 25562 31640
rect 29546 31628 29552 31680
rect 29604 31668 29610 31680
rect 30193 31671 30251 31677
rect 30193 31668 30205 31671
rect 29604 31640 30205 31668
rect 29604 31628 29610 31640
rect 30193 31637 30205 31640
rect 30239 31637 30251 31671
rect 30301 31668 30329 31776
rect 30377 31773 30389 31807
rect 30423 31773 30435 31807
rect 30377 31767 30435 31773
rect 30469 31807 30527 31813
rect 30469 31773 30481 31807
rect 30515 31804 30527 31807
rect 30745 31807 30803 31813
rect 30515 31776 30604 31804
rect 30515 31773 30527 31776
rect 30469 31767 30527 31773
rect 30576 31668 30604 31776
rect 30745 31773 30757 31807
rect 30791 31804 30803 31807
rect 30834 31804 30840 31816
rect 30791 31776 30840 31804
rect 30791 31773 30803 31776
rect 30745 31767 30803 31773
rect 30834 31764 30840 31776
rect 30892 31764 30898 31816
rect 30926 31764 30932 31816
rect 30984 31804 30990 31816
rect 31389 31807 31447 31813
rect 31389 31804 31401 31807
rect 30984 31776 31401 31804
rect 30984 31764 30990 31776
rect 31389 31773 31401 31776
rect 31435 31773 31447 31807
rect 31389 31767 31447 31773
rect 31478 31764 31484 31816
rect 31536 31804 31542 31816
rect 31536 31776 31581 31804
rect 31536 31764 31542 31776
rect 31754 31764 31760 31816
rect 31812 31804 31818 31816
rect 32217 31807 32275 31813
rect 32217 31804 32229 31807
rect 31812 31776 32229 31804
rect 31812 31764 31818 31776
rect 32217 31773 32229 31776
rect 32263 31773 32275 31807
rect 32217 31767 32275 31773
rect 32306 31764 32312 31816
rect 32364 31804 32370 31816
rect 32401 31807 32459 31813
rect 32401 31804 32413 31807
rect 32364 31776 32413 31804
rect 32364 31764 32370 31776
rect 32401 31773 32413 31776
rect 32447 31773 32459 31807
rect 33042 31804 33048 31816
rect 33003 31776 33048 31804
rect 32401 31767 32459 31773
rect 33042 31764 33048 31776
rect 33100 31764 33106 31816
rect 33229 31807 33287 31813
rect 33229 31804 33241 31807
rect 33152 31776 33241 31804
rect 32950 31696 32956 31748
rect 33008 31736 33014 31748
rect 33152 31736 33180 31776
rect 33229 31773 33241 31776
rect 33275 31773 33287 31807
rect 33870 31804 33876 31816
rect 33831 31776 33876 31804
rect 33229 31767 33287 31773
rect 33870 31764 33876 31776
rect 33928 31764 33934 31816
rect 34164 31813 34192 31844
rect 36630 31832 36636 31844
rect 36688 31832 36694 31884
rect 37568 31881 37596 31912
rect 37553 31875 37611 31881
rect 37553 31841 37565 31875
rect 37599 31841 37611 31875
rect 37553 31835 37611 31841
rect 37642 31832 37648 31884
rect 37700 31872 37706 31884
rect 37921 31875 37979 31881
rect 37921 31872 37933 31875
rect 37700 31844 37933 31872
rect 37700 31832 37706 31844
rect 37921 31841 37933 31844
rect 37967 31841 37979 31875
rect 37921 31835 37979 31841
rect 34149 31807 34207 31813
rect 34149 31773 34161 31807
rect 34195 31773 34207 31807
rect 34149 31767 34207 31773
rect 34698 31764 34704 31816
rect 34756 31804 34762 31816
rect 35345 31807 35403 31813
rect 35345 31804 35357 31807
rect 34756 31776 35357 31804
rect 34756 31764 34762 31776
rect 35345 31773 35357 31776
rect 35391 31804 35403 31807
rect 36541 31807 36599 31813
rect 35391 31776 36216 31804
rect 35391 31773 35403 31776
rect 35345 31767 35403 31773
rect 34054 31736 34060 31748
rect 33008 31708 33180 31736
rect 33967 31708 34060 31736
rect 33008 31696 33014 31708
rect 34054 31696 34060 31708
rect 34112 31736 34118 31748
rect 34716 31736 34744 31764
rect 34112 31708 34744 31736
rect 34112 31696 34118 31708
rect 35986 31696 35992 31748
rect 36044 31736 36050 31748
rect 36081 31739 36139 31745
rect 36081 31736 36093 31739
rect 36044 31708 36093 31736
rect 36044 31696 36050 31708
rect 36081 31705 36093 31708
rect 36127 31705 36139 31739
rect 36188 31736 36216 31776
rect 36541 31773 36553 31807
rect 36587 31804 36599 31807
rect 36722 31804 36728 31816
rect 36587 31776 36728 31804
rect 36587 31773 36599 31776
rect 36541 31767 36599 31773
rect 36722 31764 36728 31776
rect 36780 31764 36786 31816
rect 37366 31764 37372 31816
rect 37424 31804 37430 31816
rect 37461 31807 37519 31813
rect 37461 31804 37473 31807
rect 37424 31776 37473 31804
rect 37424 31764 37430 31776
rect 37461 31773 37473 31776
rect 37507 31773 37519 31807
rect 37461 31767 37519 31773
rect 38473 31807 38531 31813
rect 38473 31773 38485 31807
rect 38519 31804 38531 31807
rect 51718 31804 51724 31816
rect 38519 31776 51724 31804
rect 38519 31773 38531 31776
rect 38473 31767 38531 31773
rect 38488 31736 38516 31767
rect 51718 31764 51724 31776
rect 51776 31764 51782 31816
rect 36188 31708 38516 31736
rect 36081 31699 36139 31705
rect 31018 31668 31024 31680
rect 30301 31640 31024 31668
rect 30193 31631 30251 31637
rect 31018 31628 31024 31640
rect 31076 31628 31082 31680
rect 31386 31628 31392 31680
rect 31444 31668 31450 31680
rect 32674 31668 32680 31680
rect 31444 31640 32680 31668
rect 31444 31628 31450 31640
rect 32674 31628 32680 31640
rect 32732 31668 32738 31680
rect 33410 31668 33416 31680
rect 32732 31640 33416 31668
rect 32732 31628 32738 31640
rect 33410 31628 33416 31640
rect 33468 31628 33474 31680
rect 37274 31668 37280 31680
rect 37235 31640 37280 31668
rect 37274 31628 37280 31640
rect 37332 31628 37338 31680
rect 1104 31578 54372 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 54372 31578
rect 1104 31504 54372 31526
rect 16022 31464 16028 31476
rect 15983 31436 16028 31464
rect 16022 31424 16028 31436
rect 16080 31424 16086 31476
rect 17681 31467 17739 31473
rect 17681 31433 17693 31467
rect 17727 31464 17739 31467
rect 18046 31464 18052 31476
rect 17727 31436 18052 31464
rect 17727 31433 17739 31436
rect 17681 31427 17739 31433
rect 18046 31424 18052 31436
rect 18104 31424 18110 31476
rect 18414 31424 18420 31476
rect 18472 31424 18478 31476
rect 22741 31467 22799 31473
rect 22741 31464 22753 31467
rect 22112 31436 22753 31464
rect 18432 31396 18460 31424
rect 18248 31368 18460 31396
rect 16942 31328 16948 31340
rect 16903 31300 16948 31328
rect 16942 31288 16948 31300
rect 17000 31288 17006 31340
rect 17129 31331 17187 31337
rect 17129 31297 17141 31331
rect 17175 31328 17187 31331
rect 17218 31328 17224 31340
rect 17175 31300 17224 31328
rect 17175 31297 17187 31300
rect 17129 31291 17187 31297
rect 17218 31288 17224 31300
rect 17276 31288 17282 31340
rect 17586 31328 17592 31340
rect 17547 31300 17592 31328
rect 17586 31288 17592 31300
rect 17644 31288 17650 31340
rect 17773 31331 17831 31337
rect 17773 31297 17785 31331
rect 17819 31328 17831 31331
rect 17954 31328 17960 31340
rect 17819 31300 17960 31328
rect 17819 31297 17831 31300
rect 17773 31291 17831 31297
rect 17954 31288 17960 31300
rect 18012 31288 18018 31340
rect 18248 31337 18276 31368
rect 18233 31331 18291 31337
rect 18233 31297 18245 31331
rect 18279 31297 18291 31331
rect 18396 31331 18454 31337
rect 18396 31328 18408 31331
rect 18233 31291 18291 31297
rect 18340 31300 18408 31328
rect 18340 31260 18368 31300
rect 18396 31297 18408 31300
rect 18442 31297 18454 31331
rect 18396 31291 18454 31297
rect 18506 31288 18512 31340
rect 18564 31328 18570 31340
rect 18690 31337 18696 31340
rect 18647 31331 18696 31337
rect 18564 31300 18609 31328
rect 18564 31288 18570 31300
rect 18647 31297 18659 31331
rect 18693 31297 18696 31331
rect 18647 31291 18696 31297
rect 18690 31288 18696 31291
rect 18748 31288 18754 31340
rect 19518 31328 19524 31340
rect 19479 31300 19524 31328
rect 19518 31288 19524 31300
rect 19576 31288 19582 31340
rect 20533 31331 20591 31337
rect 20533 31328 20545 31331
rect 19904 31300 20545 31328
rect 19610 31260 19616 31272
rect 16960 31232 18368 31260
rect 19571 31232 19616 31260
rect 16960 31136 16988 31232
rect 19610 31220 19616 31232
rect 19668 31220 19674 31272
rect 19904 31269 19932 31300
rect 20533 31297 20545 31300
rect 20579 31328 20591 31331
rect 20714 31328 20720 31340
rect 20579 31300 20720 31328
rect 20579 31297 20591 31300
rect 20533 31291 20591 31297
rect 20714 31288 20720 31300
rect 20772 31288 20778 31340
rect 22112 31337 22140 31436
rect 22741 31433 22753 31436
rect 22787 31464 22799 31467
rect 23474 31464 23480 31476
rect 22787 31436 23480 31464
rect 22787 31433 22799 31436
rect 22741 31427 22799 31433
rect 23474 31424 23480 31436
rect 23532 31424 23538 31476
rect 23661 31467 23719 31473
rect 23661 31433 23673 31467
rect 23707 31464 23719 31467
rect 23750 31464 23756 31476
rect 23707 31436 23756 31464
rect 23707 31433 23719 31436
rect 23661 31427 23719 31433
rect 23750 31424 23756 31436
rect 23808 31424 23814 31476
rect 25866 31424 25872 31476
rect 25924 31464 25930 31476
rect 25961 31467 26019 31473
rect 25961 31464 25973 31467
rect 25924 31436 25973 31464
rect 25924 31424 25930 31436
rect 25961 31433 25973 31436
rect 26007 31433 26019 31467
rect 32950 31464 32956 31476
rect 25961 31427 26019 31433
rect 31312 31436 32956 31464
rect 22646 31396 22652 31408
rect 22607 31368 22652 31396
rect 22646 31356 22652 31368
rect 22704 31356 22710 31408
rect 23569 31399 23627 31405
rect 23569 31365 23581 31399
rect 23615 31396 23627 31399
rect 24670 31396 24676 31408
rect 23615 31368 24676 31396
rect 23615 31365 23627 31368
rect 23569 31359 23627 31365
rect 24670 31356 24676 31368
rect 24728 31356 24734 31408
rect 21913 31331 21971 31337
rect 21913 31297 21925 31331
rect 21959 31297 21971 31331
rect 21913 31291 21971 31297
rect 22097 31331 22155 31337
rect 22097 31297 22109 31331
rect 22143 31297 22155 31331
rect 22554 31328 22560 31340
rect 22515 31300 22560 31328
rect 22097 31291 22155 31297
rect 19889 31263 19947 31269
rect 19889 31229 19901 31263
rect 19935 31229 19947 31263
rect 20438 31260 20444 31272
rect 20399 31232 20444 31260
rect 19889 31223 19947 31229
rect 20438 31220 20444 31232
rect 20496 31220 20502 31272
rect 21928 31260 21956 31291
rect 22554 31288 22560 31300
rect 22612 31288 22618 31340
rect 22833 31331 22891 31337
rect 22833 31297 22845 31331
rect 22879 31328 22891 31331
rect 23198 31328 23204 31340
rect 22879 31300 23204 31328
rect 22879 31297 22891 31300
rect 22833 31291 22891 31297
rect 23198 31288 23204 31300
rect 23256 31288 23262 31340
rect 23750 31328 23756 31340
rect 23711 31300 23756 31328
rect 23750 31288 23756 31300
rect 23808 31288 23814 31340
rect 24489 31331 24547 31337
rect 24489 31297 24501 31331
rect 24535 31297 24547 31331
rect 24489 31291 24547 31297
rect 25409 31331 25467 31337
rect 25409 31297 25421 31331
rect 25455 31328 25467 31331
rect 25498 31328 25504 31340
rect 25455 31300 25504 31328
rect 25455 31297 25467 31300
rect 25409 31291 25467 31297
rect 22186 31260 22192 31272
rect 21928 31232 22192 31260
rect 22186 31220 22192 31232
rect 22244 31260 22250 31272
rect 23293 31263 23351 31269
rect 23293 31260 23305 31263
rect 22244 31232 23305 31260
rect 22244 31220 22250 31232
rect 23293 31229 23305 31232
rect 23339 31229 23351 31263
rect 23293 31223 23351 31229
rect 23382 31220 23388 31272
rect 23440 31260 23446 31272
rect 24504 31260 24532 31291
rect 25498 31288 25504 31300
rect 25556 31288 25562 31340
rect 25682 31328 25688 31340
rect 25643 31300 25688 31328
rect 25682 31288 25688 31300
rect 25740 31288 25746 31340
rect 25774 31288 25780 31340
rect 25832 31328 25838 31340
rect 26970 31328 26976 31340
rect 25832 31300 25877 31328
rect 26931 31300 26976 31328
rect 25832 31288 25838 31300
rect 26970 31288 26976 31300
rect 27028 31288 27034 31340
rect 27246 31328 27252 31340
rect 27207 31300 27252 31328
rect 27246 31288 27252 31300
rect 27304 31288 27310 31340
rect 28902 31288 28908 31340
rect 28960 31328 28966 31340
rect 29365 31331 29423 31337
rect 29365 31328 29377 31331
rect 28960 31300 29377 31328
rect 28960 31288 28966 31300
rect 29365 31297 29377 31300
rect 29411 31297 29423 31331
rect 29546 31328 29552 31340
rect 29507 31300 29552 31328
rect 29365 31291 29423 31297
rect 23440 31232 24532 31260
rect 29380 31260 29408 31291
rect 29546 31288 29552 31300
rect 29604 31288 29610 31340
rect 31312 31337 31340 31436
rect 32950 31424 32956 31436
rect 33008 31424 33014 31476
rect 33781 31467 33839 31473
rect 33781 31433 33793 31467
rect 33827 31464 33839 31467
rect 33870 31464 33876 31476
rect 33827 31436 33876 31464
rect 33827 31433 33839 31436
rect 33781 31427 33839 31433
rect 33870 31424 33876 31436
rect 33928 31424 33934 31476
rect 35897 31467 35955 31473
rect 35897 31464 35909 31467
rect 34348 31436 35909 31464
rect 31573 31399 31631 31405
rect 31573 31365 31585 31399
rect 31619 31396 31631 31399
rect 34348 31396 34376 31436
rect 35897 31433 35909 31436
rect 35943 31433 35955 31467
rect 37642 31464 37648 31476
rect 37603 31436 37648 31464
rect 35897 31427 35955 31433
rect 37642 31424 37648 31436
rect 37700 31424 37706 31476
rect 31619 31368 31754 31396
rect 31619 31365 31631 31368
rect 31573 31359 31631 31365
rect 31297 31331 31355 31337
rect 31297 31297 31309 31331
rect 31343 31297 31355 31331
rect 31726 31328 31754 31368
rect 33152 31368 34376 31396
rect 33152 31340 33180 31368
rect 32125 31331 32183 31337
rect 32125 31328 32137 31331
rect 31726 31300 32137 31328
rect 31297 31291 31355 31297
rect 32125 31297 32137 31300
rect 32171 31297 32183 31331
rect 32125 31291 32183 31297
rect 32214 31288 32220 31340
rect 32272 31328 32278 31340
rect 32490 31328 32496 31340
rect 32272 31300 32317 31328
rect 32451 31300 32496 31328
rect 32272 31288 32278 31300
rect 32490 31288 32496 31300
rect 32548 31288 32554 31340
rect 33134 31328 33140 31340
rect 33047 31300 33140 31328
rect 33134 31288 33140 31300
rect 33192 31288 33198 31340
rect 34054 31328 34060 31340
rect 34015 31300 34060 31328
rect 34054 31288 34060 31300
rect 34112 31288 34118 31340
rect 34149 31331 34207 31337
rect 34149 31297 34161 31331
rect 34195 31297 34207 31331
rect 34149 31291 34207 31297
rect 34241 31331 34299 31337
rect 34241 31297 34253 31331
rect 34287 31328 34299 31331
rect 34348 31328 34376 31368
rect 35253 31399 35311 31405
rect 35253 31365 35265 31399
rect 35299 31396 35311 31399
rect 35710 31396 35716 31408
rect 35299 31368 35716 31396
rect 35299 31365 35311 31368
rect 35253 31359 35311 31365
rect 35710 31356 35716 31368
rect 35768 31356 35774 31408
rect 37274 31396 37280 31408
rect 36372 31368 37280 31396
rect 34287 31300 34376 31328
rect 34425 31331 34483 31337
rect 34287 31297 34299 31300
rect 34241 31291 34299 31297
rect 34425 31297 34437 31331
rect 34471 31297 34483 31331
rect 34425 31291 34483 31297
rect 35069 31331 35127 31337
rect 35069 31297 35081 31331
rect 35115 31328 35127 31331
rect 35434 31328 35440 31340
rect 35115 31300 35440 31328
rect 35115 31297 35127 31300
rect 35069 31291 35127 31297
rect 30009 31263 30067 31269
rect 30009 31260 30021 31263
rect 29380 31232 30021 31260
rect 23440 31220 23446 31232
rect 30009 31229 30021 31232
rect 30055 31229 30067 31263
rect 30009 31223 30067 31229
rect 31573 31263 31631 31269
rect 31573 31229 31585 31263
rect 31619 31260 31631 31263
rect 31846 31260 31852 31272
rect 31619 31232 31852 31260
rect 31619 31229 31631 31232
rect 31573 31223 31631 31229
rect 31846 31220 31852 31232
rect 31904 31220 31910 31272
rect 32309 31263 32367 31269
rect 32309 31229 32321 31263
rect 32355 31260 32367 31263
rect 32766 31260 32772 31272
rect 32355 31232 32772 31260
rect 32355 31229 32367 31232
rect 32309 31223 32367 31229
rect 20901 31195 20959 31201
rect 20901 31161 20913 31195
rect 20947 31192 20959 31195
rect 25501 31195 25559 31201
rect 25501 31192 25513 31195
rect 20947 31164 25513 31192
rect 20947 31161 20959 31164
rect 20901 31155 20959 31161
rect 25501 31161 25513 31164
rect 25547 31161 25559 31195
rect 25501 31155 25559 31161
rect 27982 31152 27988 31204
rect 28040 31192 28046 31204
rect 28040 31164 29960 31192
rect 28040 31152 28046 31164
rect 16942 31124 16948 31136
rect 16903 31096 16948 31124
rect 16942 31084 16948 31096
rect 17000 31084 17006 31136
rect 18874 31124 18880 31136
rect 18835 31096 18880 31124
rect 18874 31084 18880 31096
rect 18932 31084 18938 31136
rect 22002 31124 22008 31136
rect 21963 31096 22008 31124
rect 22002 31084 22008 31096
rect 22060 31084 22066 31136
rect 24029 31127 24087 31133
rect 24029 31093 24041 31127
rect 24075 31124 24087 31127
rect 24210 31124 24216 31136
rect 24075 31096 24216 31124
rect 24075 31093 24087 31096
rect 24029 31087 24087 31093
rect 24210 31084 24216 31096
rect 24268 31084 24274 31136
rect 24578 31124 24584 31136
rect 24539 31096 24584 31124
rect 24578 31084 24584 31096
rect 24636 31084 24642 31136
rect 28350 31124 28356 31136
rect 28311 31096 28356 31124
rect 28350 31084 28356 31096
rect 28408 31084 28414 31136
rect 29549 31127 29607 31133
rect 29549 31093 29561 31127
rect 29595 31124 29607 31127
rect 29822 31124 29828 31136
rect 29595 31096 29828 31124
rect 29595 31093 29607 31096
rect 29549 31087 29607 31093
rect 29822 31084 29828 31096
rect 29880 31084 29886 31136
rect 29932 31124 29960 31164
rect 30374 31152 30380 31204
rect 30432 31192 30438 31204
rect 30745 31195 30803 31201
rect 30745 31192 30757 31195
rect 30432 31164 30757 31192
rect 30432 31152 30438 31164
rect 30745 31161 30757 31164
rect 30791 31192 30803 31195
rect 30834 31192 30840 31204
rect 30791 31164 30840 31192
rect 30791 31161 30803 31164
rect 30745 31155 30803 31161
rect 30834 31152 30840 31164
rect 30892 31152 30898 31204
rect 31389 31195 31447 31201
rect 31389 31161 31401 31195
rect 31435 31192 31447 31195
rect 31754 31192 31760 31204
rect 31435 31164 31760 31192
rect 31435 31161 31447 31164
rect 31389 31155 31447 31161
rect 31754 31152 31760 31164
rect 31812 31192 31818 31204
rect 31938 31192 31944 31204
rect 31812 31164 31944 31192
rect 31812 31152 31818 31164
rect 31938 31152 31944 31164
rect 31996 31152 32002 31204
rect 32324 31124 32352 31223
rect 32766 31220 32772 31232
rect 32824 31220 32830 31272
rect 33321 31263 33379 31269
rect 33321 31229 33333 31263
rect 33367 31260 33379 31263
rect 33410 31260 33416 31272
rect 33367 31232 33416 31260
rect 33367 31229 33379 31232
rect 33321 31223 33379 31229
rect 33410 31220 33416 31232
rect 33468 31220 33474 31272
rect 33778 31220 33784 31272
rect 33836 31260 33842 31272
rect 34164 31260 34192 31291
rect 34440 31260 34468 31291
rect 35434 31288 35440 31300
rect 35492 31288 35498 31340
rect 36262 31328 36268 31340
rect 36223 31300 36268 31328
rect 36262 31288 36268 31300
rect 36320 31288 36326 31340
rect 34698 31260 34704 31272
rect 33836 31232 34192 31260
rect 34348 31232 34704 31260
rect 33836 31220 33842 31232
rect 33428 31192 33456 31220
rect 34348 31192 34376 31232
rect 34698 31220 34704 31232
rect 34756 31220 34762 31272
rect 36372 31269 36400 31368
rect 37274 31356 37280 31368
rect 37332 31356 37338 31408
rect 36538 31288 36544 31340
rect 36596 31328 36602 31340
rect 37737 31331 37795 31337
rect 37737 31328 37749 31331
rect 36596 31300 37749 31328
rect 36596 31288 36602 31300
rect 37737 31297 37749 31300
rect 37783 31297 37795 31331
rect 37737 31291 37795 31297
rect 36357 31263 36415 31269
rect 36357 31229 36369 31263
rect 36403 31229 36415 31263
rect 36357 31223 36415 31229
rect 37277 31263 37335 31269
rect 37277 31229 37289 31263
rect 37323 31229 37335 31263
rect 37277 31223 37335 31229
rect 33428 31164 34376 31192
rect 35437 31195 35495 31201
rect 35437 31161 35449 31195
rect 35483 31192 35495 31195
rect 36446 31192 36452 31204
rect 35483 31164 36452 31192
rect 35483 31161 35495 31164
rect 35437 31155 35495 31161
rect 36446 31152 36452 31164
rect 36504 31192 36510 31204
rect 37292 31192 37320 31223
rect 36504 31164 37320 31192
rect 36504 31152 36510 31164
rect 32490 31124 32496 31136
rect 29932 31096 32352 31124
rect 32451 31096 32496 31124
rect 32490 31084 32496 31096
rect 32548 31084 32554 31136
rect 32950 31124 32956 31136
rect 32911 31096 32956 31124
rect 32950 31084 32956 31096
rect 33008 31084 33014 31136
rect 36630 31084 36636 31136
rect 36688 31124 36694 31136
rect 37461 31127 37519 31133
rect 37461 31124 37473 31127
rect 36688 31096 37473 31124
rect 36688 31084 36694 31096
rect 37461 31093 37473 31096
rect 37507 31093 37519 31127
rect 38194 31124 38200 31136
rect 38155 31096 38200 31124
rect 37461 31087 37519 31093
rect 38194 31084 38200 31096
rect 38252 31084 38258 31136
rect 1104 31034 54372 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 54372 31034
rect 1104 30960 54372 30982
rect 21637 30923 21695 30929
rect 21637 30889 21649 30923
rect 21683 30920 21695 30923
rect 22186 30920 22192 30932
rect 21683 30892 22192 30920
rect 21683 30889 21695 30892
rect 21637 30883 21695 30889
rect 22186 30880 22192 30892
rect 22244 30880 22250 30932
rect 23385 30923 23443 30929
rect 23385 30889 23397 30923
rect 23431 30920 23443 30923
rect 23658 30920 23664 30932
rect 23431 30892 23664 30920
rect 23431 30889 23443 30892
rect 23385 30883 23443 30889
rect 23658 30880 23664 30892
rect 23716 30880 23722 30932
rect 25682 30880 25688 30932
rect 25740 30920 25746 30932
rect 25961 30923 26019 30929
rect 25961 30920 25973 30923
rect 25740 30892 25973 30920
rect 25740 30880 25746 30892
rect 25961 30889 25973 30892
rect 26007 30889 26019 30923
rect 25961 30883 26019 30889
rect 26050 30880 26056 30932
rect 26108 30920 26114 30932
rect 27249 30923 27307 30929
rect 26108 30892 26153 30920
rect 26108 30880 26114 30892
rect 27249 30889 27261 30923
rect 27295 30920 27307 30923
rect 27338 30920 27344 30932
rect 27295 30892 27344 30920
rect 27295 30889 27307 30892
rect 27249 30883 27307 30889
rect 18601 30855 18659 30861
rect 18601 30821 18613 30855
rect 18647 30852 18659 30855
rect 19610 30852 19616 30864
rect 18647 30824 19616 30852
rect 18647 30821 18659 30824
rect 18601 30815 18659 30821
rect 19610 30812 19616 30824
rect 19668 30852 19674 30864
rect 20993 30855 21051 30861
rect 20993 30852 21005 30855
rect 19668 30824 21005 30852
rect 19668 30812 19674 30824
rect 18322 30784 18328 30796
rect 18283 30756 18328 30784
rect 18322 30744 18328 30756
rect 18380 30744 18386 30796
rect 16942 30676 16948 30728
rect 17000 30716 17006 30728
rect 19904 30725 19932 30824
rect 20993 30821 21005 30824
rect 21039 30821 21051 30855
rect 20993 30815 21051 30821
rect 22741 30855 22799 30861
rect 22741 30821 22753 30855
rect 22787 30852 22799 30855
rect 25314 30852 25320 30864
rect 22787 30824 25320 30852
rect 22787 30821 22799 30824
rect 22741 30815 22799 30821
rect 25314 30812 25320 30824
rect 25372 30812 25378 30864
rect 20349 30787 20407 30793
rect 20349 30753 20361 30787
rect 20395 30784 20407 30787
rect 20809 30787 20867 30793
rect 20809 30784 20821 30787
rect 20395 30756 20821 30784
rect 20395 30753 20407 30756
rect 20349 30747 20407 30753
rect 20809 30753 20821 30756
rect 20855 30753 20867 30787
rect 20809 30747 20867 30753
rect 22002 30744 22008 30796
rect 22060 30784 22066 30796
rect 24673 30787 24731 30793
rect 24673 30784 24685 30787
rect 22060 30756 24685 30784
rect 22060 30744 22066 30756
rect 24673 30753 24685 30756
rect 24719 30753 24731 30787
rect 24673 30747 24731 30753
rect 24946 30744 24952 30796
rect 25004 30784 25010 30796
rect 25869 30787 25927 30793
rect 25869 30784 25881 30787
rect 25004 30756 25881 30784
rect 25004 30744 25010 30756
rect 25869 30753 25881 30756
rect 25915 30784 25927 30787
rect 27264 30784 27292 30883
rect 27338 30880 27344 30892
rect 27396 30920 27402 30932
rect 28261 30923 28319 30929
rect 28261 30920 28273 30923
rect 27396 30892 28273 30920
rect 27396 30880 27402 30892
rect 28261 30889 28273 30892
rect 28307 30889 28319 30923
rect 28261 30883 28319 30889
rect 31113 30923 31171 30929
rect 31113 30889 31125 30923
rect 31159 30920 31171 30923
rect 31202 30920 31208 30932
rect 31159 30892 31208 30920
rect 31159 30889 31171 30892
rect 31113 30883 31171 30889
rect 31202 30880 31208 30892
rect 31260 30880 31266 30932
rect 31938 30920 31944 30932
rect 31899 30892 31944 30920
rect 31938 30880 31944 30892
rect 31996 30880 32002 30932
rect 32214 30880 32220 30932
rect 32272 30920 32278 30932
rect 32309 30923 32367 30929
rect 32309 30920 32321 30923
rect 32272 30892 32321 30920
rect 32272 30880 32278 30892
rect 32309 30889 32321 30892
rect 32355 30889 32367 30923
rect 32766 30920 32772 30932
rect 32727 30892 32772 30920
rect 32309 30883 32367 30889
rect 32766 30880 32772 30892
rect 32824 30880 32830 30932
rect 34698 30920 34704 30932
rect 34659 30892 34704 30920
rect 34698 30880 34704 30892
rect 34756 30880 34762 30932
rect 35621 30923 35679 30929
rect 35621 30889 35633 30923
rect 35667 30920 35679 30923
rect 36078 30920 36084 30932
rect 35667 30892 36084 30920
rect 35667 30889 35679 30892
rect 35621 30883 35679 30889
rect 36078 30880 36084 30892
rect 36136 30920 36142 30932
rect 36538 30920 36544 30932
rect 36136 30892 36544 30920
rect 36136 30880 36142 30892
rect 36538 30880 36544 30892
rect 36596 30880 36602 30932
rect 37366 30852 37372 30864
rect 36464 30824 37372 30852
rect 25915 30756 27292 30784
rect 29549 30787 29607 30793
rect 25915 30753 25927 30756
rect 25869 30747 25927 30753
rect 29549 30753 29561 30787
rect 29595 30784 29607 30787
rect 32122 30784 32128 30796
rect 29595 30756 32128 30784
rect 29595 30753 29607 30756
rect 29549 30747 29607 30753
rect 32122 30744 32128 30756
rect 32180 30744 32186 30796
rect 33778 30784 33784 30796
rect 33739 30756 33784 30784
rect 33778 30744 33784 30756
rect 33836 30744 33842 30796
rect 36354 30784 36360 30796
rect 36315 30756 36360 30784
rect 36354 30744 36360 30756
rect 36412 30744 36418 30796
rect 36464 30793 36492 30824
rect 37366 30812 37372 30824
rect 37424 30812 37430 30864
rect 36449 30787 36507 30793
rect 36449 30753 36461 30787
rect 36495 30753 36507 30787
rect 36630 30784 36636 30796
rect 36591 30756 36636 30784
rect 36449 30747 36507 30753
rect 36630 30744 36636 30756
rect 36688 30744 36694 30796
rect 18233 30719 18291 30725
rect 18233 30716 18245 30719
rect 17000 30688 18245 30716
rect 17000 30676 17006 30688
rect 18233 30685 18245 30688
rect 18279 30685 18291 30719
rect 18233 30679 18291 30685
rect 19889 30719 19947 30725
rect 19889 30685 19901 30719
rect 19935 30685 19947 30719
rect 19889 30679 19947 30685
rect 20165 30719 20223 30725
rect 20165 30685 20177 30719
rect 20211 30716 20223 30719
rect 20254 30716 20260 30728
rect 20211 30688 20260 30716
rect 20211 30685 20223 30688
rect 20165 30679 20223 30685
rect 20254 30676 20260 30688
rect 20312 30676 20318 30728
rect 21085 30719 21143 30725
rect 21085 30685 21097 30719
rect 21131 30685 21143 30719
rect 21085 30679 21143 30685
rect 19429 30651 19487 30657
rect 19429 30617 19441 30651
rect 19475 30648 19487 30651
rect 19518 30648 19524 30660
rect 19475 30620 19524 30648
rect 19475 30617 19487 30620
rect 19429 30611 19487 30617
rect 19518 30608 19524 30620
rect 19576 30648 19582 30660
rect 19981 30651 20039 30657
rect 19981 30648 19993 30651
rect 19576 30620 19993 30648
rect 19576 30608 19582 30620
rect 19981 30617 19993 30620
rect 20027 30648 20039 30651
rect 21100 30648 21128 30679
rect 21358 30676 21364 30728
rect 21416 30716 21422 30728
rect 21545 30719 21603 30725
rect 21545 30716 21557 30719
rect 21416 30688 21557 30716
rect 21416 30676 21422 30688
rect 21545 30685 21557 30688
rect 21591 30685 21603 30719
rect 21545 30679 21603 30685
rect 21729 30719 21787 30725
rect 21729 30685 21741 30719
rect 21775 30685 21787 30719
rect 23198 30716 23204 30728
rect 23159 30688 23204 30716
rect 21729 30679 21787 30685
rect 21266 30648 21272 30660
rect 20027 30620 21272 30648
rect 20027 30617 20039 30620
rect 19981 30611 20039 30617
rect 21266 30608 21272 30620
rect 21324 30648 21330 30660
rect 21744 30648 21772 30679
rect 23198 30676 23204 30688
rect 23256 30676 23262 30728
rect 23477 30719 23535 30725
rect 23477 30685 23489 30719
rect 23523 30716 23535 30719
rect 23566 30716 23572 30728
rect 23523 30688 23572 30716
rect 23523 30685 23535 30688
rect 23477 30679 23535 30685
rect 23566 30676 23572 30688
rect 23624 30716 23630 30728
rect 24578 30716 24584 30728
rect 23624 30688 24584 30716
rect 23624 30676 23630 30688
rect 24578 30676 24584 30688
rect 24636 30676 24642 30728
rect 24762 30716 24768 30728
rect 24723 30688 24768 30716
rect 24762 30676 24768 30688
rect 24820 30676 24826 30728
rect 26142 30716 26148 30728
rect 26055 30688 26148 30716
rect 26142 30676 26148 30688
rect 26200 30716 26206 30728
rect 26697 30719 26755 30725
rect 26697 30716 26709 30719
rect 26200 30688 26709 30716
rect 26200 30676 26206 30688
rect 26697 30685 26709 30688
rect 26743 30716 26755 30719
rect 28350 30716 28356 30728
rect 26743 30688 28356 30716
rect 26743 30685 26755 30688
rect 26697 30679 26755 30685
rect 28350 30676 28356 30688
rect 28408 30676 28414 30728
rect 29822 30716 29828 30728
rect 29783 30688 29828 30716
rect 29822 30676 29828 30688
rect 29880 30676 29886 30728
rect 31846 30676 31852 30728
rect 31904 30716 31910 30728
rect 31941 30719 31999 30725
rect 31941 30716 31953 30719
rect 31904 30688 31953 30716
rect 31904 30676 31910 30688
rect 31941 30685 31953 30688
rect 31987 30685 31999 30719
rect 31941 30679 31999 30685
rect 32033 30719 32091 30725
rect 32033 30685 32045 30719
rect 32079 30716 32091 30719
rect 32950 30716 32956 30728
rect 32079 30688 32956 30716
rect 32079 30685 32091 30688
rect 32033 30679 32091 30685
rect 21324 30620 21772 30648
rect 21324 30608 21330 30620
rect 2130 30540 2136 30592
rect 2188 30580 2194 30592
rect 16945 30583 17003 30589
rect 16945 30580 16957 30583
rect 2188 30552 16957 30580
rect 2188 30540 2194 30552
rect 16945 30549 16957 30552
rect 16991 30580 17003 30583
rect 17497 30583 17555 30589
rect 17497 30580 17509 30583
rect 16991 30552 17509 30580
rect 16991 30549 17003 30552
rect 16945 30543 17003 30549
rect 17497 30549 17509 30552
rect 17543 30580 17555 30583
rect 17586 30580 17592 30592
rect 17543 30552 17592 30580
rect 17543 30549 17555 30552
rect 17497 30543 17555 30549
rect 17586 30540 17592 30552
rect 17644 30540 17650 30592
rect 20806 30580 20812 30592
rect 20767 30552 20812 30580
rect 20806 30540 20812 30552
rect 20864 30540 20870 30592
rect 21744 30580 21772 30620
rect 23293 30651 23351 30657
rect 23293 30617 23305 30651
rect 23339 30648 23351 30651
rect 23750 30648 23756 30660
rect 23339 30620 23756 30648
rect 23339 30617 23351 30620
rect 23293 30611 23351 30617
rect 23750 30608 23756 30620
rect 23808 30608 23814 30660
rect 26160 30648 26188 30676
rect 23860 30620 26188 30648
rect 31956 30648 31984 30679
rect 32950 30676 32956 30688
rect 33008 30676 33014 30728
rect 33689 30719 33747 30725
rect 33689 30685 33701 30719
rect 33735 30716 33747 30719
rect 34054 30716 34060 30728
rect 33735 30688 34060 30716
rect 33735 30685 33747 30688
rect 33689 30679 33747 30685
rect 34054 30676 34060 30688
rect 34112 30676 34118 30728
rect 35434 30676 35440 30728
rect 35492 30716 35498 30728
rect 35529 30719 35587 30725
rect 35529 30716 35541 30719
rect 35492 30688 35541 30716
rect 35492 30676 35498 30688
rect 35529 30685 35541 30688
rect 35575 30685 35587 30719
rect 35710 30716 35716 30728
rect 35671 30688 35716 30716
rect 35529 30679 35587 30685
rect 32858 30648 32864 30660
rect 31956 30620 32864 30648
rect 23860 30580 23888 30620
rect 32858 30608 32864 30620
rect 32916 30648 32922 30660
rect 35544 30648 35572 30679
rect 35710 30676 35716 30688
rect 35768 30676 35774 30728
rect 36541 30719 36599 30725
rect 36541 30685 36553 30719
rect 36587 30716 36599 30719
rect 37458 30716 37464 30728
rect 36587 30688 37464 30716
rect 36587 30685 36599 30688
rect 36541 30679 36599 30685
rect 37458 30676 37464 30688
rect 37516 30676 37522 30728
rect 37277 30651 37335 30657
rect 37277 30648 37289 30651
rect 32916 30620 33364 30648
rect 35544 30620 37289 30648
rect 32916 30608 32922 30620
rect 24394 30580 24400 30592
rect 21744 30552 23888 30580
rect 24355 30552 24400 30580
rect 24394 30540 24400 30552
rect 24452 30540 24458 30592
rect 27706 30580 27712 30592
rect 27667 30552 27712 30580
rect 27706 30540 27712 30552
rect 27764 30540 27770 30592
rect 33336 30589 33364 30620
rect 37277 30617 37289 30620
rect 37323 30648 37335 30651
rect 37737 30651 37795 30657
rect 37737 30648 37749 30651
rect 37323 30620 37749 30648
rect 37323 30617 37335 30620
rect 37277 30611 37335 30617
rect 37737 30617 37749 30620
rect 37783 30617 37795 30651
rect 37737 30611 37795 30617
rect 33321 30583 33379 30589
rect 33321 30549 33333 30583
rect 33367 30549 33379 30583
rect 36170 30580 36176 30592
rect 36131 30552 36176 30580
rect 33321 30543 33379 30549
rect 36170 30540 36176 30552
rect 36228 30540 36234 30592
rect 1104 30490 54372 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 54372 30490
rect 1104 30416 54372 30438
rect 23017 30379 23075 30385
rect 23017 30345 23029 30379
rect 23063 30376 23075 30379
rect 23382 30376 23388 30388
rect 23063 30348 23388 30376
rect 23063 30345 23075 30348
rect 23017 30339 23075 30345
rect 23382 30336 23388 30348
rect 23440 30336 23446 30388
rect 23753 30379 23811 30385
rect 23753 30345 23765 30379
rect 23799 30376 23811 30379
rect 24762 30376 24768 30388
rect 23799 30348 24768 30376
rect 23799 30345 23811 30348
rect 23753 30339 23811 30345
rect 24762 30336 24768 30348
rect 24820 30336 24826 30388
rect 25685 30379 25743 30385
rect 25685 30345 25697 30379
rect 25731 30376 25743 30379
rect 25774 30376 25780 30388
rect 25731 30348 25780 30376
rect 25731 30345 25743 30348
rect 25685 30339 25743 30345
rect 25774 30336 25780 30348
rect 25832 30336 25838 30388
rect 30650 30336 30656 30388
rect 30708 30376 30714 30388
rect 31018 30376 31024 30388
rect 30708 30348 31024 30376
rect 30708 30336 30714 30348
rect 31018 30336 31024 30348
rect 31076 30336 31082 30388
rect 33505 30379 33563 30385
rect 33505 30345 33517 30379
rect 33551 30376 33563 30379
rect 34054 30376 34060 30388
rect 33551 30348 34060 30376
rect 33551 30345 33563 30348
rect 33505 30339 33563 30345
rect 34054 30336 34060 30348
rect 34112 30336 34118 30388
rect 36262 30376 36268 30388
rect 36223 30348 36268 30376
rect 36262 30336 36268 30348
rect 36320 30336 36326 30388
rect 37369 30379 37427 30385
rect 37369 30345 37381 30379
rect 37415 30376 37427 30379
rect 38194 30376 38200 30388
rect 37415 30348 38200 30376
rect 37415 30345 37427 30348
rect 37369 30339 37427 30345
rect 38194 30336 38200 30348
rect 38252 30336 38258 30388
rect 18693 30311 18751 30317
rect 18693 30277 18705 30311
rect 18739 30308 18751 30311
rect 19245 30311 19303 30317
rect 19245 30308 19257 30311
rect 18739 30280 19257 30308
rect 18739 30277 18751 30280
rect 18693 30271 18751 30277
rect 19245 30277 19257 30280
rect 19291 30308 19303 30311
rect 19426 30308 19432 30320
rect 19291 30280 19432 30308
rect 19291 30277 19303 30280
rect 19245 30271 19303 30277
rect 19426 30268 19432 30280
rect 19484 30268 19490 30320
rect 20898 30268 20904 30320
rect 20956 30308 20962 30320
rect 21450 30308 21456 30320
rect 20956 30280 21456 30308
rect 20956 30268 20962 30280
rect 21450 30268 21456 30280
rect 21508 30308 21514 30320
rect 21913 30311 21971 30317
rect 21913 30308 21925 30311
rect 21508 30280 21925 30308
rect 21508 30268 21514 30280
rect 21913 30277 21925 30280
rect 21959 30277 21971 30311
rect 21913 30271 21971 30277
rect 23474 30268 23480 30320
rect 23532 30308 23538 30320
rect 24949 30311 25007 30317
rect 24949 30308 24961 30311
rect 23532 30280 24961 30308
rect 23532 30268 23538 30280
rect 24949 30277 24961 30280
rect 24995 30277 25007 30311
rect 24949 30271 25007 30277
rect 26050 30268 26056 30320
rect 26108 30268 26114 30320
rect 32392 30311 32450 30317
rect 32392 30277 32404 30311
rect 32438 30308 32450 30311
rect 32490 30308 32496 30320
rect 32438 30280 32496 30308
rect 32438 30277 32450 30280
rect 32392 30271 32450 30277
rect 32490 30268 32496 30280
rect 32548 30268 32554 30320
rect 47578 30308 47584 30320
rect 34900 30280 47584 30308
rect 20714 30200 20720 30252
rect 20772 30240 20778 30252
rect 20809 30243 20867 30249
rect 20809 30240 20821 30243
rect 20772 30212 20821 30240
rect 20772 30200 20778 30212
rect 20809 30209 20821 30212
rect 20855 30209 20867 30243
rect 20990 30240 20996 30252
rect 20951 30212 20996 30240
rect 20809 30203 20867 30209
rect 20990 30200 20996 30212
rect 21048 30200 21054 30252
rect 21818 30240 21824 30252
rect 21779 30212 21824 30240
rect 21818 30200 21824 30212
rect 21876 30200 21882 30252
rect 22005 30243 22063 30249
rect 22005 30209 22017 30243
rect 22051 30240 22063 30243
rect 22094 30240 22100 30252
rect 22051 30212 22100 30240
rect 22051 30209 22063 30212
rect 22005 30203 22063 30209
rect 22094 30200 22100 30212
rect 22152 30200 22158 30252
rect 22925 30243 22983 30249
rect 22925 30209 22937 30243
rect 22971 30209 22983 30243
rect 22925 30203 22983 30209
rect 23109 30243 23167 30249
rect 23109 30209 23121 30243
rect 23155 30240 23167 30243
rect 23382 30240 23388 30252
rect 23155 30212 23388 30240
rect 23155 30209 23167 30212
rect 23109 30203 23167 30209
rect 20254 30132 20260 30184
rect 20312 30172 20318 30184
rect 22940 30172 22968 30203
rect 23382 30200 23388 30212
rect 23440 30200 23446 30252
rect 23566 30240 23572 30252
rect 23527 30212 23572 30240
rect 23566 30200 23572 30212
rect 23624 30200 23630 30252
rect 23750 30240 23756 30252
rect 23711 30212 23756 30240
rect 23750 30200 23756 30212
rect 23808 30200 23814 30252
rect 24213 30243 24271 30249
rect 24213 30209 24225 30243
rect 24259 30209 24271 30243
rect 24394 30240 24400 30252
rect 24355 30212 24400 30240
rect 24213 30203 24271 30209
rect 23658 30172 23664 30184
rect 20312 30144 23664 30172
rect 20312 30132 20318 30144
rect 23658 30132 23664 30144
rect 23716 30172 23722 30184
rect 23934 30172 23940 30184
rect 23716 30144 23940 30172
rect 23716 30132 23722 30144
rect 23934 30132 23940 30144
rect 23992 30132 23998 30184
rect 24228 30104 24256 30203
rect 24394 30200 24400 30212
rect 24452 30200 24458 30252
rect 24854 30240 24860 30252
rect 24815 30212 24860 30240
rect 24854 30200 24860 30212
rect 24912 30200 24918 30252
rect 25225 30243 25283 30249
rect 25225 30209 25237 30243
rect 25271 30240 25283 30243
rect 25590 30240 25596 30252
rect 25271 30212 25596 30240
rect 25271 30209 25283 30212
rect 25225 30203 25283 30209
rect 25590 30200 25596 30212
rect 25648 30200 25654 30252
rect 25869 30243 25927 30249
rect 25869 30209 25881 30243
rect 25915 30240 25927 30243
rect 26068 30240 26096 30268
rect 26234 30240 26240 30252
rect 25915 30212 26240 30240
rect 25915 30209 25927 30212
rect 25869 30203 25927 30209
rect 26234 30200 26240 30212
rect 26292 30200 26298 30252
rect 26970 30240 26976 30252
rect 26931 30212 26976 30240
rect 26970 30200 26976 30212
rect 27028 30200 27034 30252
rect 28629 30243 28687 30249
rect 28629 30209 28641 30243
rect 28675 30240 28687 30243
rect 34900 30240 34928 30280
rect 47578 30268 47584 30280
rect 47636 30268 47642 30320
rect 28675 30212 34928 30240
rect 34977 30243 35035 30249
rect 28675 30209 28687 30212
rect 28629 30203 28687 30209
rect 34977 30209 34989 30243
rect 35023 30209 35035 30243
rect 35158 30240 35164 30252
rect 35119 30212 35164 30240
rect 34977 30203 35035 30209
rect 24305 30175 24363 30181
rect 24305 30141 24317 30175
rect 24351 30172 24363 30175
rect 25041 30175 25099 30181
rect 25041 30172 25053 30175
rect 24351 30144 25053 30172
rect 24351 30141 24363 30144
rect 24305 30135 24363 30141
rect 25041 30141 25053 30144
rect 25087 30141 25099 30175
rect 25314 30172 25320 30184
rect 25041 30135 25099 30141
rect 25148 30144 25320 30172
rect 25148 30104 25176 30144
rect 25314 30132 25320 30144
rect 25372 30132 25378 30184
rect 26053 30175 26111 30181
rect 26053 30141 26065 30175
rect 26099 30172 26111 30175
rect 26142 30172 26148 30184
rect 26099 30144 26148 30172
rect 26099 30141 26111 30144
rect 26053 30135 26111 30141
rect 26142 30132 26148 30144
rect 26200 30132 26206 30184
rect 27249 30175 27307 30181
rect 27249 30172 27261 30175
rect 26252 30144 27261 30172
rect 24228 30076 25176 30104
rect 25225 30107 25283 30113
rect 25225 30073 25237 30107
rect 25271 30104 25283 30107
rect 26252 30104 26280 30144
rect 27249 30141 27261 30144
rect 27295 30141 27307 30175
rect 27249 30135 27307 30141
rect 25271 30076 26280 30104
rect 25271 30073 25283 30076
rect 25225 30067 25283 30073
rect 17954 30036 17960 30048
rect 17915 30008 17960 30036
rect 17954 29996 17960 30008
rect 18012 29996 18018 30048
rect 19797 30039 19855 30045
rect 19797 30005 19809 30039
rect 19843 30036 19855 30039
rect 20346 30036 20352 30048
rect 19843 30008 20352 30036
rect 19843 30005 19855 30008
rect 19797 29999 19855 30005
rect 20346 29996 20352 30008
rect 20404 29996 20410 30048
rect 20901 30039 20959 30045
rect 20901 30005 20913 30039
rect 20947 30036 20959 30039
rect 22002 30036 22008 30048
rect 20947 30008 22008 30036
rect 20947 30005 20959 30008
rect 20901 29999 20959 30005
rect 22002 29996 22008 30008
rect 22060 29996 22066 30048
rect 26050 29996 26056 30048
rect 26108 30036 26114 30048
rect 28644 30036 28672 30203
rect 32122 30172 32128 30184
rect 32035 30144 32128 30172
rect 32122 30132 32128 30144
rect 32180 30132 32186 30184
rect 34992 30172 35020 30203
rect 35158 30200 35164 30212
rect 35216 30200 35222 30252
rect 35253 30243 35311 30249
rect 35253 30209 35265 30243
rect 35299 30240 35311 30243
rect 35710 30240 35716 30252
rect 35299 30212 35716 30240
rect 35299 30209 35311 30212
rect 35253 30203 35311 30209
rect 35710 30200 35716 30212
rect 35768 30200 35774 30252
rect 36078 30200 36084 30252
rect 36136 30240 36142 30252
rect 36173 30243 36231 30249
rect 36173 30240 36185 30243
rect 36136 30212 36185 30240
rect 36136 30200 36142 30212
rect 36173 30209 36185 30212
rect 36219 30209 36231 30243
rect 36173 30203 36231 30209
rect 36357 30243 36415 30249
rect 36357 30209 36369 30243
rect 36403 30240 36415 30243
rect 36446 30240 36452 30252
rect 36403 30212 36452 30240
rect 36403 30209 36415 30212
rect 36357 30203 36415 30209
rect 36446 30200 36452 30212
rect 36504 30200 36510 30252
rect 52917 30243 52975 30249
rect 52917 30209 52929 30243
rect 52963 30240 52975 30243
rect 53558 30240 53564 30252
rect 52963 30212 53564 30240
rect 52963 30209 52975 30212
rect 52917 30203 52975 30209
rect 53558 30200 53564 30212
rect 53616 30200 53622 30252
rect 35802 30172 35808 30184
rect 34992 30144 35808 30172
rect 35802 30132 35808 30144
rect 35860 30132 35866 30184
rect 26108 30008 28672 30036
rect 32140 30036 32168 30132
rect 32490 30036 32496 30048
rect 32140 30008 32496 30036
rect 26108 29996 26114 30008
rect 32490 29996 32496 30008
rect 32548 29996 32554 30048
rect 35253 30039 35311 30045
rect 35253 30005 35265 30039
rect 35299 30036 35311 30039
rect 35986 30036 35992 30048
rect 35299 30008 35992 30036
rect 35299 30005 35311 30008
rect 35253 29999 35311 30005
rect 35986 29996 35992 30008
rect 36044 30036 36050 30048
rect 36446 30036 36452 30048
rect 36044 30008 36452 30036
rect 36044 29996 36050 30008
rect 36446 29996 36452 30008
rect 36504 29996 36510 30048
rect 53466 30036 53472 30048
rect 53427 30008 53472 30036
rect 53466 29996 53472 30008
rect 53524 29996 53530 30048
rect 1104 29946 54372 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 54372 29946
rect 1104 29872 54372 29894
rect 18693 29835 18751 29841
rect 18693 29801 18705 29835
rect 18739 29832 18751 29835
rect 22922 29832 22928 29844
rect 18739 29804 22928 29832
rect 18739 29801 18751 29804
rect 18693 29795 18751 29801
rect 22922 29792 22928 29804
rect 22980 29832 22986 29844
rect 23198 29832 23204 29844
rect 22980 29804 23204 29832
rect 22980 29792 22986 29804
rect 23198 29792 23204 29804
rect 23256 29792 23262 29844
rect 23569 29835 23627 29841
rect 23569 29801 23581 29835
rect 23615 29832 23627 29835
rect 23750 29832 23756 29844
rect 23615 29804 23756 29832
rect 23615 29801 23627 29804
rect 23569 29795 23627 29801
rect 23750 29792 23756 29804
rect 23808 29792 23814 29844
rect 24854 29792 24860 29844
rect 24912 29832 24918 29844
rect 25133 29835 25191 29841
rect 25133 29832 25145 29835
rect 24912 29804 25145 29832
rect 24912 29792 24918 29804
rect 25133 29801 25145 29804
rect 25179 29801 25191 29835
rect 26142 29832 26148 29844
rect 26103 29804 26148 29832
rect 25133 29795 25191 29801
rect 26142 29792 26148 29804
rect 26200 29792 26206 29844
rect 30193 29835 30251 29841
rect 30193 29801 30205 29835
rect 30239 29832 30251 29835
rect 31202 29832 31208 29844
rect 30239 29804 31208 29832
rect 30239 29801 30251 29804
rect 30193 29795 30251 29801
rect 31202 29792 31208 29804
rect 31260 29792 31266 29844
rect 33042 29832 33048 29844
rect 33003 29804 33048 29832
rect 33042 29792 33048 29804
rect 33100 29792 33106 29844
rect 33318 29792 33324 29844
rect 33376 29832 33382 29844
rect 34057 29835 34115 29841
rect 34057 29832 34069 29835
rect 33376 29804 34069 29832
rect 33376 29792 33382 29804
rect 34057 29801 34069 29804
rect 34103 29832 34115 29835
rect 34146 29832 34152 29844
rect 34103 29804 34152 29832
rect 34103 29801 34115 29804
rect 34057 29795 34115 29801
rect 34146 29792 34152 29804
rect 34204 29792 34210 29844
rect 36446 29832 36452 29844
rect 36407 29804 36452 29832
rect 36446 29792 36452 29804
rect 36504 29792 36510 29844
rect 20346 29724 20352 29776
rect 20404 29764 20410 29776
rect 20717 29767 20775 29773
rect 20717 29764 20729 29767
rect 20404 29736 20729 29764
rect 20404 29724 20410 29736
rect 20717 29733 20729 29736
rect 20763 29764 20775 29767
rect 20898 29764 20904 29776
rect 20763 29736 20904 29764
rect 20763 29733 20775 29736
rect 20717 29727 20775 29733
rect 20898 29724 20904 29736
rect 20956 29764 20962 29776
rect 23017 29767 23075 29773
rect 20956 29736 22324 29764
rect 20956 29724 20962 29736
rect 20806 29656 20812 29708
rect 20864 29696 20870 29708
rect 21177 29699 21235 29705
rect 21177 29696 21189 29699
rect 20864 29668 21189 29696
rect 20864 29656 20870 29668
rect 21177 29665 21189 29668
rect 21223 29696 21235 29699
rect 21266 29696 21272 29708
rect 21223 29668 21272 29696
rect 21223 29665 21235 29668
rect 21177 29659 21235 29665
rect 21266 29656 21272 29668
rect 21324 29656 21330 29708
rect 22189 29699 22247 29705
rect 22189 29696 22201 29699
rect 21652 29668 22201 29696
rect 1394 29628 1400 29640
rect 1355 29600 1400 29628
rect 1394 29588 1400 29600
rect 1452 29588 1458 29640
rect 19242 29588 19248 29640
rect 19300 29628 19306 29640
rect 19613 29631 19671 29637
rect 19613 29628 19625 29631
rect 19300 29600 19625 29628
rect 19300 29588 19306 29600
rect 19613 29597 19625 29600
rect 19659 29597 19671 29631
rect 19613 29591 19671 29597
rect 19797 29631 19855 29637
rect 19797 29597 19809 29631
rect 19843 29628 19855 29631
rect 19978 29628 19984 29640
rect 19843 29600 19984 29628
rect 19843 29597 19855 29600
rect 19797 29591 19855 29597
rect 19978 29588 19984 29600
rect 20036 29588 20042 29640
rect 21450 29588 21456 29640
rect 21508 29628 21514 29640
rect 21652 29637 21680 29668
rect 22189 29665 22201 29668
rect 22235 29665 22247 29699
rect 22296 29696 22324 29736
rect 23017 29733 23029 29767
rect 23063 29764 23075 29767
rect 23290 29764 23296 29776
rect 23063 29736 23296 29764
rect 23063 29733 23075 29736
rect 23017 29727 23075 29733
rect 23290 29724 23296 29736
rect 23348 29724 23354 29776
rect 24489 29767 24547 29773
rect 24489 29733 24501 29767
rect 24535 29764 24547 29767
rect 24535 29736 25636 29764
rect 24535 29733 24547 29736
rect 24489 29727 24547 29733
rect 23382 29696 23388 29708
rect 22296 29668 23388 29696
rect 22189 29659 22247 29665
rect 23382 29656 23388 29668
rect 23440 29696 23446 29708
rect 24673 29699 24731 29705
rect 23440 29668 23704 29696
rect 23440 29656 23446 29668
rect 21545 29631 21603 29637
rect 21545 29628 21557 29631
rect 21508 29600 21557 29628
rect 21508 29588 21514 29600
rect 21545 29597 21557 29600
rect 21591 29597 21603 29631
rect 21545 29591 21603 29597
rect 21637 29631 21695 29637
rect 21637 29597 21649 29631
rect 21683 29597 21695 29631
rect 21637 29591 21695 29597
rect 22002 29588 22008 29640
rect 22060 29628 22066 29640
rect 22097 29631 22155 29637
rect 22097 29628 22109 29631
rect 22060 29600 22109 29628
rect 22060 29588 22066 29600
rect 22097 29597 22109 29600
rect 22143 29597 22155 29631
rect 22097 29591 22155 29597
rect 22741 29631 22799 29637
rect 22741 29597 22753 29631
rect 22787 29628 22799 29631
rect 23106 29628 23112 29640
rect 22787 29600 23112 29628
rect 22787 29597 22799 29600
rect 22741 29591 22799 29597
rect 20162 29560 20168 29572
rect 6886 29532 20168 29560
rect 1581 29495 1639 29501
rect 1581 29461 1593 29495
rect 1627 29492 1639 29495
rect 6886 29492 6914 29532
rect 20162 29520 20168 29532
rect 20220 29520 20226 29572
rect 22278 29560 22284 29572
rect 21468 29532 22284 29560
rect 18138 29492 18144 29504
rect 1627 29464 6914 29492
rect 18099 29464 18144 29492
rect 1627 29461 1639 29464
rect 1581 29455 1639 29461
rect 18138 29452 18144 29464
rect 18196 29452 18202 29504
rect 19334 29452 19340 29504
rect 19392 29492 19398 29504
rect 21468 29501 21496 29532
rect 22278 29520 22284 29532
rect 22336 29560 22342 29572
rect 22756 29560 22784 29591
rect 23106 29588 23112 29600
rect 23164 29588 23170 29640
rect 23676 29637 23704 29668
rect 24673 29665 24685 29699
rect 24719 29696 24731 29699
rect 24946 29696 24952 29708
rect 24719 29668 24952 29696
rect 24719 29665 24731 29668
rect 24673 29659 24731 29665
rect 24946 29656 24952 29668
rect 25004 29696 25010 29708
rect 25498 29696 25504 29708
rect 25004 29668 25504 29696
rect 25004 29656 25010 29668
rect 25498 29656 25504 29668
rect 25556 29656 25562 29708
rect 23477 29631 23535 29637
rect 23477 29597 23489 29631
rect 23523 29597 23535 29631
rect 23477 29591 23535 29597
rect 23661 29631 23719 29637
rect 23661 29597 23673 29631
rect 23707 29628 23719 29631
rect 23842 29628 23848 29640
rect 23707 29600 23848 29628
rect 23707 29597 23719 29600
rect 23661 29591 23719 29597
rect 22336 29532 22784 29560
rect 23017 29563 23075 29569
rect 22336 29520 22342 29532
rect 23017 29529 23029 29563
rect 23063 29560 23075 29563
rect 23198 29560 23204 29572
rect 23063 29532 23204 29560
rect 23063 29529 23075 29532
rect 23017 29523 23075 29529
rect 23198 29520 23204 29532
rect 23256 29520 23262 29572
rect 23492 29560 23520 29591
rect 23842 29588 23848 29600
rect 23900 29628 23906 29640
rect 25608 29637 25636 29736
rect 31662 29724 31668 29776
rect 31720 29764 31726 29776
rect 31720 29736 32076 29764
rect 31720 29724 31726 29736
rect 26605 29699 26663 29705
rect 26605 29665 26617 29699
rect 26651 29696 26663 29699
rect 26970 29696 26976 29708
rect 26651 29668 26976 29696
rect 26651 29665 26663 29668
rect 26605 29659 26663 29665
rect 26970 29656 26976 29668
rect 27028 29696 27034 29708
rect 27798 29696 27804 29708
rect 27028 29668 27804 29696
rect 27028 29656 27034 29668
rect 27798 29656 27804 29668
rect 27856 29656 27862 29708
rect 31478 29656 31484 29708
rect 31536 29696 31542 29708
rect 31941 29699 31999 29705
rect 31941 29696 31953 29699
rect 31536 29668 31953 29696
rect 31536 29656 31542 29668
rect 31941 29665 31953 29668
rect 31987 29665 31999 29699
rect 32048 29696 32076 29736
rect 32766 29724 32772 29776
rect 32824 29764 32830 29776
rect 53466 29764 53472 29776
rect 32824 29736 53472 29764
rect 32824 29724 32830 29736
rect 53466 29724 53472 29736
rect 53524 29724 53530 29776
rect 33318 29696 33324 29708
rect 32048 29668 33324 29696
rect 31941 29659 31999 29665
rect 33318 29656 33324 29668
rect 33376 29656 33382 29708
rect 33778 29656 33784 29708
rect 33836 29696 33842 29708
rect 34701 29699 34759 29705
rect 34701 29696 34713 29699
rect 33836 29668 34713 29696
rect 33836 29656 33842 29668
rect 34701 29665 34713 29668
rect 34747 29665 34759 29699
rect 36170 29696 36176 29708
rect 34701 29659 34759 29665
rect 35636 29668 36176 29696
rect 24397 29631 24455 29637
rect 24397 29628 24409 29631
rect 23900 29600 24409 29628
rect 23900 29588 23906 29600
rect 24397 29597 24409 29600
rect 24443 29597 24455 29631
rect 25317 29631 25375 29637
rect 25317 29628 25329 29631
rect 24397 29591 24455 29597
rect 24688 29600 25329 29628
rect 23750 29560 23756 29572
rect 23492 29532 23756 29560
rect 23750 29520 23756 29532
rect 23808 29520 23814 29572
rect 19705 29495 19763 29501
rect 19705 29492 19717 29495
rect 19392 29464 19717 29492
rect 19392 29452 19398 29464
rect 19705 29461 19717 29464
rect 19751 29461 19763 29495
rect 19705 29455 19763 29461
rect 21453 29495 21511 29501
rect 21453 29461 21465 29495
rect 21499 29461 21511 29495
rect 22830 29492 22836 29504
rect 22791 29464 22836 29492
rect 21453 29455 21511 29461
rect 22830 29452 22836 29464
rect 22888 29452 22894 29504
rect 24412 29492 24440 29591
rect 24688 29569 24716 29600
rect 25317 29597 25329 29600
rect 25363 29597 25375 29631
rect 25317 29591 25375 29597
rect 25593 29631 25651 29637
rect 25593 29597 25605 29631
rect 25639 29628 25651 29631
rect 25774 29628 25780 29640
rect 25639 29600 25780 29628
rect 25639 29597 25651 29600
rect 25593 29591 25651 29597
rect 25774 29588 25780 29600
rect 25832 29588 25838 29640
rect 26881 29631 26939 29637
rect 26881 29597 26893 29631
rect 26927 29628 26939 29631
rect 27246 29628 27252 29640
rect 26927 29600 27252 29628
rect 26927 29597 26939 29600
rect 26881 29591 26939 29597
rect 27246 29588 27252 29600
rect 27304 29588 27310 29640
rect 28810 29628 28816 29640
rect 28771 29600 28816 29628
rect 28810 29588 28816 29600
rect 28868 29588 28874 29640
rect 28997 29631 29055 29637
rect 28997 29597 29009 29631
rect 29043 29628 29055 29631
rect 29549 29631 29607 29637
rect 29549 29628 29561 29631
rect 29043 29600 29561 29628
rect 29043 29597 29055 29600
rect 28997 29591 29055 29597
rect 29549 29597 29561 29600
rect 29595 29628 29607 29631
rect 29822 29628 29828 29640
rect 29595 29600 29828 29628
rect 29595 29597 29607 29600
rect 29549 29591 29607 29597
rect 29822 29588 29828 29600
rect 29880 29588 29886 29640
rect 31662 29588 31668 29640
rect 31720 29630 31726 29640
rect 31720 29602 31763 29630
rect 31846 29628 31852 29640
rect 31720 29588 31726 29602
rect 31807 29600 31852 29628
rect 31846 29588 31852 29600
rect 31904 29588 31910 29640
rect 32033 29631 32091 29637
rect 32033 29597 32045 29631
rect 32079 29597 32091 29631
rect 32033 29591 32091 29597
rect 32217 29631 32275 29637
rect 32217 29597 32229 29631
rect 32263 29628 32275 29631
rect 32582 29628 32588 29640
rect 32263 29600 32588 29628
rect 32263 29597 32275 29600
rect 32217 29591 32275 29597
rect 24673 29563 24731 29569
rect 24673 29529 24685 29563
rect 24719 29529 24731 29563
rect 24673 29523 24731 29529
rect 25406 29492 25412 29504
rect 24412 29464 25412 29492
rect 25406 29452 25412 29464
rect 25464 29492 25470 29504
rect 25501 29495 25559 29501
rect 25501 29492 25513 29495
rect 25464 29464 25513 29492
rect 25464 29452 25470 29464
rect 25501 29461 25513 29464
rect 25547 29492 25559 29495
rect 26050 29492 26056 29504
rect 25547 29464 26056 29492
rect 25547 29461 25559 29464
rect 25501 29455 25559 29461
rect 26050 29452 26056 29464
rect 26108 29452 26114 29504
rect 27614 29452 27620 29504
rect 27672 29492 27678 29504
rect 27985 29495 28043 29501
rect 27985 29492 27997 29495
rect 27672 29464 27997 29492
rect 27672 29452 27678 29464
rect 27985 29461 27997 29464
rect 28031 29461 28043 29495
rect 27985 29455 28043 29461
rect 28997 29495 29055 29501
rect 28997 29461 29009 29495
rect 29043 29492 29055 29495
rect 29086 29492 29092 29504
rect 29043 29464 29092 29492
rect 29043 29461 29055 29464
rect 28997 29455 29055 29461
rect 29086 29452 29092 29464
rect 29144 29452 29150 29504
rect 30374 29452 30380 29504
rect 30432 29492 30438 29504
rect 30653 29495 30711 29501
rect 30653 29492 30665 29495
rect 30432 29464 30665 29492
rect 30432 29452 30438 29464
rect 30653 29461 30665 29464
rect 30699 29461 30711 29495
rect 30653 29455 30711 29461
rect 31386 29452 31392 29504
rect 31444 29492 31450 29504
rect 32048 29492 32076 29591
rect 32582 29588 32588 29600
rect 32640 29588 32646 29640
rect 32861 29631 32919 29637
rect 32861 29597 32873 29631
rect 32907 29597 32919 29631
rect 32861 29591 32919 29597
rect 33045 29631 33103 29637
rect 33045 29597 33057 29631
rect 33091 29628 33103 29631
rect 33134 29628 33140 29640
rect 33091 29600 33140 29628
rect 33091 29597 33103 29600
rect 33045 29591 33103 29597
rect 32876 29560 32904 29591
rect 33134 29588 33140 29600
rect 33192 29588 33198 29640
rect 35636 29614 35664 29668
rect 36170 29656 36176 29668
rect 36228 29656 36234 29708
rect 35710 29588 35716 29640
rect 35768 29628 35774 29640
rect 35768 29600 35813 29628
rect 35768 29588 35774 29600
rect 36630 29588 36636 29640
rect 36688 29628 36694 29640
rect 36725 29631 36783 29637
rect 36725 29628 36737 29631
rect 36688 29600 36737 29628
rect 36688 29588 36694 29600
rect 36725 29597 36737 29600
rect 36771 29597 36783 29631
rect 36725 29591 36783 29597
rect 33410 29560 33416 29572
rect 32876 29532 33416 29560
rect 33336 29504 33364 29532
rect 33410 29520 33416 29532
rect 33468 29520 33474 29572
rect 32398 29492 32404 29504
rect 31444 29464 32076 29492
rect 32359 29464 32404 29492
rect 31444 29452 31450 29464
rect 32398 29452 32404 29464
rect 32456 29452 32462 29504
rect 33318 29452 33324 29504
rect 33376 29492 33382 29504
rect 33505 29495 33563 29501
rect 33505 29492 33517 29495
rect 33376 29464 33517 29492
rect 33376 29452 33382 29464
rect 33505 29461 33517 29464
rect 33551 29461 33563 29495
rect 36262 29492 36268 29504
rect 36223 29464 36268 29492
rect 33505 29455 33563 29461
rect 36262 29452 36268 29464
rect 36320 29452 36326 29504
rect 1104 29402 54372 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 54372 29402
rect 1104 29328 54372 29350
rect 1394 29288 1400 29300
rect 1355 29260 1400 29288
rect 1394 29248 1400 29260
rect 1452 29248 1458 29300
rect 19242 29288 19248 29300
rect 19203 29260 19248 29288
rect 19242 29248 19248 29260
rect 19300 29248 19306 29300
rect 20717 29291 20775 29297
rect 20717 29257 20729 29291
rect 20763 29288 20775 29291
rect 20806 29288 20812 29300
rect 20763 29260 20812 29288
rect 20763 29257 20775 29260
rect 20717 29251 20775 29257
rect 20806 29248 20812 29260
rect 20864 29248 20870 29300
rect 21913 29291 21971 29297
rect 21913 29257 21925 29291
rect 21959 29288 21971 29291
rect 22094 29288 22100 29300
rect 21959 29260 22100 29288
rect 21959 29257 21971 29260
rect 21913 29251 21971 29257
rect 22094 29248 22100 29260
rect 22152 29248 22158 29300
rect 23293 29291 23351 29297
rect 23293 29257 23305 29291
rect 23339 29288 23351 29291
rect 23474 29288 23480 29300
rect 23339 29260 23480 29288
rect 23339 29257 23351 29260
rect 23293 29251 23351 29257
rect 23474 29248 23480 29260
rect 23532 29248 23538 29300
rect 23842 29288 23848 29300
rect 23803 29260 23848 29288
rect 23842 29248 23848 29260
rect 23900 29248 23906 29300
rect 33594 29288 33600 29300
rect 24136 29260 33600 29288
rect 18138 29220 18144 29232
rect 18051 29192 18144 29220
rect 18138 29180 18144 29192
rect 18196 29220 18202 29232
rect 20162 29220 20168 29232
rect 18196 29192 20168 29220
rect 18196 29180 18202 29192
rect 19352 29161 19380 29192
rect 20162 29180 20168 29192
rect 20220 29220 20226 29232
rect 24136 29220 24164 29260
rect 33594 29248 33600 29260
rect 33652 29248 33658 29300
rect 33781 29291 33839 29297
rect 33781 29257 33793 29291
rect 33827 29257 33839 29291
rect 33781 29251 33839 29257
rect 20220 29192 24164 29220
rect 25117 29223 25175 29229
rect 20220 29180 20226 29192
rect 25117 29189 25129 29223
rect 25163 29220 25175 29223
rect 25317 29223 25375 29229
rect 25163 29192 25268 29220
rect 25163 29189 25175 29192
rect 25117 29183 25175 29189
rect 19153 29155 19211 29161
rect 19153 29121 19165 29155
rect 19199 29121 19211 29155
rect 19153 29115 19211 29121
rect 19337 29155 19395 29161
rect 19337 29121 19349 29155
rect 19383 29121 19395 29155
rect 19337 29115 19395 29121
rect 19981 29155 20039 29161
rect 19981 29121 19993 29155
rect 20027 29152 20039 29155
rect 20254 29152 20260 29164
rect 20027 29124 20260 29152
rect 20027 29121 20039 29124
rect 19981 29115 20039 29121
rect 17589 29087 17647 29093
rect 17589 29053 17601 29087
rect 17635 29084 17647 29087
rect 19168 29084 19196 29115
rect 19996 29084 20024 29115
rect 20254 29112 20260 29124
rect 20312 29112 20318 29164
rect 20625 29155 20683 29161
rect 20625 29121 20637 29155
rect 20671 29121 20683 29155
rect 20898 29152 20904 29164
rect 20859 29124 20904 29152
rect 20625 29115 20683 29121
rect 17635 29056 20024 29084
rect 20640 29084 20668 29115
rect 20898 29112 20904 29124
rect 20956 29112 20962 29164
rect 21726 29112 21732 29164
rect 21784 29152 21790 29164
rect 21821 29155 21879 29161
rect 21821 29152 21833 29155
rect 21784 29124 21833 29152
rect 21784 29112 21790 29124
rect 21821 29121 21833 29124
rect 21867 29121 21879 29155
rect 21821 29115 21879 29121
rect 22094 29112 22100 29164
rect 22152 29152 22158 29164
rect 22830 29152 22836 29164
rect 22152 29124 22836 29152
rect 22152 29112 22158 29124
rect 22830 29112 22836 29124
rect 22888 29152 22894 29164
rect 23017 29155 23075 29161
rect 23017 29152 23029 29155
rect 22888 29124 23029 29152
rect 22888 29112 22894 29124
rect 23017 29121 23029 29124
rect 23063 29121 23075 29155
rect 23017 29115 23075 29121
rect 23106 29112 23112 29164
rect 23164 29152 23170 29164
rect 25240 29152 25268 29192
rect 25317 29189 25329 29223
rect 25363 29220 25375 29223
rect 25406 29220 25412 29232
rect 25363 29192 25412 29220
rect 25363 29189 25375 29192
rect 25317 29183 25375 29189
rect 25406 29180 25412 29192
rect 25464 29180 25470 29232
rect 26234 29220 26240 29232
rect 25884 29192 26240 29220
rect 25774 29152 25780 29164
rect 23164 29124 23209 29152
rect 25240 29124 25780 29152
rect 23164 29112 23170 29124
rect 25774 29112 25780 29124
rect 25832 29112 25838 29164
rect 25884 29152 25912 29192
rect 26234 29180 26240 29192
rect 26292 29180 26298 29232
rect 31570 29220 31576 29232
rect 31220 29192 31576 29220
rect 25953 29155 26011 29161
rect 25953 29152 25965 29155
rect 25884 29124 25965 29152
rect 25953 29121 25965 29124
rect 25999 29121 26011 29155
rect 25953 29115 26011 29121
rect 26050 29112 26056 29164
rect 26108 29152 26114 29164
rect 26973 29155 27031 29161
rect 26108 29124 26153 29152
rect 26108 29112 26114 29124
rect 26973 29121 26985 29155
rect 27019 29121 27031 29155
rect 26973 29115 27031 29121
rect 27157 29155 27215 29161
rect 27157 29121 27169 29155
rect 27203 29152 27215 29155
rect 27203 29124 27476 29152
rect 27203 29121 27215 29124
rect 27157 29115 27215 29121
rect 23290 29084 23296 29096
rect 20640 29056 20760 29084
rect 23251 29056 23296 29084
rect 17635 29053 17647 29056
rect 17589 29047 17647 29053
rect 20732 29028 20760 29056
rect 23290 29044 23296 29056
rect 23348 29044 23354 29096
rect 24489 29087 24547 29093
rect 24489 29053 24501 29087
rect 24535 29084 24547 29087
rect 26142 29084 26148 29096
rect 24535 29056 26148 29084
rect 24535 29053 24547 29056
rect 24489 29047 24547 29053
rect 26142 29044 26148 29056
rect 26200 29044 26206 29096
rect 26237 29087 26295 29093
rect 26237 29053 26249 29087
rect 26283 29084 26295 29087
rect 26326 29084 26332 29096
rect 26283 29056 26332 29084
rect 26283 29053 26295 29056
rect 26237 29047 26295 29053
rect 26326 29044 26332 29056
rect 26384 29044 26390 29096
rect 18693 29019 18751 29025
rect 18693 28985 18705 29019
rect 18739 29016 18751 29019
rect 20346 29016 20352 29028
rect 18739 28988 20352 29016
rect 18739 28985 18751 28988
rect 18693 28979 18751 28985
rect 20346 28976 20352 28988
rect 20404 28976 20410 29028
rect 20714 28976 20720 29028
rect 20772 28976 20778 29028
rect 22002 28976 22008 29028
rect 22060 29016 22066 29028
rect 22189 29019 22247 29025
rect 22189 29016 22201 29019
rect 22060 28988 22201 29016
rect 22060 28976 22066 28988
rect 22189 28985 22201 28988
rect 22235 28985 22247 29019
rect 22189 28979 22247 28985
rect 24854 28976 24860 29028
rect 24912 29016 24918 29028
rect 26988 29016 27016 29115
rect 27448 29028 27476 29124
rect 27798 29112 27804 29164
rect 27856 29152 27862 29164
rect 28445 29155 28503 29161
rect 28445 29152 28457 29155
rect 27856 29124 28457 29152
rect 27856 29112 27862 29124
rect 28445 29121 28457 29124
rect 28491 29121 28503 29155
rect 28445 29115 28503 29121
rect 28534 29112 28540 29164
rect 28592 29152 28598 29164
rect 31220 29161 31248 29192
rect 31570 29180 31576 29192
rect 31628 29180 31634 29232
rect 33796 29220 33824 29251
rect 33870 29248 33876 29300
rect 33928 29288 33934 29300
rect 53374 29288 53380 29300
rect 33928 29260 53380 29288
rect 33928 29248 33934 29260
rect 53374 29248 53380 29260
rect 53432 29248 53438 29300
rect 33796 29192 34928 29220
rect 28701 29155 28759 29161
rect 28701 29152 28713 29155
rect 28592 29124 28713 29152
rect 28592 29112 28598 29124
rect 28701 29121 28713 29124
rect 28747 29121 28759 29155
rect 28701 29115 28759 29121
rect 30745 29155 30803 29161
rect 30745 29121 30757 29155
rect 30791 29152 30803 29155
rect 31205 29155 31263 29161
rect 31205 29152 31217 29155
rect 30791 29124 31217 29152
rect 30791 29121 30803 29124
rect 30745 29115 30803 29121
rect 31205 29121 31217 29124
rect 31251 29121 31263 29155
rect 31205 29115 31263 29121
rect 31294 29112 31300 29164
rect 31352 29152 31358 29164
rect 31389 29155 31447 29161
rect 31389 29152 31401 29155
rect 31352 29124 31401 29152
rect 31352 29112 31358 29124
rect 31389 29121 31401 29124
rect 31435 29121 31447 29155
rect 31389 29115 31447 29121
rect 32030 29112 32036 29164
rect 32088 29152 32094 29164
rect 32125 29155 32183 29161
rect 32125 29152 32137 29155
rect 32088 29124 32137 29152
rect 32088 29112 32094 29124
rect 32125 29121 32137 29124
rect 32171 29121 32183 29155
rect 32125 29115 32183 29121
rect 32582 29112 32588 29164
rect 32640 29152 32646 29164
rect 34900 29161 34928 29192
rect 32677 29155 32735 29161
rect 32677 29152 32689 29155
rect 32640 29124 32689 29152
rect 32640 29112 32646 29124
rect 32677 29121 32689 29124
rect 32723 29121 32735 29155
rect 33587 29155 33645 29161
rect 33587 29152 33599 29155
rect 32677 29115 32735 29121
rect 33520 29124 33599 29152
rect 24912 28988 25912 29016
rect 24912 28976 24918 28988
rect 19794 28948 19800 28960
rect 19755 28920 19800 28948
rect 19794 28908 19800 28920
rect 19852 28908 19858 28960
rect 20898 28948 20904 28960
rect 20859 28920 20904 28948
rect 20898 28908 20904 28920
rect 20956 28908 20962 28960
rect 22281 28951 22339 28957
rect 22281 28917 22293 28951
rect 22327 28948 22339 28951
rect 22370 28948 22376 28960
rect 22327 28920 22376 28948
rect 22327 28917 22339 28920
rect 22281 28911 22339 28917
rect 22370 28908 22376 28920
rect 22428 28908 22434 28960
rect 22554 28948 22560 28960
rect 22515 28920 22560 28948
rect 22554 28908 22560 28920
rect 22612 28908 22618 28960
rect 24946 28948 24952 28960
rect 24907 28920 24952 28948
rect 24946 28908 24952 28920
rect 25004 28908 25010 28960
rect 25130 28948 25136 28960
rect 25091 28920 25136 28948
rect 25130 28908 25136 28920
rect 25188 28908 25194 28960
rect 25498 28908 25504 28960
rect 25556 28948 25562 28960
rect 25777 28951 25835 28957
rect 25777 28948 25789 28951
rect 25556 28920 25789 28948
rect 25556 28908 25562 28920
rect 25777 28917 25789 28920
rect 25823 28917 25835 28951
rect 25884 28948 25912 28988
rect 26160 28988 27016 29016
rect 26160 28948 26188 28988
rect 27430 28976 27436 29028
rect 27488 29016 27494 29028
rect 27617 29019 27675 29025
rect 27617 29016 27629 29019
rect 27488 28988 27629 29016
rect 27488 28976 27494 28988
rect 27617 28985 27629 28988
rect 27663 29016 27675 29019
rect 27706 29016 27712 29028
rect 27663 28988 27712 29016
rect 27663 28985 27675 28988
rect 27617 28979 27675 28985
rect 27706 28976 27712 28988
rect 27764 28976 27770 29028
rect 29638 29016 29644 29028
rect 29380 28988 29644 29016
rect 26970 28948 26976 28960
rect 25884 28920 26188 28948
rect 26931 28920 26976 28948
rect 25777 28911 25835 28917
rect 26970 28908 26976 28920
rect 27028 28908 27034 28960
rect 28718 28908 28724 28960
rect 28776 28948 28782 28960
rect 29380 28948 29408 28988
rect 29638 28976 29644 28988
rect 29696 29016 29702 29028
rect 29822 29016 29828 29028
rect 29696 28988 29828 29016
rect 29696 28976 29702 28988
rect 29822 28976 29828 28988
rect 29880 28976 29886 29028
rect 31294 28976 31300 29028
rect 31352 29016 31358 29028
rect 31481 29019 31539 29025
rect 31481 29016 31493 29019
rect 31352 28988 31493 29016
rect 31352 28976 31358 28988
rect 31481 28985 31493 28988
rect 31527 28985 31539 29019
rect 33520 29016 33548 29124
rect 33587 29121 33599 29124
rect 33633 29121 33645 29155
rect 33587 29115 33645 29121
rect 33781 29155 33839 29161
rect 33781 29121 33793 29155
rect 33827 29152 33839 29155
rect 34885 29155 34943 29161
rect 33827 29124 34836 29152
rect 33827 29121 33839 29124
rect 33781 29115 33839 29121
rect 34333 29087 34391 29093
rect 34333 29053 34345 29087
rect 34379 29084 34391 29087
rect 34422 29084 34428 29096
rect 34379 29056 34428 29084
rect 34379 29053 34391 29056
rect 34333 29047 34391 29053
rect 34422 29044 34428 29056
rect 34480 29044 34486 29096
rect 34808 29084 34836 29124
rect 34885 29121 34897 29155
rect 34931 29121 34943 29155
rect 34885 29115 34943 29121
rect 35253 29155 35311 29161
rect 35253 29121 35265 29155
rect 35299 29152 35311 29155
rect 35805 29155 35863 29161
rect 35805 29152 35817 29155
rect 35299 29124 35817 29152
rect 35299 29121 35311 29124
rect 35253 29115 35311 29121
rect 35805 29121 35817 29124
rect 35851 29121 35863 29155
rect 35805 29115 35863 29121
rect 35989 29155 36047 29161
rect 35989 29121 36001 29155
rect 36035 29152 36047 29155
rect 36170 29152 36176 29164
rect 36035 29124 36176 29152
rect 36035 29121 36047 29124
rect 35989 29115 36047 29121
rect 36170 29112 36176 29124
rect 36228 29112 36234 29164
rect 35342 29084 35348 29096
rect 34808 29056 35348 29084
rect 35342 29044 35348 29056
rect 35400 29044 35406 29096
rect 35618 29044 35624 29096
rect 35676 29084 35682 29096
rect 36081 29087 36139 29093
rect 36081 29084 36093 29087
rect 35676 29056 36093 29084
rect 35676 29044 35682 29056
rect 36081 29053 36093 29056
rect 36127 29053 36139 29087
rect 36446 29084 36452 29096
rect 36407 29056 36452 29084
rect 36081 29047 36139 29053
rect 36446 29044 36452 29056
rect 36504 29044 36510 29096
rect 35802 29016 35808 29028
rect 33520 28988 35808 29016
rect 31481 28979 31539 28985
rect 35802 28976 35808 28988
rect 35860 28976 35866 29028
rect 28776 28920 29408 28948
rect 28776 28908 28782 28920
rect 30650 28908 30656 28960
rect 30708 28948 30714 28960
rect 31938 28948 31944 28960
rect 30708 28920 31944 28948
rect 30708 28908 30714 28920
rect 31938 28908 31944 28920
rect 31996 28908 32002 28960
rect 32217 28951 32275 28957
rect 32217 28917 32229 28951
rect 32263 28948 32275 28951
rect 33962 28948 33968 28960
rect 32263 28920 33968 28948
rect 32263 28917 32275 28920
rect 32217 28911 32275 28917
rect 33962 28908 33968 28920
rect 34020 28908 34026 28960
rect 1104 28858 54372 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 54372 28858
rect 1104 28784 54372 28806
rect 18509 28747 18567 28753
rect 18509 28713 18521 28747
rect 18555 28744 18567 28747
rect 18874 28744 18880 28756
rect 18555 28716 18880 28744
rect 18555 28713 18567 28716
rect 18509 28707 18567 28713
rect 18874 28704 18880 28716
rect 18932 28744 18938 28756
rect 19426 28744 19432 28756
rect 18932 28716 19432 28744
rect 18932 28704 18938 28716
rect 19426 28704 19432 28716
rect 19484 28704 19490 28756
rect 21266 28744 21272 28756
rect 19536 28716 20116 28744
rect 21227 28716 21272 28744
rect 18782 28636 18788 28688
rect 18840 28676 18846 28688
rect 19536 28676 19564 28716
rect 18840 28648 19564 28676
rect 19705 28679 19763 28685
rect 18840 28636 18846 28648
rect 19705 28645 19717 28679
rect 19751 28676 19763 28679
rect 19978 28676 19984 28688
rect 19751 28648 19984 28676
rect 19751 28645 19763 28648
rect 19705 28639 19763 28645
rect 19978 28636 19984 28648
rect 20036 28636 20042 28688
rect 20088 28676 20116 28716
rect 21266 28704 21272 28716
rect 21324 28704 21330 28756
rect 28261 28747 28319 28753
rect 22066 28716 27844 28744
rect 22066 28676 22094 28716
rect 20088 28648 22094 28676
rect 23658 28636 23664 28688
rect 23716 28676 23722 28688
rect 25130 28676 25136 28688
rect 23716 28648 25136 28676
rect 23716 28636 23722 28648
rect 18693 28611 18751 28617
rect 18693 28577 18705 28611
rect 18739 28608 18751 28611
rect 19334 28608 19340 28620
rect 18739 28580 19340 28608
rect 18739 28577 18751 28580
rect 18693 28571 18751 28577
rect 19334 28568 19340 28580
rect 19392 28568 19398 28620
rect 20070 28608 20076 28620
rect 19536 28580 20076 28608
rect 17218 28500 17224 28552
rect 17276 28540 17282 28552
rect 19536 28549 19564 28580
rect 20070 28568 20076 28580
rect 20128 28568 20134 28620
rect 20441 28611 20499 28617
rect 20441 28577 20453 28611
rect 20487 28608 20499 28611
rect 21361 28611 21419 28617
rect 21361 28608 21373 28611
rect 20487 28580 21373 28608
rect 20487 28577 20499 28580
rect 20441 28571 20499 28577
rect 21361 28577 21373 28580
rect 21407 28577 21419 28611
rect 21361 28571 21419 28577
rect 18417 28543 18475 28549
rect 18417 28540 18429 28543
rect 17276 28512 18429 28540
rect 17276 28500 17282 28512
rect 18417 28509 18429 28512
rect 18463 28540 18475 28543
rect 19521 28543 19579 28549
rect 19521 28540 19533 28543
rect 18463 28512 19533 28540
rect 18463 28509 18475 28512
rect 18417 28503 18475 28509
rect 19521 28509 19533 28512
rect 19567 28509 19579 28543
rect 19521 28503 19579 28509
rect 19610 28500 19616 28552
rect 19668 28540 19674 28552
rect 19668 28512 19713 28540
rect 19668 28500 19674 28512
rect 19794 28500 19800 28552
rect 19852 28540 19858 28552
rect 20809 28543 20867 28549
rect 19852 28512 19897 28540
rect 19852 28500 19858 28512
rect 20809 28509 20821 28543
rect 20855 28540 20867 28543
rect 20898 28540 20904 28552
rect 20855 28512 20904 28540
rect 20855 28509 20867 28512
rect 20809 28503 20867 28509
rect 20898 28500 20904 28512
rect 20956 28500 20962 28552
rect 21266 28540 21272 28552
rect 21227 28512 21272 28540
rect 21266 28500 21272 28512
rect 21324 28500 21330 28552
rect 21376 28540 21404 28571
rect 22094 28540 22100 28552
rect 21376 28512 22100 28540
rect 22094 28500 22100 28512
rect 22152 28540 22158 28552
rect 22152 28512 22197 28540
rect 22152 28500 22158 28512
rect 22278 28500 22284 28552
rect 22336 28540 22342 28552
rect 22557 28543 22615 28549
rect 22336 28512 22381 28540
rect 22336 28500 22342 28512
rect 22557 28509 22569 28543
rect 22603 28509 22615 28543
rect 22557 28503 22615 28509
rect 18693 28475 18751 28481
rect 18693 28441 18705 28475
rect 18739 28472 18751 28475
rect 20625 28475 20683 28481
rect 18739 28444 20300 28472
rect 18739 28441 18751 28444
rect 18693 28435 18751 28441
rect 19334 28404 19340 28416
rect 19295 28376 19340 28404
rect 19334 28364 19340 28376
rect 19392 28364 19398 28416
rect 20272 28404 20300 28444
rect 20625 28441 20637 28475
rect 20671 28472 20683 28475
rect 22002 28472 22008 28484
rect 20671 28444 22008 28472
rect 20671 28441 20683 28444
rect 20625 28435 20683 28441
rect 22002 28432 22008 28444
rect 22060 28472 22066 28484
rect 22572 28472 22600 28503
rect 22060 28444 22600 28472
rect 22741 28475 22799 28481
rect 22060 28432 22066 28444
rect 22741 28441 22753 28475
rect 22787 28472 22799 28475
rect 23106 28472 23112 28484
rect 22787 28444 23112 28472
rect 22787 28441 22799 28444
rect 22741 28435 22799 28441
rect 23106 28432 23112 28444
rect 23164 28472 23170 28484
rect 23201 28475 23259 28481
rect 23201 28472 23213 28475
rect 23164 28444 23213 28472
rect 23164 28432 23170 28444
rect 23201 28441 23213 28444
rect 23247 28441 23259 28475
rect 23382 28472 23388 28484
rect 23343 28444 23388 28472
rect 23201 28435 23259 28441
rect 23382 28432 23388 28444
rect 23440 28432 23446 28484
rect 20806 28404 20812 28416
rect 20272 28376 20812 28404
rect 20806 28364 20812 28376
rect 20864 28364 20870 28416
rect 21637 28407 21695 28413
rect 21637 28373 21649 28407
rect 21683 28404 21695 28407
rect 22646 28404 22652 28416
rect 21683 28376 22652 28404
rect 21683 28373 21695 28376
rect 21637 28367 21695 28373
rect 22646 28364 22652 28376
rect 22704 28364 22710 28416
rect 23569 28407 23627 28413
rect 23569 28373 23581 28407
rect 23615 28404 23627 28407
rect 23934 28404 23940 28416
rect 23615 28376 23940 28404
rect 23615 28373 23627 28376
rect 23569 28367 23627 28373
rect 23934 28364 23940 28376
rect 23992 28364 23998 28416
rect 24118 28364 24124 28416
rect 24176 28404 24182 28416
rect 24857 28407 24915 28413
rect 24857 28404 24869 28407
rect 24176 28376 24869 28404
rect 24176 28364 24182 28376
rect 24857 28373 24869 28376
rect 24903 28373 24915 28407
rect 24964 28404 24992 28648
rect 25130 28636 25136 28648
rect 25188 28636 25194 28688
rect 25314 28676 25320 28688
rect 25240 28648 25320 28676
rect 25240 28617 25268 28648
rect 25314 28636 25320 28648
rect 25372 28636 25378 28688
rect 27816 28676 27844 28716
rect 28261 28713 28273 28747
rect 28307 28744 28319 28747
rect 28534 28744 28540 28756
rect 28307 28716 28540 28744
rect 28307 28713 28319 28716
rect 28261 28707 28319 28713
rect 28534 28704 28540 28716
rect 28592 28704 28598 28756
rect 30469 28747 30527 28753
rect 28644 28716 30420 28744
rect 28644 28676 28672 28716
rect 29549 28679 29607 28685
rect 29549 28676 29561 28679
rect 27816 28648 28672 28676
rect 28736 28648 29561 28676
rect 25041 28611 25099 28617
rect 25041 28577 25053 28611
rect 25087 28577 25099 28611
rect 25041 28571 25099 28577
rect 25225 28611 25283 28617
rect 25225 28577 25237 28611
rect 25271 28577 25283 28611
rect 27798 28608 27804 28620
rect 27759 28580 27804 28608
rect 25225 28571 25283 28577
rect 25056 28472 25084 28571
rect 27798 28568 27804 28580
rect 27856 28568 27862 28620
rect 28736 28617 28764 28648
rect 29549 28645 29561 28648
rect 29595 28645 29607 28679
rect 29549 28639 29607 28645
rect 28721 28611 28779 28617
rect 28721 28577 28733 28611
rect 28767 28577 28779 28611
rect 28721 28571 28779 28577
rect 25130 28500 25136 28552
rect 25188 28540 25194 28552
rect 25188 28512 25233 28540
rect 25188 28500 25194 28512
rect 25314 28500 25320 28552
rect 25372 28540 25378 28552
rect 25372 28512 25417 28540
rect 25372 28500 25378 28512
rect 26970 28500 26976 28552
rect 27028 28540 27034 28552
rect 27534 28543 27592 28549
rect 27534 28540 27546 28543
rect 27028 28512 27546 28540
rect 27028 28500 27034 28512
rect 27534 28509 27546 28512
rect 27580 28509 27592 28543
rect 28442 28540 28448 28552
rect 28403 28512 28448 28540
rect 27534 28503 27592 28509
rect 28442 28500 28448 28512
rect 28500 28500 28506 28552
rect 28629 28543 28687 28549
rect 28629 28509 28641 28543
rect 28675 28540 28687 28543
rect 28994 28540 29000 28552
rect 28675 28512 29000 28540
rect 28675 28509 28687 28512
rect 28629 28503 28687 28509
rect 28994 28500 29000 28512
rect 29052 28500 29058 28552
rect 29822 28540 29828 28552
rect 29783 28512 29828 28540
rect 29822 28500 29828 28512
rect 29880 28500 29886 28552
rect 30285 28543 30343 28549
rect 30285 28509 30297 28543
rect 30331 28509 30343 28543
rect 30392 28540 30420 28716
rect 30469 28713 30481 28747
rect 30515 28744 30527 28747
rect 32306 28744 32312 28756
rect 30515 28716 32312 28744
rect 30515 28713 30527 28716
rect 30469 28707 30527 28713
rect 32306 28704 32312 28716
rect 32364 28744 32370 28756
rect 32582 28744 32588 28756
rect 32364 28716 32588 28744
rect 32364 28704 32370 28716
rect 32582 28704 32588 28716
rect 32640 28704 32646 28756
rect 35802 28744 35808 28756
rect 35763 28716 35808 28744
rect 35802 28704 35808 28716
rect 35860 28704 35866 28756
rect 35526 28636 35532 28688
rect 35584 28676 35590 28688
rect 36633 28679 36691 28685
rect 36633 28676 36645 28679
rect 35584 28648 36645 28676
rect 35584 28636 35590 28648
rect 36633 28645 36645 28648
rect 36679 28676 36691 28679
rect 37185 28679 37243 28685
rect 37185 28676 37197 28679
rect 36679 28648 37197 28676
rect 36679 28645 36691 28648
rect 36633 28639 36691 28645
rect 37185 28645 37197 28648
rect 37231 28676 37243 28679
rect 37826 28676 37832 28688
rect 37231 28648 37832 28676
rect 37231 28645 37243 28648
rect 37185 28639 37243 28645
rect 37826 28636 37832 28648
rect 37884 28636 37890 28688
rect 32490 28608 32496 28620
rect 32451 28580 32496 28608
rect 32490 28568 32496 28580
rect 32548 28568 32554 28620
rect 33229 28611 33287 28617
rect 33229 28577 33241 28611
rect 33275 28608 33287 28611
rect 33410 28608 33416 28620
rect 33275 28580 33416 28608
rect 33275 28577 33287 28580
rect 33229 28571 33287 28577
rect 33410 28568 33416 28580
rect 33468 28568 33474 28620
rect 34057 28611 34115 28617
rect 34057 28577 34069 28611
rect 34103 28608 34115 28611
rect 36262 28608 36268 28620
rect 34103 28580 35112 28608
rect 34103 28577 34115 28580
rect 34057 28571 34115 28577
rect 32237 28543 32295 28549
rect 30392 28512 31892 28540
rect 30285 28503 30343 28509
rect 25406 28472 25412 28484
rect 25056 28444 25412 28472
rect 25406 28432 25412 28444
rect 25464 28432 25470 28484
rect 27798 28432 27804 28484
rect 27856 28472 27862 28484
rect 29549 28475 29607 28481
rect 29549 28472 29561 28475
rect 27856 28444 29561 28472
rect 27856 28432 27862 28444
rect 29549 28441 29561 28444
rect 29595 28441 29607 28475
rect 30300 28472 30328 28503
rect 30374 28472 30380 28484
rect 30300 28444 30380 28472
rect 29549 28435 29607 28441
rect 30374 28432 30380 28444
rect 30432 28432 30438 28484
rect 31864 28472 31892 28512
rect 32237 28509 32249 28543
rect 32283 28540 32295 28543
rect 32398 28540 32404 28552
rect 32283 28512 32404 28540
rect 32283 28509 32295 28512
rect 32237 28503 32295 28509
rect 32398 28500 32404 28512
rect 32456 28500 32462 28552
rect 32950 28540 32956 28552
rect 32911 28512 32956 28540
rect 32950 28500 32956 28512
rect 33008 28500 33014 28552
rect 33962 28540 33968 28552
rect 33923 28512 33968 28540
rect 33962 28500 33968 28512
rect 34020 28500 34026 28552
rect 34149 28543 34207 28549
rect 34149 28509 34161 28543
rect 34195 28540 34207 28543
rect 34974 28540 34980 28552
rect 34195 28512 34836 28540
rect 34935 28512 34980 28540
rect 34195 28509 34207 28512
rect 34149 28503 34207 28509
rect 34701 28475 34759 28481
rect 34701 28472 34713 28475
rect 31864 28444 34713 28472
rect 34701 28441 34713 28444
rect 34747 28441 34759 28475
rect 34701 28435 34759 28441
rect 26326 28404 26332 28416
rect 24964 28376 26332 28404
rect 24857 28367 24915 28373
rect 26326 28364 26332 28376
rect 26384 28404 26390 28416
rect 26421 28407 26479 28413
rect 26421 28404 26433 28407
rect 26384 28376 26433 28404
rect 26384 28364 26390 28376
rect 26421 28373 26433 28376
rect 26467 28373 26479 28407
rect 26421 28367 26479 28373
rect 28074 28364 28080 28416
rect 28132 28404 28138 28416
rect 29733 28407 29791 28413
rect 29733 28404 29745 28407
rect 28132 28376 29745 28404
rect 28132 28364 28138 28376
rect 29733 28373 29745 28376
rect 29779 28373 29791 28407
rect 29733 28367 29791 28373
rect 30834 28364 30840 28416
rect 30892 28404 30898 28416
rect 31113 28407 31171 28413
rect 31113 28404 31125 28407
rect 30892 28376 31125 28404
rect 30892 28364 30898 28376
rect 31113 28373 31125 28376
rect 31159 28373 31171 28407
rect 31113 28367 31171 28373
rect 31386 28364 31392 28416
rect 31444 28404 31450 28416
rect 31570 28404 31576 28416
rect 31444 28376 31576 28404
rect 31444 28364 31450 28376
rect 31570 28364 31576 28376
rect 31628 28364 31634 28416
rect 34808 28404 34836 28512
rect 34974 28500 34980 28512
rect 35032 28500 35038 28552
rect 35084 28549 35112 28580
rect 35176 28580 36268 28608
rect 35176 28549 35204 28580
rect 36262 28568 36268 28580
rect 36320 28568 36326 28620
rect 35069 28543 35127 28549
rect 35069 28509 35081 28543
rect 35115 28509 35127 28543
rect 35069 28503 35127 28509
rect 35161 28543 35219 28549
rect 35161 28509 35173 28543
rect 35207 28509 35219 28543
rect 35342 28540 35348 28552
rect 35303 28512 35348 28540
rect 35161 28503 35219 28509
rect 35342 28500 35348 28512
rect 35400 28500 35406 28552
rect 35894 28500 35900 28552
rect 35952 28540 35958 28552
rect 36173 28543 36231 28549
rect 36173 28540 36185 28543
rect 35952 28512 36185 28540
rect 35952 28500 35958 28512
rect 36173 28509 36185 28512
rect 36219 28540 36231 28543
rect 37737 28543 37795 28549
rect 37737 28540 37749 28543
rect 36219 28512 37749 28540
rect 36219 28509 36231 28512
rect 36173 28503 36231 28509
rect 37737 28509 37749 28512
rect 37783 28509 37795 28543
rect 37737 28503 37795 28509
rect 35526 28432 35532 28484
rect 35584 28472 35590 28484
rect 35989 28475 36047 28481
rect 35989 28472 36001 28475
rect 35584 28444 36001 28472
rect 35584 28432 35590 28444
rect 35989 28441 36001 28444
rect 36035 28441 36047 28475
rect 35989 28435 36047 28441
rect 35894 28404 35900 28416
rect 34808 28376 35900 28404
rect 35894 28364 35900 28376
rect 35952 28364 35958 28416
rect 1104 28314 54372 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 54372 28314
rect 1104 28240 54372 28262
rect 19705 28203 19763 28209
rect 19705 28169 19717 28203
rect 19751 28200 19763 28203
rect 19978 28200 19984 28212
rect 19751 28172 19984 28200
rect 19751 28169 19763 28172
rect 19705 28163 19763 28169
rect 19978 28160 19984 28172
rect 20036 28160 20042 28212
rect 20901 28203 20959 28209
rect 20901 28169 20913 28203
rect 20947 28200 20959 28203
rect 22002 28200 22008 28212
rect 20947 28172 22008 28200
rect 20947 28169 20959 28172
rect 20901 28163 20959 28169
rect 22002 28160 22008 28172
rect 22060 28160 22066 28212
rect 22370 28160 22376 28212
rect 22428 28200 22434 28212
rect 23201 28203 23259 28209
rect 23201 28200 23213 28203
rect 22428 28172 23213 28200
rect 22428 28160 22434 28172
rect 23201 28169 23213 28172
rect 23247 28200 23259 28203
rect 23382 28200 23388 28212
rect 23247 28172 23388 28200
rect 23247 28169 23259 28172
rect 23201 28163 23259 28169
rect 23382 28160 23388 28172
rect 23440 28160 23446 28212
rect 23934 28200 23940 28212
rect 23895 28172 23940 28200
rect 23934 28160 23940 28172
rect 23992 28160 23998 28212
rect 25314 28200 25320 28212
rect 25275 28172 25320 28200
rect 25314 28160 25320 28172
rect 25372 28160 25378 28212
rect 26326 28200 26332 28212
rect 26287 28172 26332 28200
rect 26326 28160 26332 28172
rect 26384 28160 26390 28212
rect 27798 28200 27804 28212
rect 27759 28172 27804 28200
rect 27798 28160 27804 28172
rect 27856 28160 27862 28212
rect 30469 28203 30527 28209
rect 30469 28169 30481 28203
rect 30515 28169 30527 28203
rect 30469 28163 30527 28169
rect 31573 28203 31631 28209
rect 31573 28169 31585 28203
rect 31619 28200 31631 28203
rect 31846 28200 31852 28212
rect 31619 28172 31852 28200
rect 31619 28169 31631 28172
rect 31573 28163 31631 28169
rect 19245 28135 19303 28141
rect 19245 28101 19257 28135
rect 19291 28132 19303 28135
rect 20346 28132 20352 28144
rect 19291 28104 20352 28132
rect 19291 28101 19303 28104
rect 19245 28095 19303 28101
rect 20346 28092 20352 28104
rect 20404 28132 20410 28144
rect 20533 28135 20591 28141
rect 20533 28132 20545 28135
rect 20404 28104 20545 28132
rect 20404 28092 20410 28104
rect 20533 28101 20545 28104
rect 20579 28101 20591 28135
rect 20533 28095 20591 28101
rect 20714 28092 20720 28144
rect 20772 28141 20778 28144
rect 20772 28135 20791 28141
rect 20779 28101 20791 28135
rect 20772 28095 20791 28101
rect 20772 28092 20778 28095
rect 21910 28092 21916 28144
rect 21968 28132 21974 28144
rect 22189 28135 22247 28141
rect 22189 28132 22201 28135
rect 21968 28104 22201 28132
rect 21968 28092 21974 28104
rect 22189 28101 22201 28104
rect 22235 28132 22247 28135
rect 23658 28132 23664 28144
rect 22235 28104 23664 28132
rect 22235 28101 22247 28104
rect 22189 28095 22247 28101
rect 23658 28092 23664 28104
rect 23716 28092 23722 28144
rect 24118 28132 24124 28144
rect 24079 28104 24124 28132
rect 24118 28092 24124 28104
rect 24176 28092 24182 28144
rect 25501 28135 25559 28141
rect 25501 28101 25513 28135
rect 25547 28132 25559 28135
rect 25590 28132 25596 28144
rect 25547 28104 25596 28132
rect 25547 28101 25559 28104
rect 25501 28095 25559 28101
rect 19889 28067 19947 28073
rect 19889 28033 19901 28067
rect 19935 28064 19947 28067
rect 20162 28064 20168 28076
rect 19935 28036 20168 28064
rect 19935 28033 19947 28036
rect 19889 28027 19947 28033
rect 20162 28024 20168 28036
rect 20220 28024 20226 28076
rect 22002 28064 22008 28076
rect 21963 28036 22008 28064
rect 22002 28024 22008 28036
rect 22060 28024 22066 28076
rect 22281 28067 22339 28073
rect 22281 28033 22293 28067
rect 22327 28033 22339 28067
rect 23106 28064 23112 28076
rect 23067 28036 23112 28064
rect 22281 28027 22339 28033
rect 18693 27999 18751 28005
rect 18693 27965 18705 27999
rect 18739 27996 18751 27999
rect 20073 27999 20131 28005
rect 20073 27996 20085 27999
rect 18739 27968 20085 27996
rect 18739 27965 18751 27968
rect 18693 27959 18751 27965
rect 20073 27965 20085 27968
rect 20119 27996 20131 27999
rect 20254 27996 20260 28008
rect 20119 27968 20260 27996
rect 20119 27965 20131 27968
rect 20073 27959 20131 27965
rect 20254 27956 20260 27968
rect 20312 27956 20318 28008
rect 21450 27956 21456 28008
rect 21508 27996 21514 28008
rect 22296 27996 22324 28027
rect 23106 28024 23112 28036
rect 23164 28024 23170 28076
rect 23382 28064 23388 28076
rect 23343 28036 23388 28064
rect 23382 28024 23388 28036
rect 23440 28024 23446 28076
rect 23845 28067 23903 28073
rect 23845 28033 23857 28067
rect 23891 28033 23903 28067
rect 24578 28064 24584 28076
rect 24539 28036 24584 28064
rect 23845 28027 23903 28033
rect 23860 27996 23888 28027
rect 24578 28024 24584 28036
rect 24636 28024 24642 28076
rect 24673 28067 24731 28073
rect 24673 28033 24685 28067
rect 24719 28064 24731 28067
rect 24946 28064 24952 28076
rect 24719 28036 24952 28064
rect 24719 28033 24731 28036
rect 24673 28027 24731 28033
rect 24946 28024 24952 28036
rect 25004 28024 25010 28076
rect 25516 28064 25544 28095
rect 25590 28092 25596 28104
rect 25648 28092 25654 28144
rect 26142 28092 26148 28144
rect 26200 28132 26206 28144
rect 27065 28135 27123 28141
rect 27065 28132 27077 28135
rect 26200 28104 27077 28132
rect 26200 28092 26206 28104
rect 27065 28101 27077 28104
rect 27111 28101 27123 28135
rect 28718 28132 28724 28144
rect 28679 28104 28724 28132
rect 27065 28095 27123 28101
rect 28718 28092 28724 28104
rect 28776 28092 28782 28144
rect 28810 28092 28816 28144
rect 28868 28132 28874 28144
rect 28905 28135 28963 28141
rect 28905 28132 28917 28135
rect 28868 28104 28917 28132
rect 28868 28092 28874 28104
rect 28905 28101 28917 28104
rect 28951 28101 28963 28135
rect 30484 28132 30512 28163
rect 31846 28160 31852 28172
rect 31904 28160 31910 28212
rect 35342 28160 35348 28212
rect 35400 28200 35406 28212
rect 35529 28203 35587 28209
rect 35529 28200 35541 28203
rect 35400 28172 35541 28200
rect 35400 28160 35406 28172
rect 35529 28169 35541 28172
rect 35575 28169 35587 28203
rect 35529 28163 35587 28169
rect 36265 28203 36323 28209
rect 36265 28169 36277 28203
rect 36311 28200 36323 28203
rect 36446 28200 36452 28212
rect 36311 28172 36452 28200
rect 36311 28169 36323 28172
rect 36265 28163 36323 28169
rect 36446 28160 36452 28172
rect 36504 28160 36510 28212
rect 37826 28200 37832 28212
rect 37787 28172 37832 28200
rect 37826 28160 37832 28172
rect 37884 28160 37890 28212
rect 31205 28135 31263 28141
rect 31205 28132 31217 28135
rect 30484 28104 31217 28132
rect 28905 28095 28963 28101
rect 31205 28101 31217 28104
rect 31251 28101 31263 28135
rect 31205 28095 31263 28101
rect 31294 28092 31300 28144
rect 31352 28132 31358 28144
rect 32122 28132 32128 28144
rect 31352 28104 32128 28132
rect 31352 28092 31358 28104
rect 32122 28092 32128 28104
rect 32180 28092 32186 28144
rect 33962 28092 33968 28144
rect 34020 28132 34026 28144
rect 35069 28135 35127 28141
rect 34020 28104 35020 28132
rect 34020 28092 34026 28104
rect 25240 28036 25544 28064
rect 24762 27996 24768 28008
rect 21508 27968 22324 27996
rect 23400 27968 23888 27996
rect 24136 27968 24768 27996
rect 21508 27956 21514 27968
rect 23400 27937 23428 27968
rect 24136 27937 24164 27968
rect 24762 27956 24768 27968
rect 24820 27956 24826 28008
rect 24857 27999 24915 28005
rect 24857 27965 24869 27999
rect 24903 27996 24915 27999
rect 25240 27996 25268 28036
rect 25866 28024 25872 28076
rect 25924 28064 25930 28076
rect 26973 28067 27031 28073
rect 26973 28064 26985 28067
rect 25924 28036 26985 28064
rect 25924 28024 25930 28036
rect 26973 28033 26985 28036
rect 27019 28033 27031 28067
rect 26973 28027 27031 28033
rect 27249 28067 27307 28073
rect 27249 28033 27261 28067
rect 27295 28064 27307 28067
rect 27430 28064 27436 28076
rect 27295 28036 27436 28064
rect 27295 28033 27307 28036
rect 27249 28027 27307 28033
rect 27430 28024 27436 28036
rect 27488 28024 27494 28076
rect 28074 28064 28080 28076
rect 28035 28036 28080 28064
rect 28074 28024 28080 28036
rect 28132 28024 28138 28076
rect 29822 28064 29828 28076
rect 29012 28036 29828 28064
rect 24903 27968 25268 27996
rect 27801 27999 27859 28005
rect 24903 27965 24915 27968
rect 24857 27959 24915 27965
rect 27801 27965 27813 27999
rect 27847 27996 27859 27999
rect 27890 27996 27896 28008
rect 27847 27968 27896 27996
rect 27847 27965 27859 27968
rect 27801 27959 27859 27965
rect 23385 27931 23443 27937
rect 23385 27897 23397 27931
rect 23431 27897 23443 27931
rect 23385 27891 23443 27897
rect 24121 27931 24179 27937
rect 24121 27897 24133 27931
rect 24167 27897 24179 27931
rect 24872 27928 24900 27959
rect 27890 27956 27896 27968
rect 27948 27956 27954 28008
rect 27985 27999 28043 28005
rect 27985 27965 27997 27999
rect 28031 27996 28043 27999
rect 29012 27996 29040 28036
rect 29822 28024 29828 28036
rect 29880 28024 29886 28076
rect 30101 28067 30159 28073
rect 30101 28033 30113 28067
rect 30147 28064 30159 28067
rect 30834 28064 30840 28076
rect 30147 28036 30840 28064
rect 30147 28033 30159 28036
rect 30101 28027 30159 28033
rect 30834 28024 30840 28036
rect 30892 28024 30898 28076
rect 30926 28024 30932 28076
rect 30984 28064 30990 28076
rect 31077 28067 31135 28073
rect 30984 28036 31029 28064
rect 30984 28024 30990 28036
rect 31077 28033 31089 28067
rect 31123 28064 31135 28067
rect 31435 28067 31493 28073
rect 31123 28036 31248 28064
rect 31123 28033 31135 28036
rect 31077 28027 31135 28033
rect 28031 27968 29040 27996
rect 28031 27965 28043 27968
rect 27985 27959 28043 27965
rect 29086 27956 29092 28008
rect 29144 27996 29150 28008
rect 30009 27999 30067 28005
rect 30009 27996 30021 27999
rect 29144 27968 30021 27996
rect 29144 27956 29150 27968
rect 30009 27965 30021 27968
rect 30055 27965 30067 27999
rect 31220 27996 31248 28036
rect 31435 28033 31447 28067
rect 31481 28064 31493 28067
rect 31570 28064 31576 28076
rect 31481 28036 31576 28064
rect 31481 28033 31493 28036
rect 31435 28027 31493 28033
rect 31570 28024 31576 28036
rect 31628 28024 31634 28076
rect 32306 28064 32312 28076
rect 32267 28036 32312 28064
rect 32306 28024 32312 28036
rect 32364 28024 32370 28076
rect 32674 28024 32680 28076
rect 32732 28064 32738 28076
rect 32769 28067 32827 28073
rect 32769 28064 32781 28067
rect 32732 28036 32781 28064
rect 32732 28024 32738 28036
rect 32769 28033 32781 28036
rect 32815 28033 32827 28067
rect 32769 28027 32827 28033
rect 32953 28067 33011 28073
rect 32953 28033 32965 28067
rect 32999 28033 33011 28067
rect 32953 28027 33011 28033
rect 32030 27996 32036 28008
rect 31220 27968 32036 27996
rect 30009 27959 30067 27965
rect 32030 27956 32036 27968
rect 32088 27956 32094 28008
rect 24121 27891 24179 27897
rect 24688 27900 24900 27928
rect 20717 27863 20775 27869
rect 20717 27829 20729 27863
rect 20763 27860 20775 27863
rect 20806 27860 20812 27872
rect 20763 27832 20812 27860
rect 20763 27829 20775 27832
rect 20717 27823 20775 27829
rect 20806 27820 20812 27832
rect 20864 27820 20870 27872
rect 21266 27820 21272 27872
rect 21324 27860 21330 27872
rect 21821 27863 21879 27869
rect 21821 27860 21833 27863
rect 21324 27832 21833 27860
rect 21324 27820 21330 27832
rect 21821 27829 21833 27832
rect 21867 27829 21879 27863
rect 21821 27823 21879 27829
rect 23198 27820 23204 27872
rect 23256 27860 23262 27872
rect 24688 27860 24716 27900
rect 24946 27888 24952 27940
rect 25004 27928 25010 27940
rect 25869 27931 25927 27937
rect 25869 27928 25881 27931
rect 25004 27900 25881 27928
rect 25004 27888 25010 27900
rect 25869 27897 25881 27900
rect 25915 27928 25927 27931
rect 26050 27928 26056 27940
rect 25915 27900 26056 27928
rect 25915 27897 25927 27900
rect 25869 27891 25927 27897
rect 26050 27888 26056 27900
rect 26108 27888 26114 27940
rect 27246 27928 27252 27940
rect 27207 27900 27252 27928
rect 27246 27888 27252 27900
rect 27304 27888 27310 27940
rect 28442 27888 28448 27940
rect 28500 27928 28506 27940
rect 28500 27900 29500 27928
rect 28500 27888 28506 27900
rect 23256 27832 24716 27860
rect 24765 27863 24823 27869
rect 23256 27820 23262 27832
rect 24765 27829 24777 27863
rect 24811 27860 24823 27863
rect 25314 27860 25320 27872
rect 24811 27832 25320 27860
rect 24811 27829 24823 27832
rect 24765 27823 24823 27829
rect 25314 27820 25320 27832
rect 25372 27820 25378 27872
rect 25498 27860 25504 27872
rect 25459 27832 25504 27860
rect 25498 27820 25504 27832
rect 25556 27820 25562 27872
rect 28537 27863 28595 27869
rect 28537 27829 28549 27863
rect 28583 27860 28595 27863
rect 28718 27860 28724 27872
rect 28583 27832 28724 27860
rect 28583 27829 28595 27832
rect 28537 27823 28595 27829
rect 28718 27820 28724 27832
rect 28776 27820 28782 27872
rect 29472 27869 29500 27900
rect 30374 27888 30380 27940
rect 30432 27928 30438 27940
rect 30926 27928 30932 27940
rect 30432 27900 30932 27928
rect 30432 27888 30438 27900
rect 30926 27888 30932 27900
rect 30984 27888 30990 27940
rect 31018 27888 31024 27940
rect 31076 27928 31082 27940
rect 31662 27928 31668 27940
rect 31076 27900 31668 27928
rect 31076 27888 31082 27900
rect 31662 27888 31668 27900
rect 31720 27928 31726 27940
rect 32968 27928 32996 28027
rect 34422 28024 34428 28076
rect 34480 28024 34486 28076
rect 34992 28064 35020 28104
rect 35069 28101 35081 28135
rect 35115 28132 35127 28135
rect 35618 28132 35624 28144
rect 35115 28104 35624 28132
rect 35115 28101 35127 28104
rect 35069 28095 35127 28101
rect 35618 28092 35624 28104
rect 35676 28092 35682 28144
rect 36004 28104 36400 28132
rect 35526 28064 35532 28076
rect 34992 28036 35532 28064
rect 35526 28024 35532 28036
rect 35584 28024 35590 28076
rect 35713 28067 35771 28073
rect 35713 28033 35725 28067
rect 35759 28064 35771 28067
rect 35894 28064 35900 28076
rect 35759 28036 35900 28064
rect 35759 28033 35771 28036
rect 35713 28027 35771 28033
rect 35894 28024 35900 28036
rect 35952 28024 35958 28076
rect 34238 27996 34244 28008
rect 34199 27968 34244 27996
rect 34238 27956 34244 27968
rect 34296 27956 34302 28008
rect 34440 27996 34468 28024
rect 36004 27996 36032 28104
rect 36372 28073 36400 28104
rect 36173 28067 36231 28073
rect 36173 28033 36185 28067
rect 36219 28033 36231 28067
rect 36173 28027 36231 28033
rect 36357 28067 36415 28073
rect 36357 28033 36369 28067
rect 36403 28064 36415 28067
rect 36446 28064 36452 28076
rect 36403 28036 36452 28064
rect 36403 28033 36415 28036
rect 36357 28027 36415 28033
rect 34440 27968 36032 27996
rect 34054 27928 34060 27940
rect 31720 27900 32996 27928
rect 33152 27900 34060 27928
rect 31720 27888 31726 27900
rect 29457 27863 29515 27869
rect 29457 27829 29469 27863
rect 29503 27860 29515 27863
rect 33152 27860 33180 27900
rect 34054 27888 34060 27900
rect 34112 27888 34118 27940
rect 34256 27928 34284 27956
rect 36188 27928 36216 28027
rect 36446 28024 36452 28036
rect 36504 28024 36510 28076
rect 53374 27996 53380 28008
rect 53335 27968 53380 27996
rect 53374 27956 53380 27968
rect 53432 27956 53438 28008
rect 53650 27996 53656 28008
rect 53611 27968 53656 27996
rect 53650 27956 53656 27968
rect 53708 27956 53714 28008
rect 37277 27931 37335 27937
rect 37277 27928 37289 27931
rect 34256 27900 37289 27928
rect 37277 27897 37289 27900
rect 37323 27928 37335 27931
rect 37550 27928 37556 27940
rect 37323 27900 37556 27928
rect 37323 27897 37335 27900
rect 37277 27891 37335 27897
rect 37550 27888 37556 27900
rect 37608 27888 37614 27940
rect 29503 27832 33180 27860
rect 29503 27829 29515 27832
rect 29457 27823 29515 27829
rect 1104 27770 54372 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 54372 27770
rect 1104 27696 54372 27718
rect 18874 27616 18880 27668
rect 18932 27656 18938 27668
rect 19521 27659 19579 27665
rect 19521 27656 19533 27659
rect 18932 27628 19533 27656
rect 18932 27616 18938 27628
rect 19521 27625 19533 27628
rect 19567 27625 19579 27659
rect 19521 27619 19579 27625
rect 21358 27616 21364 27668
rect 21416 27656 21422 27668
rect 21637 27659 21695 27665
rect 21637 27656 21649 27659
rect 21416 27628 21649 27656
rect 21416 27616 21422 27628
rect 21637 27625 21649 27628
rect 21683 27656 21695 27659
rect 22370 27656 22376 27668
rect 21683 27628 22376 27656
rect 21683 27625 21695 27628
rect 21637 27619 21695 27625
rect 22370 27616 22376 27628
rect 22428 27616 22434 27668
rect 23382 27616 23388 27668
rect 23440 27656 23446 27668
rect 25682 27656 25688 27668
rect 23440 27628 25688 27656
rect 23440 27616 23446 27628
rect 25682 27616 25688 27628
rect 25740 27616 25746 27668
rect 27890 27656 27896 27668
rect 27851 27628 27896 27656
rect 27890 27616 27896 27628
rect 27948 27616 27954 27668
rect 31294 27656 31300 27668
rect 31255 27628 31300 27656
rect 31294 27616 31300 27628
rect 31352 27616 31358 27668
rect 36446 27656 36452 27668
rect 31404 27628 32628 27656
rect 36407 27628 36452 27656
rect 19889 27591 19947 27597
rect 19889 27557 19901 27591
rect 19935 27588 19947 27591
rect 20714 27588 20720 27600
rect 19935 27560 20720 27588
rect 19935 27557 19947 27560
rect 19889 27551 19947 27557
rect 20714 27548 20720 27560
rect 20772 27548 20778 27600
rect 22925 27591 22983 27597
rect 22925 27557 22937 27591
rect 22971 27588 22983 27591
rect 25593 27591 25651 27597
rect 25593 27588 25605 27591
rect 22971 27560 25605 27588
rect 22971 27557 22983 27560
rect 22925 27551 22983 27557
rect 25593 27557 25605 27560
rect 25639 27557 25651 27591
rect 25866 27588 25872 27600
rect 25827 27560 25872 27588
rect 25593 27551 25651 27557
rect 25866 27548 25872 27560
rect 25924 27548 25930 27600
rect 26329 27591 26387 27597
rect 26329 27557 26341 27591
rect 26375 27588 26387 27591
rect 28810 27588 28816 27600
rect 26375 27560 28816 27588
rect 26375 27557 26387 27560
rect 26329 27551 26387 27557
rect 21450 27520 21456 27532
rect 21411 27492 21456 27520
rect 21450 27480 21456 27492
rect 21508 27480 21514 27532
rect 23658 27480 23664 27532
rect 23716 27520 23722 27532
rect 23753 27523 23811 27529
rect 23753 27520 23765 27523
rect 23716 27492 23765 27520
rect 23716 27480 23722 27492
rect 23753 27489 23765 27492
rect 23799 27489 23811 27523
rect 23753 27483 23811 27489
rect 24673 27523 24731 27529
rect 24673 27489 24685 27523
rect 24719 27520 24731 27523
rect 25501 27523 25559 27529
rect 25501 27520 25513 27523
rect 24719 27492 25513 27520
rect 24719 27489 24731 27492
rect 24673 27483 24731 27489
rect 25501 27489 25513 27492
rect 25547 27489 25559 27523
rect 26344 27520 26372 27551
rect 28810 27548 28816 27560
rect 28868 27548 28874 27600
rect 28994 27588 29000 27600
rect 28955 27560 29000 27588
rect 28994 27548 29000 27560
rect 29052 27548 29058 27600
rect 29638 27588 29644 27600
rect 29599 27560 29644 27588
rect 29638 27548 29644 27560
rect 29696 27548 29702 27600
rect 30926 27548 30932 27600
rect 30984 27588 30990 27600
rect 31404 27588 31432 27628
rect 30984 27560 31432 27588
rect 30984 27548 30990 27560
rect 31478 27548 31484 27600
rect 31536 27588 31542 27600
rect 31536 27560 31581 27588
rect 31536 27548 31542 27560
rect 25501 27483 25559 27489
rect 25608 27492 26372 27520
rect 1673 27455 1731 27461
rect 1673 27421 1685 27455
rect 1719 27421 1731 27455
rect 1673 27415 1731 27421
rect 1688 27384 1716 27415
rect 19426 27412 19432 27464
rect 19484 27452 19490 27464
rect 19521 27455 19579 27461
rect 19521 27452 19533 27455
rect 19484 27424 19533 27452
rect 19484 27412 19490 27424
rect 19521 27421 19533 27424
rect 19567 27421 19579 27455
rect 19521 27415 19579 27421
rect 19705 27455 19763 27461
rect 19705 27421 19717 27455
rect 19751 27452 19763 27455
rect 20070 27452 20076 27464
rect 19751 27424 20076 27452
rect 19751 27421 19763 27424
rect 19705 27415 19763 27421
rect 20070 27412 20076 27424
rect 20128 27412 20134 27464
rect 20717 27455 20775 27461
rect 20717 27421 20729 27455
rect 20763 27452 20775 27455
rect 21082 27452 21088 27464
rect 20763 27424 21088 27452
rect 20763 27421 20775 27424
rect 20717 27415 20775 27421
rect 21082 27412 21088 27424
rect 21140 27452 21146 27464
rect 21361 27455 21419 27461
rect 21361 27452 21373 27455
rect 21140 27424 21373 27452
rect 21140 27412 21146 27424
rect 21361 27421 21373 27424
rect 21407 27452 21419 27455
rect 21910 27452 21916 27464
rect 21407 27424 21916 27452
rect 21407 27421 21419 27424
rect 21361 27415 21419 27421
rect 21910 27412 21916 27424
rect 21968 27412 21974 27464
rect 22554 27412 22560 27464
rect 22612 27452 22618 27464
rect 22741 27455 22799 27461
rect 22741 27452 22753 27455
rect 22612 27424 22753 27452
rect 22612 27412 22618 27424
rect 22741 27421 22753 27424
rect 22787 27421 22799 27455
rect 22741 27415 22799 27421
rect 24118 27412 24124 27464
rect 24176 27452 24182 27464
rect 24581 27455 24639 27461
rect 24581 27452 24593 27455
rect 24176 27424 24593 27452
rect 24176 27412 24182 27424
rect 24581 27421 24593 27424
rect 24627 27421 24639 27455
rect 24581 27415 24639 27421
rect 25225 27455 25283 27461
rect 25225 27421 25237 27455
rect 25271 27421 25283 27455
rect 25225 27415 25283 27421
rect 2225 27387 2283 27393
rect 2225 27384 2237 27387
rect 1688 27356 2237 27384
rect 2225 27353 2237 27356
rect 2271 27384 2283 27387
rect 16574 27384 16580 27396
rect 2271 27356 16580 27384
rect 2271 27353 2283 27356
rect 2225 27347 2283 27353
rect 16574 27344 16580 27356
rect 16632 27344 16638 27396
rect 22186 27344 22192 27396
rect 22244 27384 22250 27396
rect 22373 27387 22431 27393
rect 22373 27384 22385 27387
rect 22244 27356 22385 27384
rect 22244 27344 22250 27356
rect 22373 27353 22385 27356
rect 22419 27353 22431 27387
rect 22646 27384 22652 27396
rect 22607 27356 22652 27384
rect 22373 27347 22431 27353
rect 22646 27344 22652 27356
rect 22704 27344 22710 27396
rect 1486 27316 1492 27328
rect 1447 27288 1492 27316
rect 1486 27276 1492 27288
rect 1544 27276 1550 27328
rect 22278 27276 22284 27328
rect 22336 27316 22342 27328
rect 22557 27319 22615 27325
rect 22557 27316 22569 27319
rect 22336 27288 22569 27316
rect 22336 27276 22342 27288
rect 22557 27285 22569 27288
rect 22603 27285 22615 27319
rect 24596 27316 24624 27415
rect 25240 27384 25268 27415
rect 25314 27412 25320 27464
rect 25372 27452 25378 27464
rect 25409 27455 25467 27461
rect 25409 27452 25421 27455
rect 25372 27424 25421 27452
rect 25372 27412 25378 27424
rect 25409 27421 25421 27424
rect 25455 27421 25467 27455
rect 25409 27415 25467 27421
rect 25608 27384 25636 27492
rect 27614 27480 27620 27532
rect 27672 27480 27678 27532
rect 29546 27480 29552 27532
rect 29604 27520 29610 27532
rect 30193 27523 30251 27529
rect 30193 27520 30205 27523
rect 29604 27492 30205 27520
rect 29604 27480 29610 27492
rect 30193 27489 30205 27492
rect 30239 27489 30251 27523
rect 30193 27483 30251 27489
rect 30653 27523 30711 27529
rect 30653 27489 30665 27523
rect 30699 27520 30711 27523
rect 31570 27520 31576 27532
rect 30699 27492 31576 27520
rect 30699 27489 30711 27492
rect 30653 27483 30711 27489
rect 31570 27480 31576 27492
rect 31628 27480 31634 27532
rect 31938 27520 31944 27532
rect 31899 27492 31944 27520
rect 31938 27480 31944 27492
rect 31996 27480 32002 27532
rect 25682 27412 25688 27464
rect 25740 27452 25746 27464
rect 25740 27424 25785 27452
rect 25740 27412 25746 27424
rect 26050 27412 26056 27464
rect 26108 27452 26114 27464
rect 26513 27455 26571 27461
rect 26513 27452 26525 27455
rect 26108 27424 26525 27452
rect 26108 27412 26114 27424
rect 26513 27421 26525 27424
rect 26559 27421 26571 27455
rect 26513 27415 26571 27421
rect 26602 27412 26608 27464
rect 26660 27452 26666 27464
rect 27632 27452 27660 27480
rect 26660 27424 27660 27452
rect 26660 27412 26666 27424
rect 28166 27412 28172 27464
rect 28224 27452 28230 27464
rect 28353 27455 28411 27461
rect 28353 27452 28365 27455
rect 28224 27424 28365 27452
rect 28224 27412 28230 27424
rect 28353 27421 28365 27424
rect 28399 27421 28411 27455
rect 28718 27452 28724 27464
rect 28679 27424 28724 27452
rect 28353 27415 28411 27421
rect 28718 27412 28724 27424
rect 28776 27412 28782 27464
rect 28813 27455 28871 27461
rect 28813 27421 28825 27455
rect 28859 27452 28871 27455
rect 29086 27452 29092 27464
rect 28859 27424 29092 27452
rect 28859 27421 28871 27424
rect 28813 27415 28871 27421
rect 29086 27412 29092 27424
rect 29144 27412 29150 27464
rect 30006 27412 30012 27464
rect 30064 27452 30070 27464
rect 30285 27455 30343 27461
rect 30285 27452 30297 27455
rect 30064 27424 30297 27452
rect 30064 27412 30070 27424
rect 30285 27421 30297 27424
rect 30331 27452 30343 27455
rect 32122 27452 32128 27464
rect 30331 27424 31356 27452
rect 32083 27424 32128 27452
rect 30331 27421 30343 27424
rect 30285 27415 30343 27421
rect 25240 27356 25636 27384
rect 25884 27356 27568 27384
rect 25884 27316 25912 27356
rect 24596 27288 25912 27316
rect 22557 27279 22615 27285
rect 25958 27276 25964 27328
rect 26016 27316 26022 27328
rect 27157 27319 27215 27325
rect 27157 27316 27169 27319
rect 26016 27288 27169 27316
rect 26016 27276 26022 27288
rect 27157 27285 27169 27288
rect 27203 27285 27215 27319
rect 27540 27316 27568 27356
rect 27614 27344 27620 27396
rect 27672 27384 27678 27396
rect 28491 27387 28549 27393
rect 28491 27384 28503 27387
rect 27672 27356 28503 27384
rect 27672 27344 27678 27356
rect 28491 27353 28503 27356
rect 28537 27353 28549 27387
rect 28491 27347 28549 27353
rect 28626 27344 28632 27396
rect 28684 27384 28690 27396
rect 28684 27356 28729 27384
rect 28684 27344 28690 27356
rect 31018 27344 31024 27396
rect 31076 27384 31082 27396
rect 31113 27387 31171 27393
rect 31113 27384 31125 27387
rect 31076 27356 31125 27384
rect 31076 27344 31082 27356
rect 31113 27353 31125 27356
rect 31159 27353 31171 27387
rect 31328 27384 31356 27424
rect 32122 27412 32128 27424
rect 32180 27412 32186 27464
rect 32398 27412 32404 27464
rect 32456 27452 32462 27464
rect 32600 27452 32628 27628
rect 36446 27616 36452 27628
rect 36504 27656 36510 27668
rect 37001 27659 37059 27665
rect 37001 27656 37013 27659
rect 36504 27628 37013 27656
rect 36504 27616 36510 27628
rect 37001 27625 37013 27628
rect 37047 27625 37059 27659
rect 37550 27656 37556 27668
rect 37511 27628 37556 27656
rect 37001 27619 37059 27625
rect 37550 27616 37556 27628
rect 37608 27616 37614 27668
rect 53650 27656 53656 27668
rect 53611 27628 53656 27656
rect 53650 27616 53656 27628
rect 53708 27616 53714 27668
rect 34146 27480 34152 27532
rect 34204 27520 34210 27532
rect 34793 27523 34851 27529
rect 34793 27520 34805 27523
rect 34204 27492 34805 27520
rect 34204 27480 34210 27492
rect 34793 27489 34805 27492
rect 34839 27489 34851 27523
rect 34793 27483 34851 27489
rect 32677 27455 32735 27461
rect 32677 27452 32689 27455
rect 32456 27424 32689 27452
rect 32456 27412 32462 27424
rect 32677 27421 32689 27424
rect 32723 27452 32735 27455
rect 33778 27452 33784 27464
rect 32723 27424 33784 27452
rect 32723 27421 32735 27424
rect 32677 27415 32735 27421
rect 33778 27412 33784 27424
rect 33836 27412 33842 27464
rect 35342 27452 35348 27464
rect 35303 27424 35348 27452
rect 35342 27412 35348 27424
rect 35400 27412 35406 27464
rect 31478 27384 31484 27396
rect 31328 27356 31484 27384
rect 31113 27347 31171 27353
rect 31478 27344 31484 27356
rect 31536 27344 31542 27396
rect 27798 27316 27804 27328
rect 27540 27288 27804 27316
rect 27157 27279 27215 27285
rect 27798 27276 27804 27288
rect 27856 27276 27862 27328
rect 30374 27276 30380 27328
rect 30432 27316 30438 27328
rect 31313 27319 31371 27325
rect 31313 27316 31325 27319
rect 30432 27288 31325 27316
rect 30432 27276 30438 27288
rect 31313 27285 31325 27288
rect 31359 27285 31371 27319
rect 35894 27316 35900 27328
rect 35855 27288 35900 27316
rect 31313 27279 31371 27285
rect 35894 27276 35900 27288
rect 35952 27276 35958 27328
rect 37550 27276 37556 27328
rect 37608 27316 37614 27328
rect 41506 27316 41512 27328
rect 37608 27288 41512 27316
rect 37608 27276 37614 27288
rect 41506 27276 41512 27288
rect 41564 27276 41570 27328
rect 1104 27226 54372 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 54372 27226
rect 1104 27152 54372 27174
rect 20162 27072 20168 27124
rect 20220 27112 20226 27124
rect 20349 27115 20407 27121
rect 20349 27112 20361 27115
rect 20220 27084 20361 27112
rect 20220 27072 20226 27084
rect 20349 27081 20361 27084
rect 20395 27081 20407 27115
rect 20349 27075 20407 27081
rect 22649 27115 22707 27121
rect 22649 27081 22661 27115
rect 22695 27112 22707 27115
rect 24118 27112 24124 27124
rect 22695 27084 24124 27112
rect 22695 27081 22707 27084
rect 22649 27075 22707 27081
rect 24118 27072 24124 27084
rect 24176 27072 24182 27124
rect 24305 27115 24363 27121
rect 24305 27081 24317 27115
rect 24351 27112 24363 27115
rect 25130 27112 25136 27124
rect 24351 27084 25136 27112
rect 24351 27081 24363 27084
rect 24305 27075 24363 27081
rect 25130 27072 25136 27084
rect 25188 27072 25194 27124
rect 25406 27072 25412 27124
rect 25464 27112 25470 27124
rect 25501 27115 25559 27121
rect 25501 27112 25513 27115
rect 25464 27084 25513 27112
rect 25464 27072 25470 27084
rect 25501 27081 25513 27084
rect 25547 27081 25559 27115
rect 26142 27112 26148 27124
rect 26103 27084 26148 27112
rect 25501 27075 25559 27081
rect 26142 27072 26148 27084
rect 26200 27072 26206 27124
rect 28626 27112 28632 27124
rect 27549 27084 28632 27112
rect 19889 27047 19947 27053
rect 19889 27013 19901 27047
rect 19935 27044 19947 27047
rect 20254 27044 20260 27056
rect 19935 27016 20260 27044
rect 19935 27013 19947 27016
rect 19889 27007 19947 27013
rect 20254 27004 20260 27016
rect 20312 27004 20318 27056
rect 21269 27047 21327 27053
rect 21269 27013 21281 27047
rect 21315 27044 21327 27047
rect 23198 27044 23204 27056
rect 21315 27016 22324 27044
rect 23159 27016 23204 27044
rect 21315 27013 21327 27016
rect 21269 27007 21327 27013
rect 22296 26988 22324 27016
rect 23198 27004 23204 27016
rect 23256 27004 23262 27056
rect 25317 27047 25375 27053
rect 25317 27044 25329 27047
rect 24228 27016 25329 27044
rect 24228 26988 24256 27016
rect 25317 27013 25329 27016
rect 25363 27013 25375 27047
rect 25317 27007 25375 27013
rect 25590 27004 25596 27056
rect 25648 27044 25654 27056
rect 27549 27044 27577 27084
rect 28626 27072 28632 27084
rect 28684 27072 28690 27124
rect 29546 27112 29552 27124
rect 29507 27084 29552 27112
rect 29546 27072 29552 27084
rect 29604 27072 29610 27124
rect 30374 27112 30380 27124
rect 30335 27084 30380 27112
rect 30374 27072 30380 27084
rect 30432 27072 30438 27124
rect 30834 27072 30840 27124
rect 30892 27112 30898 27124
rect 31481 27115 31539 27121
rect 31481 27112 31493 27115
rect 30892 27084 31493 27112
rect 30892 27072 30898 27084
rect 25648 27016 27577 27044
rect 25648 27004 25654 27016
rect 27614 27004 27620 27056
rect 27672 27044 27678 27056
rect 27672 27016 29408 27044
rect 27672 27004 27678 27016
rect 20990 26976 20996 26988
rect 20951 26948 20996 26976
rect 20990 26936 20996 26948
rect 21048 26936 21054 26988
rect 21085 26979 21143 26985
rect 21085 26945 21097 26979
rect 21131 26976 21143 26979
rect 21450 26976 21456 26988
rect 21131 26948 21456 26976
rect 21131 26945 21143 26948
rect 21085 26939 21143 26945
rect 21450 26936 21456 26948
rect 21508 26936 21514 26988
rect 22186 26976 22192 26988
rect 22147 26948 22192 26976
rect 22186 26936 22192 26948
rect 22244 26936 22250 26988
rect 22278 26936 22284 26988
rect 22336 26976 22342 26988
rect 22465 26979 22523 26985
rect 22336 26948 22381 26976
rect 22336 26936 22342 26948
rect 22465 26945 22477 26979
rect 22511 26976 22523 26979
rect 22554 26976 22560 26988
rect 22511 26948 22560 26976
rect 22511 26945 22523 26948
rect 22465 26939 22523 26945
rect 22554 26936 22560 26948
rect 22612 26936 22618 26988
rect 24210 26976 24216 26988
rect 24171 26948 24216 26976
rect 24210 26936 24216 26948
rect 24268 26936 24274 26988
rect 24397 26979 24455 26985
rect 24397 26945 24409 26979
rect 24443 26976 24455 26979
rect 24486 26976 24492 26988
rect 24443 26948 24492 26976
rect 24443 26945 24455 26948
rect 24397 26939 24455 26945
rect 24486 26936 24492 26948
rect 24544 26976 24550 26988
rect 25133 26979 25191 26985
rect 25133 26976 25145 26979
rect 24544 26948 25145 26976
rect 24544 26936 24550 26948
rect 25133 26945 25145 26948
rect 25179 26945 25191 26979
rect 26234 26976 26240 26988
rect 26195 26948 26240 26976
rect 25133 26939 25191 26945
rect 26234 26936 26240 26948
rect 26292 26936 26298 26988
rect 26421 26979 26479 26985
rect 26421 26945 26433 26979
rect 26467 26945 26479 26979
rect 26421 26939 26479 26945
rect 21266 26908 21272 26920
rect 21227 26880 21272 26908
rect 21266 26868 21272 26880
rect 21324 26868 21330 26920
rect 22373 26911 22431 26917
rect 22373 26877 22385 26911
rect 22419 26908 22431 26911
rect 22646 26908 22652 26920
rect 22419 26880 22652 26908
rect 22419 26877 22431 26880
rect 22373 26871 22431 26877
rect 22646 26868 22652 26880
rect 22704 26868 22710 26920
rect 23753 26911 23811 26917
rect 23753 26877 23765 26911
rect 23799 26908 23811 26911
rect 25222 26908 25228 26920
rect 23799 26880 25228 26908
rect 23799 26877 23811 26880
rect 23753 26871 23811 26877
rect 25222 26868 25228 26880
rect 25280 26868 25286 26920
rect 26142 26868 26148 26920
rect 26200 26908 26206 26920
rect 26436 26908 26464 26939
rect 27338 26936 27344 26988
rect 27396 26976 27402 26988
rect 27433 26979 27491 26985
rect 27433 26976 27445 26979
rect 27396 26948 27445 26976
rect 27396 26936 27402 26948
rect 27433 26945 27445 26948
rect 27479 26945 27491 26979
rect 27890 26976 27896 26988
rect 27851 26948 27896 26976
rect 27433 26939 27491 26945
rect 27890 26936 27896 26948
rect 27948 26936 27954 26988
rect 27982 26936 27988 26988
rect 28040 26976 28046 26988
rect 28169 26979 28227 26985
rect 28040 26948 28085 26976
rect 28040 26936 28046 26948
rect 28169 26945 28181 26979
rect 28215 26976 28227 26979
rect 28258 26976 28264 26988
rect 28215 26948 28264 26976
rect 28215 26945 28227 26948
rect 28169 26939 28227 26945
rect 26973 26911 27031 26917
rect 26973 26908 26985 26911
rect 26200 26880 26985 26908
rect 26200 26868 26206 26880
rect 26973 26877 26985 26880
rect 27019 26877 27031 26911
rect 28184 26908 28212 26939
rect 28258 26936 28264 26948
rect 28316 26936 28322 26988
rect 29380 26985 29408 27016
rect 30116 27016 31064 27044
rect 30116 26988 30144 27016
rect 29365 26979 29423 26985
rect 29365 26945 29377 26979
rect 29411 26945 29423 26979
rect 30098 26976 30104 26988
rect 30059 26948 30104 26976
rect 29365 26939 29423 26945
rect 30098 26936 30104 26948
rect 30156 26936 30162 26988
rect 31036 26985 31064 27016
rect 30837 26979 30895 26985
rect 30837 26976 30849 26979
rect 30208 26948 30849 26976
rect 29178 26908 29184 26920
rect 26973 26871 27031 26877
rect 27080 26880 28212 26908
rect 29139 26880 29184 26908
rect 26418 26800 26424 26852
rect 26476 26840 26482 26852
rect 27080 26840 27108 26880
rect 29178 26868 29184 26880
rect 29236 26868 29242 26920
rect 29270 26868 29276 26920
rect 29328 26908 29334 26920
rect 30208 26908 30236 26948
rect 30837 26945 30849 26948
rect 30883 26945 30895 26979
rect 30837 26939 30895 26945
rect 31021 26979 31079 26985
rect 31021 26945 31033 26979
rect 31067 26945 31079 26979
rect 31021 26939 31079 26945
rect 30374 26908 30380 26920
rect 29328 26880 30236 26908
rect 30335 26880 30380 26908
rect 29328 26868 29334 26880
rect 30374 26868 30380 26880
rect 30432 26868 30438 26920
rect 31312 26908 31340 27084
rect 31481 27081 31493 27084
rect 31527 27081 31539 27115
rect 31481 27075 31539 27081
rect 32585 27115 32643 27121
rect 32585 27081 32597 27115
rect 32631 27112 32643 27115
rect 32950 27112 32956 27124
rect 32631 27084 32956 27112
rect 32631 27081 32643 27084
rect 32585 27075 32643 27081
rect 32950 27072 32956 27084
rect 33008 27072 33014 27124
rect 32122 27004 32128 27056
rect 32180 27044 32186 27056
rect 32217 27047 32275 27053
rect 32217 27044 32229 27047
rect 32180 27016 32229 27044
rect 32180 27004 32186 27016
rect 32217 27013 32229 27016
rect 32263 27013 32275 27047
rect 32398 27044 32404 27056
rect 32359 27016 32404 27044
rect 32217 27007 32275 27013
rect 32398 27004 32404 27016
rect 32456 27004 32462 27056
rect 33778 27004 33784 27056
rect 33836 27044 33842 27056
rect 34885 27047 34943 27053
rect 34885 27044 34897 27047
rect 33836 27016 34897 27044
rect 33836 27004 33842 27016
rect 34885 27013 34897 27016
rect 34931 27013 34943 27047
rect 34885 27007 34943 27013
rect 31478 26936 31484 26988
rect 31536 26976 31542 26988
rect 33137 26979 33195 26985
rect 33137 26976 33149 26979
rect 31536 26948 33149 26976
rect 31536 26936 31542 26948
rect 33137 26945 33149 26948
rect 33183 26945 33195 26979
rect 33137 26939 33195 26945
rect 33965 26979 34023 26985
rect 33965 26945 33977 26979
rect 34011 26976 34023 26979
rect 34330 26976 34336 26988
rect 34011 26948 34336 26976
rect 34011 26945 34023 26948
rect 33965 26939 34023 26945
rect 34330 26936 34336 26948
rect 34388 26976 34394 26988
rect 34606 26976 34612 26988
rect 34388 26948 34612 26976
rect 34388 26936 34394 26948
rect 34606 26936 34612 26948
rect 34664 26936 34670 26988
rect 35713 26979 35771 26985
rect 35713 26945 35725 26979
rect 35759 26976 35771 26979
rect 36078 26976 36084 26988
rect 35759 26948 36084 26976
rect 35759 26945 35771 26948
rect 35713 26939 35771 26945
rect 36078 26936 36084 26948
rect 36136 26936 36142 26988
rect 34054 26908 34060 26920
rect 31312 26880 34060 26908
rect 34054 26868 34060 26880
rect 34112 26868 34118 26920
rect 28166 26840 28172 26852
rect 26476 26812 27108 26840
rect 28127 26812 28172 26840
rect 26476 26800 26482 26812
rect 28166 26800 28172 26812
rect 28224 26800 28230 26852
rect 29822 26800 29828 26852
rect 29880 26840 29886 26852
rect 30837 26843 30895 26849
rect 30837 26840 30849 26843
rect 29880 26812 30849 26840
rect 29880 26800 29886 26812
rect 30837 26809 30849 26812
rect 30883 26809 30895 26843
rect 30837 26803 30895 26809
rect 25958 26772 25964 26784
rect 25919 26744 25964 26772
rect 25958 26732 25964 26744
rect 26016 26732 26022 26784
rect 27154 26772 27160 26784
rect 27115 26744 27160 26772
rect 27154 26732 27160 26744
rect 27212 26732 27218 26784
rect 30190 26772 30196 26784
rect 30151 26744 30196 26772
rect 30190 26732 30196 26744
rect 30248 26732 30254 26784
rect 35894 26732 35900 26784
rect 35952 26772 35958 26784
rect 36173 26775 36231 26781
rect 36173 26772 36185 26775
rect 35952 26744 36185 26772
rect 35952 26732 35958 26744
rect 36173 26741 36185 26744
rect 36219 26741 36231 26775
rect 36173 26735 36231 26741
rect 1104 26682 54372 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 54372 26682
rect 1104 26608 54372 26630
rect 22097 26571 22155 26577
rect 22097 26537 22109 26571
rect 22143 26568 22155 26571
rect 22186 26568 22192 26580
rect 22143 26540 22192 26568
rect 22143 26537 22155 26540
rect 22097 26531 22155 26537
rect 22186 26528 22192 26540
rect 22244 26528 22250 26580
rect 24486 26568 24492 26580
rect 24447 26540 24492 26568
rect 24486 26528 24492 26540
rect 24544 26528 24550 26580
rect 25958 26568 25964 26580
rect 25919 26540 25964 26568
rect 25958 26528 25964 26540
rect 26016 26528 26022 26580
rect 27614 26568 27620 26580
rect 27575 26540 27620 26568
rect 27614 26528 27620 26540
rect 27672 26528 27678 26580
rect 28074 26528 28080 26580
rect 28132 26568 28138 26580
rect 28169 26571 28227 26577
rect 28169 26568 28181 26571
rect 28132 26540 28181 26568
rect 28132 26528 28138 26540
rect 28169 26537 28181 26540
rect 28215 26537 28227 26571
rect 28169 26531 28227 26537
rect 28997 26571 29055 26577
rect 28997 26537 29009 26571
rect 29043 26568 29055 26571
rect 30190 26568 30196 26580
rect 29043 26540 30196 26568
rect 29043 26537 29055 26540
rect 28997 26531 29055 26537
rect 30190 26528 30196 26540
rect 30248 26568 30254 26580
rect 30377 26571 30435 26577
rect 30377 26568 30389 26571
rect 30248 26540 30389 26568
rect 30248 26528 30254 26540
rect 30377 26537 30389 26540
rect 30423 26537 30435 26571
rect 30377 26531 30435 26537
rect 30745 26571 30803 26577
rect 30745 26537 30757 26571
rect 30791 26568 30803 26571
rect 31294 26568 31300 26580
rect 30791 26540 31300 26568
rect 30791 26537 30803 26540
rect 30745 26531 30803 26537
rect 31294 26528 31300 26540
rect 31352 26528 31358 26580
rect 31662 26528 31668 26580
rect 31720 26568 31726 26580
rect 32493 26571 32551 26577
rect 31720 26540 31984 26568
rect 31720 26528 31726 26540
rect 20441 26503 20499 26509
rect 20441 26469 20453 26503
rect 20487 26500 20499 26503
rect 21450 26500 21456 26512
rect 20487 26472 21456 26500
rect 20487 26469 20499 26472
rect 20441 26463 20499 26469
rect 21450 26460 21456 26472
rect 21508 26460 21514 26512
rect 22741 26503 22799 26509
rect 22741 26469 22753 26503
rect 22787 26500 22799 26503
rect 22787 26472 27660 26500
rect 22787 26469 22799 26472
rect 22741 26463 22799 26469
rect 19334 26392 19340 26444
rect 19392 26432 19398 26444
rect 19981 26435 20039 26441
rect 19981 26432 19993 26435
rect 19392 26404 19993 26432
rect 19392 26392 19398 26404
rect 19981 26401 19993 26404
rect 20027 26432 20039 26435
rect 20162 26432 20168 26444
rect 20027 26404 20168 26432
rect 20027 26401 20039 26404
rect 19981 26395 20039 26401
rect 20162 26392 20168 26404
rect 20220 26392 20226 26444
rect 21726 26392 21732 26444
rect 21784 26432 21790 26444
rect 21913 26435 21971 26441
rect 21913 26432 21925 26435
rect 21784 26404 21925 26432
rect 21784 26392 21790 26404
rect 21913 26401 21925 26404
rect 21959 26401 21971 26435
rect 21913 26395 21971 26401
rect 25501 26435 25559 26441
rect 25501 26401 25513 26435
rect 25547 26432 25559 26435
rect 25866 26432 25872 26444
rect 25547 26404 25872 26432
rect 25547 26401 25559 26404
rect 25501 26395 25559 26401
rect 20070 26364 20076 26376
rect 20031 26336 20076 26364
rect 20070 26324 20076 26336
rect 20128 26324 20134 26376
rect 21821 26367 21879 26373
rect 21821 26333 21833 26367
rect 21867 26333 21879 26367
rect 21928 26364 21956 26395
rect 25866 26392 25872 26404
rect 25924 26392 25930 26444
rect 26142 26432 26148 26444
rect 26103 26404 26148 26432
rect 26142 26392 26148 26404
rect 26200 26392 26206 26444
rect 26418 26432 26424 26444
rect 26379 26404 26424 26432
rect 26418 26392 26424 26404
rect 26476 26392 26482 26444
rect 27154 26432 27160 26444
rect 26988 26404 27160 26432
rect 22649 26367 22707 26373
rect 22649 26364 22661 26367
rect 21928 26336 22661 26364
rect 21821 26327 21879 26333
rect 22649 26333 22661 26336
rect 22695 26333 22707 26367
rect 22649 26327 22707 26333
rect 22833 26367 22891 26373
rect 22833 26333 22845 26367
rect 22879 26333 22891 26367
rect 24394 26364 24400 26376
rect 24355 26336 24400 26364
rect 22833 26327 22891 26333
rect 21836 26296 21864 26327
rect 22462 26296 22468 26308
rect 21836 26268 22468 26296
rect 22462 26256 22468 26268
rect 22520 26296 22526 26308
rect 22848 26296 22876 26327
rect 24394 26324 24400 26336
rect 24452 26324 24458 26376
rect 24581 26367 24639 26373
rect 24581 26333 24593 26367
rect 24627 26364 24639 26367
rect 24854 26364 24860 26376
rect 24627 26336 24860 26364
rect 24627 26333 24639 26336
rect 24581 26327 24639 26333
rect 24854 26324 24860 26336
rect 24912 26324 24918 26376
rect 25406 26324 25412 26376
rect 25464 26364 25470 26376
rect 26050 26364 26056 26376
rect 25464 26336 26056 26364
rect 25464 26324 25470 26336
rect 26050 26324 26056 26336
rect 26108 26364 26114 26376
rect 26237 26367 26295 26373
rect 26237 26364 26249 26367
rect 26108 26336 26249 26364
rect 26108 26324 26114 26336
rect 26237 26333 26249 26336
rect 26283 26333 26295 26367
rect 26237 26327 26295 26333
rect 23750 26296 23756 26308
rect 22520 26268 22876 26296
rect 23711 26268 23756 26296
rect 22520 26256 22526 26268
rect 23750 26256 23756 26268
rect 23808 26256 23814 26308
rect 21082 26228 21088 26240
rect 21043 26200 21088 26228
rect 21082 26188 21088 26200
rect 21140 26188 21146 26240
rect 26252 26228 26280 26327
rect 26326 26324 26332 26376
rect 26384 26364 26390 26376
rect 26988 26373 27016 26404
rect 27154 26392 27160 26404
rect 27212 26392 27218 26444
rect 26973 26367 27031 26373
rect 26384 26336 26429 26364
rect 26384 26324 26390 26336
rect 26973 26333 26985 26367
rect 27019 26333 27031 26367
rect 26973 26327 27031 26333
rect 27062 26324 27068 26376
rect 27120 26364 27126 26376
rect 27448 26367 27506 26373
rect 27120 26336 27165 26364
rect 27120 26324 27126 26336
rect 27448 26333 27460 26367
rect 27494 26364 27506 26367
rect 27632 26364 27660 26472
rect 28258 26460 28264 26512
rect 28316 26500 28322 26512
rect 30650 26500 30656 26512
rect 28316 26472 30656 26500
rect 28316 26460 28322 26472
rect 30650 26460 30656 26472
rect 30708 26460 30714 26512
rect 27798 26392 27804 26444
rect 27856 26432 27862 26444
rect 27856 26404 28304 26432
rect 27856 26392 27862 26404
rect 28276 26373 28304 26404
rect 30190 26392 30196 26444
rect 30248 26432 30254 26444
rect 30469 26435 30527 26441
rect 30469 26432 30481 26435
rect 30248 26404 30481 26432
rect 30248 26392 30254 26404
rect 30469 26401 30481 26404
rect 30515 26401 30527 26435
rect 30469 26395 30527 26401
rect 28077 26367 28135 26373
rect 28077 26364 28089 26367
rect 27494 26336 27568 26364
rect 27632 26336 28089 26364
rect 27494 26333 27506 26336
rect 27448 26327 27506 26333
rect 26344 26296 26372 26324
rect 27249 26299 27307 26305
rect 27249 26296 27261 26299
rect 26344 26268 27261 26296
rect 27249 26265 27261 26268
rect 27295 26265 27307 26299
rect 27249 26259 27307 26265
rect 27341 26299 27399 26305
rect 27341 26265 27353 26299
rect 27387 26265 27399 26299
rect 27540 26296 27568 26336
rect 28077 26333 28089 26336
rect 28123 26333 28135 26367
rect 28077 26327 28135 26333
rect 28261 26367 28319 26373
rect 28261 26333 28273 26367
rect 28307 26364 28319 26367
rect 28721 26367 28779 26373
rect 28721 26364 28733 26367
rect 28307 26336 28733 26364
rect 28307 26333 28319 26336
rect 28261 26327 28319 26333
rect 28721 26333 28733 26336
rect 28767 26333 28779 26367
rect 28721 26327 28779 26333
rect 28997 26367 29055 26373
rect 28997 26333 29009 26367
rect 29043 26364 29055 26367
rect 29270 26364 29276 26376
rect 29043 26336 29276 26364
rect 29043 26333 29055 26336
rect 28997 26327 29055 26333
rect 27614 26296 27620 26308
rect 27540 26268 27620 26296
rect 27341 26259 27399 26265
rect 27356 26228 27384 26259
rect 27614 26256 27620 26268
rect 27672 26256 27678 26308
rect 28092 26296 28120 26327
rect 29270 26324 29276 26336
rect 29328 26324 29334 26376
rect 29638 26324 29644 26376
rect 29696 26364 29702 26376
rect 29917 26367 29975 26373
rect 29917 26364 29929 26367
rect 29696 26336 29929 26364
rect 29696 26324 29702 26336
rect 29917 26333 29929 26336
rect 29963 26333 29975 26367
rect 30374 26364 30380 26376
rect 30335 26336 30380 26364
rect 29917 26327 29975 26333
rect 30374 26324 30380 26336
rect 30432 26324 30438 26376
rect 31205 26367 31263 26373
rect 31205 26364 31217 26367
rect 30576 26336 31217 26364
rect 28813 26299 28871 26305
rect 28813 26296 28825 26299
rect 28092 26268 28825 26296
rect 28813 26265 28825 26268
rect 28859 26265 28871 26299
rect 29730 26296 29736 26308
rect 29691 26268 29736 26296
rect 28813 26259 28871 26265
rect 29730 26256 29736 26268
rect 29788 26256 29794 26308
rect 29546 26228 29552 26240
rect 26252 26200 27384 26228
rect 29507 26200 29552 26228
rect 29546 26188 29552 26200
rect 29604 26188 29610 26240
rect 29748 26228 29776 26256
rect 30576 26228 30604 26336
rect 31205 26333 31217 26336
rect 31251 26333 31263 26367
rect 31386 26364 31392 26376
rect 31347 26336 31392 26364
rect 31205 26327 31263 26333
rect 31220 26296 31248 26327
rect 31386 26324 31392 26336
rect 31444 26364 31450 26376
rect 31956 26373 31984 26540
rect 32493 26537 32505 26571
rect 32539 26568 32551 26571
rect 32766 26568 32772 26580
rect 32539 26540 32772 26568
rect 32539 26537 32551 26540
rect 32493 26531 32551 26537
rect 32766 26528 32772 26540
rect 32824 26528 32830 26580
rect 33778 26528 33784 26580
rect 33836 26568 33842 26580
rect 34057 26571 34115 26577
rect 34057 26568 34069 26571
rect 33836 26540 34069 26568
rect 33836 26528 33842 26540
rect 34057 26537 34069 26540
rect 34103 26537 34115 26571
rect 34057 26531 34115 26537
rect 34054 26392 34060 26444
rect 34112 26432 34118 26444
rect 34793 26435 34851 26441
rect 34793 26432 34805 26435
rect 34112 26404 34805 26432
rect 34112 26392 34118 26404
rect 34793 26401 34805 26404
rect 34839 26432 34851 26435
rect 52822 26432 52828 26444
rect 34839 26404 52828 26432
rect 34839 26401 34851 26404
rect 34793 26395 34851 26401
rect 52822 26392 52828 26404
rect 52880 26392 52886 26444
rect 31941 26367 31999 26373
rect 31444 26336 31892 26364
rect 31444 26324 31450 26336
rect 31754 26296 31760 26308
rect 31220 26268 31760 26296
rect 31754 26256 31760 26268
rect 31812 26256 31818 26308
rect 31864 26296 31892 26336
rect 31941 26333 31953 26367
rect 31987 26364 31999 26367
rect 32953 26367 33011 26373
rect 32953 26364 32965 26367
rect 31987 26336 32965 26364
rect 31987 26333 31999 26336
rect 31941 26327 31999 26333
rect 32953 26333 32965 26336
rect 32999 26333 33011 26367
rect 32953 26327 33011 26333
rect 35342 26324 35348 26376
rect 35400 26364 35406 26376
rect 35621 26367 35679 26373
rect 35621 26364 35633 26367
rect 35400 26336 35633 26364
rect 35400 26324 35406 26336
rect 35621 26333 35633 26336
rect 35667 26364 35679 26367
rect 53374 26364 53380 26376
rect 35667 26336 53380 26364
rect 35667 26333 35679 26336
rect 35621 26327 35679 26333
rect 53374 26324 53380 26336
rect 53432 26324 53438 26376
rect 33318 26296 33324 26308
rect 31864 26268 33324 26296
rect 33318 26256 33324 26268
rect 33376 26296 33382 26308
rect 33597 26299 33655 26305
rect 33597 26296 33609 26299
rect 33376 26268 33609 26296
rect 33376 26256 33382 26268
rect 33597 26265 33609 26268
rect 33643 26296 33655 26299
rect 36078 26296 36084 26308
rect 33643 26268 35940 26296
rect 36039 26268 36084 26296
rect 33643 26265 33655 26268
rect 33597 26259 33655 26265
rect 31294 26228 31300 26240
rect 29748 26200 30604 26228
rect 31255 26200 31300 26228
rect 31294 26188 31300 26200
rect 31352 26188 31358 26240
rect 35912 26228 35940 26268
rect 36078 26256 36084 26268
rect 36136 26256 36142 26308
rect 52454 26296 52460 26308
rect 36188 26268 52460 26296
rect 36188 26228 36216 26268
rect 52454 26256 52460 26268
rect 52512 26256 52518 26308
rect 35912 26200 36216 26228
rect 1104 26138 54372 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 54372 26138
rect 1104 26064 54372 26086
rect 20070 26024 20076 26036
rect 20031 25996 20076 26024
rect 20070 25984 20076 25996
rect 20128 25984 20134 26036
rect 24394 26024 24400 26036
rect 24355 25996 24400 26024
rect 24394 25984 24400 25996
rect 24452 25984 24458 26036
rect 24854 26024 24860 26036
rect 24815 25996 24860 26024
rect 24854 25984 24860 25996
rect 24912 25984 24918 26036
rect 26234 25984 26240 26036
rect 26292 26024 26298 26036
rect 26329 26027 26387 26033
rect 26329 26024 26341 26027
rect 26292 25996 26341 26024
rect 26292 25984 26298 25996
rect 26329 25993 26341 25996
rect 26375 25993 26387 26027
rect 26329 25987 26387 25993
rect 27062 25984 27068 26036
rect 27120 26024 27126 26036
rect 27525 26027 27583 26033
rect 27120 25996 27292 26024
rect 27120 25984 27126 25996
rect 19334 25916 19340 25968
rect 19392 25956 19398 25968
rect 24213 25959 24271 25965
rect 24213 25956 24225 25959
rect 19392 25928 20668 25956
rect 19392 25916 19398 25928
rect 19978 25888 19984 25900
rect 19939 25860 19984 25888
rect 19978 25848 19984 25860
rect 20036 25848 20042 25900
rect 20640 25897 20668 25928
rect 22940 25928 24225 25956
rect 20165 25891 20223 25897
rect 20165 25857 20177 25891
rect 20211 25888 20223 25891
rect 20625 25891 20683 25897
rect 20211 25860 20300 25888
rect 20211 25857 20223 25860
rect 20165 25851 20223 25857
rect 19334 25644 19340 25696
rect 19392 25684 19398 25696
rect 19429 25687 19487 25693
rect 19429 25684 19441 25687
rect 19392 25656 19441 25684
rect 19392 25644 19398 25656
rect 19429 25653 19441 25656
rect 19475 25653 19487 25687
rect 19429 25647 19487 25653
rect 20162 25644 20168 25696
rect 20220 25684 20226 25696
rect 20272 25684 20300 25860
rect 20625 25857 20637 25891
rect 20671 25857 20683 25891
rect 20625 25851 20683 25857
rect 20809 25891 20867 25897
rect 20809 25857 20821 25891
rect 20855 25888 20867 25891
rect 22186 25888 22192 25900
rect 20855 25860 22192 25888
rect 20855 25857 20867 25860
rect 20809 25851 20867 25857
rect 22186 25848 22192 25860
rect 22244 25888 22250 25900
rect 22940 25897 22968 25928
rect 24213 25925 24225 25928
rect 24259 25956 24271 25959
rect 24872 25956 24900 25984
rect 27154 25956 27160 25968
rect 24259 25928 24808 25956
rect 24872 25928 26372 25956
rect 24259 25925 24271 25928
rect 24213 25919 24271 25925
rect 22925 25891 22983 25897
rect 22925 25888 22937 25891
rect 22244 25860 22937 25888
rect 22244 25848 22250 25860
rect 22925 25857 22937 25860
rect 22971 25857 22983 25891
rect 22925 25851 22983 25857
rect 23658 25848 23664 25900
rect 23716 25888 23722 25900
rect 24029 25891 24087 25897
rect 24029 25888 24041 25891
rect 23716 25860 24041 25888
rect 23716 25848 23722 25860
rect 24029 25857 24041 25860
rect 24075 25857 24087 25891
rect 24029 25851 24087 25857
rect 24044 25820 24072 25851
rect 24670 25848 24676 25900
rect 24728 25888 24734 25900
rect 24780 25888 24808 25928
rect 25976 25897 26004 25928
rect 26344 25900 26372 25928
rect 27080 25928 27160 25956
rect 24857 25891 24915 25897
rect 24857 25888 24869 25891
rect 24728 25860 24869 25888
rect 24728 25848 24734 25860
rect 24857 25857 24869 25860
rect 24903 25857 24915 25891
rect 24857 25851 24915 25857
rect 25041 25891 25099 25897
rect 25041 25857 25053 25891
rect 25087 25857 25099 25891
rect 25041 25851 25099 25857
rect 25961 25891 26019 25897
rect 25961 25857 25973 25891
rect 26007 25857 26019 25891
rect 25961 25851 26019 25857
rect 24578 25820 24584 25832
rect 24044 25792 24584 25820
rect 24578 25780 24584 25792
rect 24636 25820 24642 25832
rect 25056 25820 25084 25851
rect 26050 25848 26056 25900
rect 26108 25888 26114 25900
rect 26145 25891 26203 25897
rect 26145 25888 26157 25891
rect 26108 25860 26157 25888
rect 26108 25848 26114 25860
rect 26145 25857 26157 25860
rect 26191 25857 26203 25891
rect 26145 25851 26203 25857
rect 24636 25792 25084 25820
rect 24636 25780 24642 25792
rect 23569 25755 23627 25761
rect 23569 25721 23581 25755
rect 23615 25752 23627 25755
rect 25682 25752 25688 25764
rect 23615 25724 25688 25752
rect 23615 25721 23627 25724
rect 23569 25715 23627 25721
rect 25682 25712 25688 25724
rect 25740 25712 25746 25764
rect 26160 25752 26188 25851
rect 26326 25848 26332 25900
rect 26384 25848 26390 25900
rect 27080 25897 27108 25928
rect 27154 25916 27160 25928
rect 27212 25916 27218 25968
rect 27264 25956 27292 25996
rect 27525 25993 27537 26027
rect 27571 26024 27583 26027
rect 27890 26024 27896 26036
rect 27571 25996 27896 26024
rect 27571 25993 27583 25996
rect 27525 25987 27583 25993
rect 27890 25984 27896 25996
rect 27948 25984 27954 26036
rect 27982 25984 27988 26036
rect 28040 26024 28046 26036
rect 28721 26027 28779 26033
rect 28721 26024 28733 26027
rect 28040 25996 28733 26024
rect 28040 25984 28046 25996
rect 28721 25993 28733 25996
rect 28767 25993 28779 26027
rect 30190 26024 30196 26036
rect 30151 25996 30196 26024
rect 28721 25987 28779 25993
rect 30190 25984 30196 25996
rect 30248 25984 30254 26036
rect 32766 26024 32772 26036
rect 32727 25996 32772 26024
rect 32766 25984 32772 25996
rect 32824 25984 32830 26036
rect 33318 26024 33324 26036
rect 33279 25996 33324 26024
rect 33318 25984 33324 25996
rect 33376 25984 33382 26036
rect 33778 26024 33784 26036
rect 33739 25996 33784 26024
rect 33778 25984 33784 25996
rect 33836 25984 33842 26036
rect 34330 26024 34336 26036
rect 34291 25996 34336 26024
rect 34330 25984 34336 25996
rect 34388 25984 34394 26036
rect 28000 25956 28028 25984
rect 27264 25928 28028 25956
rect 29362 25916 29368 25968
rect 29420 25956 29426 25968
rect 29638 25956 29644 25968
rect 29420 25928 29644 25956
rect 29420 25916 29426 25928
rect 29638 25916 29644 25928
rect 29696 25956 29702 25968
rect 31021 25959 31079 25965
rect 29696 25928 29868 25956
rect 29696 25916 29702 25928
rect 27065 25891 27123 25897
rect 27065 25857 27077 25891
rect 27111 25857 27123 25891
rect 27065 25851 27123 25857
rect 27430 25848 27436 25900
rect 27488 25888 27494 25900
rect 27985 25891 28043 25897
rect 27985 25888 27997 25891
rect 27488 25860 27997 25888
rect 27488 25848 27494 25860
rect 27985 25857 27997 25860
rect 28031 25857 28043 25891
rect 27985 25851 28043 25857
rect 28721 25891 28779 25897
rect 28721 25857 28733 25891
rect 28767 25857 28779 25891
rect 28721 25851 28779 25857
rect 28905 25891 28963 25897
rect 28905 25857 28917 25891
rect 28951 25888 28963 25891
rect 29546 25888 29552 25900
rect 28951 25860 29552 25888
rect 28951 25857 28963 25860
rect 28905 25851 28963 25857
rect 26344 25820 26372 25848
rect 27157 25823 27215 25829
rect 27157 25820 27169 25823
rect 26344 25792 27169 25820
rect 27157 25789 27169 25792
rect 27203 25789 27215 25823
rect 27157 25783 27215 25789
rect 27249 25823 27307 25829
rect 27249 25789 27261 25823
rect 27295 25789 27307 25823
rect 27249 25783 27307 25789
rect 27264 25752 27292 25783
rect 27338 25780 27344 25832
rect 27396 25820 27402 25832
rect 27614 25820 27620 25832
rect 27396 25792 27620 25820
rect 27396 25780 27402 25792
rect 27614 25780 27620 25792
rect 27672 25780 27678 25832
rect 28736 25820 28764 25851
rect 29546 25848 29552 25860
rect 29604 25848 29610 25900
rect 29840 25897 29868 25928
rect 31021 25925 31033 25959
rect 31067 25956 31079 25959
rect 31067 25928 31754 25956
rect 31067 25925 31079 25928
rect 31021 25919 31079 25925
rect 31726 25900 31754 25928
rect 29825 25891 29883 25897
rect 29825 25857 29837 25891
rect 29871 25857 29883 25891
rect 30006 25888 30012 25900
rect 29967 25860 30012 25888
rect 29825 25851 29883 25857
rect 29178 25820 29184 25832
rect 28736 25792 29184 25820
rect 29178 25780 29184 25792
rect 29236 25820 29242 25832
rect 29638 25820 29644 25832
rect 29236 25792 29644 25820
rect 29236 25780 29242 25792
rect 29638 25780 29644 25792
rect 29696 25780 29702 25832
rect 26160 25724 27292 25752
rect 29840 25752 29868 25851
rect 30006 25848 30012 25860
rect 30064 25848 30070 25900
rect 31205 25891 31263 25897
rect 31205 25857 31217 25891
rect 31251 25888 31263 25891
rect 31386 25888 31392 25900
rect 31251 25860 31392 25888
rect 31251 25857 31263 25860
rect 31205 25851 31263 25857
rect 31386 25848 31392 25860
rect 31444 25848 31450 25900
rect 31726 25860 31760 25900
rect 31754 25848 31760 25860
rect 31812 25888 31818 25900
rect 32766 25888 32772 25900
rect 31812 25860 32772 25888
rect 31812 25848 31818 25860
rect 32766 25848 32772 25860
rect 32824 25848 32830 25900
rect 29840 25724 31754 25752
rect 20717 25687 20775 25693
rect 20717 25684 20729 25687
rect 20220 25656 20729 25684
rect 20220 25644 20226 25656
rect 20717 25653 20729 25656
rect 20763 25653 20775 25687
rect 20717 25647 20775 25653
rect 21082 25644 21088 25696
rect 21140 25684 21146 25696
rect 21821 25687 21879 25693
rect 21821 25684 21833 25687
rect 21140 25656 21833 25684
rect 21140 25644 21146 25656
rect 21821 25653 21833 25656
rect 21867 25653 21879 25687
rect 22462 25684 22468 25696
rect 22423 25656 22468 25684
rect 21821 25647 21879 25653
rect 22462 25644 22468 25656
rect 22520 25644 22526 25696
rect 30466 25644 30472 25696
rect 30524 25684 30530 25696
rect 30837 25687 30895 25693
rect 30837 25684 30849 25687
rect 30524 25656 30849 25684
rect 30524 25644 30530 25656
rect 30837 25653 30849 25656
rect 30883 25653 30895 25687
rect 31726 25684 31754 25724
rect 32214 25684 32220 25696
rect 31726 25656 32220 25684
rect 30837 25647 30895 25653
rect 32214 25644 32220 25656
rect 32272 25644 32278 25696
rect 1104 25594 54372 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 54372 25594
rect 1104 25520 54372 25542
rect 19981 25483 20039 25489
rect 19981 25449 19993 25483
rect 20027 25480 20039 25483
rect 21177 25483 21235 25489
rect 20027 25452 20576 25480
rect 20027 25449 20039 25452
rect 19981 25443 20039 25449
rect 20070 25412 20076 25424
rect 19720 25384 20076 25412
rect 19720 25285 19748 25384
rect 20070 25372 20076 25384
rect 20128 25372 20134 25424
rect 20162 25344 20168 25356
rect 20123 25316 20168 25344
rect 20162 25304 20168 25316
rect 20220 25304 20226 25356
rect 20548 25344 20576 25452
rect 21177 25449 21189 25483
rect 21223 25480 21235 25483
rect 21726 25480 21732 25492
rect 21223 25452 21732 25480
rect 21223 25449 21235 25452
rect 21177 25443 21235 25449
rect 21726 25440 21732 25452
rect 21784 25440 21790 25492
rect 24670 25480 24676 25492
rect 24631 25452 24676 25480
rect 24670 25440 24676 25452
rect 24728 25440 24734 25492
rect 25590 25440 25596 25492
rect 25648 25480 25654 25492
rect 25777 25483 25835 25489
rect 25777 25480 25789 25483
rect 25648 25452 25789 25480
rect 25648 25440 25654 25452
rect 25777 25449 25789 25452
rect 25823 25449 25835 25483
rect 27154 25480 27160 25492
rect 27115 25452 27160 25480
rect 25777 25443 25835 25449
rect 27154 25440 27160 25452
rect 27212 25440 27218 25492
rect 28997 25483 29055 25489
rect 28997 25449 29009 25483
rect 29043 25480 29055 25483
rect 29270 25480 29276 25492
rect 29043 25452 29276 25480
rect 29043 25449 29055 25452
rect 28997 25443 29055 25449
rect 29270 25440 29276 25452
rect 29328 25440 29334 25492
rect 29638 25480 29644 25492
rect 29599 25452 29644 25480
rect 29638 25440 29644 25452
rect 29696 25440 29702 25492
rect 32033 25483 32091 25489
rect 32033 25449 32045 25483
rect 32079 25480 32091 25483
rect 32214 25480 32220 25492
rect 32079 25452 32220 25480
rect 32079 25449 32091 25452
rect 32033 25443 32091 25449
rect 32214 25440 32220 25452
rect 32272 25480 32278 25492
rect 51442 25480 51448 25492
rect 32272 25452 51448 25480
rect 32272 25440 32278 25452
rect 51442 25440 51448 25452
rect 51500 25440 51506 25492
rect 52822 25480 52828 25492
rect 52783 25452 52828 25480
rect 52822 25440 52828 25452
rect 52880 25440 52886 25492
rect 26421 25415 26479 25421
rect 26421 25381 26433 25415
rect 26467 25412 26479 25415
rect 27338 25412 27344 25424
rect 26467 25384 27344 25412
rect 26467 25381 26479 25384
rect 26421 25375 26479 25381
rect 27338 25372 27344 25384
rect 27396 25372 27402 25424
rect 32585 25415 32643 25421
rect 32585 25381 32597 25415
rect 32631 25412 32643 25415
rect 32766 25412 32772 25424
rect 32631 25384 32772 25412
rect 32631 25381 32643 25384
rect 32585 25375 32643 25381
rect 32766 25372 32772 25384
rect 32824 25372 32830 25424
rect 20717 25347 20775 25353
rect 20717 25344 20729 25347
rect 20548 25316 20729 25344
rect 20717 25313 20729 25316
rect 20763 25344 20775 25347
rect 20898 25344 20904 25356
rect 20763 25316 20904 25344
rect 20763 25313 20775 25316
rect 20717 25307 20775 25313
rect 20898 25304 20904 25316
rect 20956 25304 20962 25356
rect 26602 25344 26608 25356
rect 26344 25316 26608 25344
rect 26344 25288 26372 25316
rect 26602 25304 26608 25316
rect 26660 25344 26666 25356
rect 27617 25347 27675 25353
rect 27617 25344 27629 25347
rect 26660 25316 27629 25344
rect 26660 25304 26666 25316
rect 19705 25279 19763 25285
rect 19705 25245 19717 25279
rect 19751 25245 19763 25279
rect 19705 25239 19763 25245
rect 19797 25279 19855 25285
rect 19797 25245 19809 25279
rect 19843 25276 19855 25279
rect 19978 25276 19984 25288
rect 19843 25248 19984 25276
rect 19843 25245 19855 25248
rect 19797 25239 19855 25245
rect 19978 25236 19984 25248
rect 20036 25236 20042 25288
rect 20806 25276 20812 25288
rect 20767 25248 20812 25276
rect 20806 25236 20812 25248
rect 20864 25236 20870 25288
rect 26326 25276 26332 25288
rect 25148 25248 26332 25276
rect 1854 25208 1860 25220
rect 1815 25180 1860 25208
rect 1854 25168 1860 25180
rect 1912 25168 1918 25220
rect 1949 25143 2007 25149
rect 1949 25109 1961 25143
rect 1995 25140 2007 25143
rect 16482 25140 16488 25152
rect 1995 25112 16488 25140
rect 1995 25109 2007 25112
rect 1949 25103 2007 25109
rect 16482 25100 16488 25112
rect 16540 25100 16546 25152
rect 21729 25143 21787 25149
rect 21729 25109 21741 25143
rect 21775 25140 21787 25143
rect 22186 25140 22192 25152
rect 21775 25112 22192 25140
rect 21775 25109 21787 25112
rect 21729 25103 21787 25109
rect 22186 25100 22192 25112
rect 22244 25100 22250 25152
rect 22462 25100 22468 25152
rect 22520 25140 22526 25152
rect 22925 25143 22983 25149
rect 22925 25140 22937 25143
rect 22520 25112 22937 25140
rect 22520 25100 22526 25112
rect 22925 25109 22937 25112
rect 22971 25140 22983 25143
rect 24486 25140 24492 25152
rect 22971 25112 24492 25140
rect 22971 25109 22983 25112
rect 22925 25103 22983 25109
rect 24486 25100 24492 25112
rect 24544 25140 24550 25152
rect 25148 25149 25176 25248
rect 26326 25236 26332 25248
rect 26384 25236 26390 25288
rect 27172 25285 27200 25316
rect 27617 25313 27629 25316
rect 27663 25313 27675 25347
rect 30006 25344 30012 25356
rect 27617 25307 27675 25313
rect 29012 25316 30012 25344
rect 29012 25285 29040 25316
rect 30006 25304 30012 25316
rect 30064 25304 30070 25356
rect 30466 25344 30472 25356
rect 30427 25316 30472 25344
rect 30466 25304 30472 25316
rect 30524 25344 30530 25356
rect 30524 25316 31524 25344
rect 30524 25304 30530 25316
rect 26513 25279 26571 25285
rect 26513 25245 26525 25279
rect 26559 25276 26571 25279
rect 26973 25279 27031 25285
rect 26973 25276 26985 25279
rect 26559 25248 26985 25276
rect 26559 25245 26571 25248
rect 26513 25239 26571 25245
rect 26973 25245 26985 25248
rect 27019 25245 27031 25279
rect 26973 25239 27031 25245
rect 27157 25279 27215 25285
rect 27157 25245 27169 25279
rect 27203 25245 27215 25279
rect 27157 25239 27215 25245
rect 28813 25279 28871 25285
rect 28813 25245 28825 25279
rect 28859 25245 28871 25279
rect 28813 25239 28871 25245
rect 28997 25279 29055 25285
rect 28997 25245 29009 25279
rect 29043 25245 29055 25279
rect 28997 25239 29055 25245
rect 26988 25208 27016 25239
rect 27614 25208 27620 25220
rect 26988 25180 27620 25208
rect 27614 25168 27620 25180
rect 27672 25168 27678 25220
rect 28828 25208 28856 25239
rect 29362 25236 29368 25288
rect 29420 25276 29426 25288
rect 29549 25279 29607 25285
rect 29549 25276 29561 25279
rect 29420 25248 29561 25276
rect 29420 25236 29426 25248
rect 29549 25245 29561 25248
rect 29595 25245 29607 25279
rect 29730 25276 29736 25288
rect 29691 25248 29736 25276
rect 29549 25239 29607 25245
rect 29730 25236 29736 25248
rect 29788 25236 29794 25288
rect 30377 25279 30435 25285
rect 30377 25245 30389 25279
rect 30423 25245 30435 25279
rect 30377 25239 30435 25245
rect 30837 25279 30895 25285
rect 30837 25245 30849 25279
rect 30883 25276 30895 25279
rect 31294 25276 31300 25288
rect 30883 25248 31300 25276
rect 30883 25245 30895 25248
rect 30837 25239 30895 25245
rect 29380 25208 29408 25236
rect 28828 25180 29408 25208
rect 30392 25208 30420 25239
rect 31294 25236 31300 25248
rect 31352 25236 31358 25288
rect 31496 25285 31524 25316
rect 31481 25279 31539 25285
rect 31481 25245 31493 25279
rect 31527 25245 31539 25279
rect 31481 25239 31539 25245
rect 52822 25236 52828 25288
rect 52880 25276 52886 25288
rect 53377 25279 53435 25285
rect 53377 25276 53389 25279
rect 52880 25248 53389 25276
rect 52880 25236 52886 25248
rect 53377 25245 53389 25248
rect 53423 25245 53435 25279
rect 53377 25239 53435 25245
rect 30466 25208 30472 25220
rect 30392 25180 30472 25208
rect 30466 25168 30472 25180
rect 30524 25168 30530 25220
rect 25133 25143 25191 25149
rect 25133 25140 25145 25143
rect 24544 25112 25145 25140
rect 24544 25100 24550 25112
rect 25133 25109 25145 25112
rect 25179 25109 25191 25143
rect 28258 25140 28264 25152
rect 28219 25112 28264 25140
rect 25133 25103 25191 25109
rect 28258 25100 28264 25112
rect 28316 25100 28322 25152
rect 30193 25143 30251 25149
rect 30193 25109 30205 25143
rect 30239 25140 30251 25143
rect 30742 25140 30748 25152
rect 30239 25112 30748 25140
rect 30239 25109 30251 25112
rect 30193 25103 30251 25109
rect 30742 25100 30748 25112
rect 30800 25100 30806 25152
rect 31294 25140 31300 25152
rect 31255 25112 31300 25140
rect 31294 25100 31300 25112
rect 31352 25100 31358 25152
rect 53558 25140 53564 25152
rect 53519 25112 53564 25140
rect 53558 25100 53564 25112
rect 53616 25100 53622 25152
rect 1104 25050 54372 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 54372 25050
rect 1104 24976 54372 24998
rect 1673 24939 1731 24945
rect 1673 24905 1685 24939
rect 1719 24936 1731 24939
rect 1854 24936 1860 24948
rect 1719 24908 1860 24936
rect 1719 24905 1731 24908
rect 1673 24899 1731 24905
rect 1854 24896 1860 24908
rect 1912 24896 1918 24948
rect 19889 24939 19947 24945
rect 19889 24905 19901 24939
rect 19935 24936 19947 24939
rect 19978 24936 19984 24948
rect 19935 24908 19984 24936
rect 19935 24905 19947 24908
rect 19889 24899 19947 24905
rect 19978 24896 19984 24908
rect 20036 24896 20042 24948
rect 20806 24896 20812 24948
rect 20864 24936 20870 24948
rect 21821 24939 21879 24945
rect 21821 24936 21833 24939
rect 20864 24908 21833 24936
rect 20864 24896 20870 24908
rect 21821 24905 21833 24908
rect 21867 24905 21879 24939
rect 24578 24936 24584 24948
rect 24539 24908 24584 24936
rect 21821 24899 21879 24905
rect 24578 24896 24584 24908
rect 24636 24936 24642 24948
rect 25133 24939 25191 24945
rect 25133 24936 25145 24939
rect 24636 24908 25145 24936
rect 24636 24896 24642 24908
rect 25133 24905 25145 24908
rect 25179 24905 25191 24939
rect 25133 24899 25191 24905
rect 25682 24896 25688 24948
rect 25740 24936 25746 24948
rect 25961 24939 26019 24945
rect 25961 24936 25973 24939
rect 25740 24908 25973 24936
rect 25740 24896 25746 24908
rect 25961 24905 25973 24908
rect 26007 24905 26019 24939
rect 25961 24899 26019 24905
rect 29181 24939 29239 24945
rect 29181 24905 29193 24939
rect 29227 24936 29239 24939
rect 29362 24936 29368 24948
rect 29227 24908 29368 24936
rect 29227 24905 29239 24908
rect 29181 24899 29239 24905
rect 29362 24896 29368 24908
rect 29420 24896 29426 24948
rect 29641 24939 29699 24945
rect 29641 24905 29653 24939
rect 29687 24936 29699 24939
rect 30006 24936 30012 24948
rect 29687 24908 30012 24936
rect 29687 24905 29699 24908
rect 29641 24899 29699 24905
rect 30006 24896 30012 24908
rect 30064 24896 30070 24948
rect 32217 24939 32275 24945
rect 32217 24905 32229 24939
rect 32263 24936 32275 24939
rect 32766 24936 32772 24948
rect 32263 24908 32772 24936
rect 32263 24905 32275 24908
rect 32217 24899 32275 24905
rect 32766 24896 32772 24908
rect 32824 24896 32830 24948
rect 20714 24868 20720 24880
rect 20180 24840 20720 24868
rect 20073 24803 20131 24809
rect 20073 24769 20085 24803
rect 20119 24800 20131 24803
rect 20180 24800 20208 24840
rect 20714 24828 20720 24840
rect 20772 24868 20778 24880
rect 22186 24868 22192 24880
rect 20772 24840 22192 24868
rect 20772 24828 20778 24840
rect 22186 24828 22192 24840
rect 22244 24828 22250 24880
rect 30466 24868 30472 24880
rect 29932 24840 30472 24868
rect 20119 24772 20208 24800
rect 20257 24803 20315 24809
rect 20119 24769 20131 24772
rect 20073 24763 20131 24769
rect 20257 24769 20269 24803
rect 20303 24769 20315 24803
rect 20898 24800 20904 24812
rect 20859 24772 20904 24800
rect 20257 24763 20315 24769
rect 20272 24732 20300 24763
rect 20898 24760 20904 24772
rect 20956 24760 20962 24812
rect 21266 24800 21272 24812
rect 21227 24772 21272 24800
rect 21266 24760 21272 24772
rect 21324 24800 21330 24812
rect 21821 24803 21879 24809
rect 21821 24800 21833 24803
rect 21324 24772 21833 24800
rect 21324 24760 21330 24772
rect 21821 24769 21833 24772
rect 21867 24769 21879 24803
rect 22002 24800 22008 24812
rect 21963 24772 22008 24800
rect 21821 24763 21879 24769
rect 22002 24760 22008 24772
rect 22060 24760 22066 24812
rect 27065 24803 27123 24809
rect 27065 24769 27077 24803
rect 27111 24800 27123 24803
rect 28258 24800 28264 24812
rect 27111 24772 28264 24800
rect 27111 24769 27123 24772
rect 27065 24763 27123 24769
rect 28258 24760 28264 24772
rect 28316 24760 28322 24812
rect 19352 24704 20300 24732
rect 21085 24735 21143 24741
rect 19352 24608 19380 24704
rect 21085 24701 21097 24735
rect 21131 24732 21143 24735
rect 21358 24732 21364 24744
rect 21131 24704 21364 24732
rect 21131 24701 21143 24704
rect 21085 24695 21143 24701
rect 21358 24692 21364 24704
rect 21416 24692 21422 24744
rect 29932 24741 29960 24840
rect 30466 24828 30472 24840
rect 30524 24828 30530 24880
rect 31294 24868 31300 24880
rect 30668 24840 31300 24868
rect 30009 24803 30067 24809
rect 30009 24769 30021 24803
rect 30055 24800 30067 24803
rect 30668 24800 30696 24840
rect 31294 24828 31300 24840
rect 31352 24828 31358 24880
rect 30055 24772 30696 24800
rect 30055 24769 30067 24772
rect 30009 24763 30067 24769
rect 30742 24760 30748 24812
rect 30800 24800 30806 24812
rect 31021 24803 31079 24809
rect 31021 24800 31033 24803
rect 30800 24772 31033 24800
rect 30800 24760 30806 24772
rect 31021 24769 31033 24772
rect 31067 24769 31079 24803
rect 31021 24763 31079 24769
rect 29917 24735 29975 24741
rect 29917 24701 29929 24735
rect 29963 24701 29975 24735
rect 29917 24695 29975 24701
rect 21177 24667 21235 24673
rect 21177 24633 21189 24667
rect 21223 24664 21235 24667
rect 29932 24664 29960 24695
rect 30466 24692 30472 24744
rect 30524 24732 30530 24744
rect 30929 24735 30987 24741
rect 30929 24732 30941 24735
rect 30524 24704 30941 24732
rect 30524 24692 30530 24704
rect 30929 24701 30941 24704
rect 30975 24701 30987 24735
rect 30929 24695 30987 24701
rect 21223 24636 29960 24664
rect 21223 24633 21235 24636
rect 21177 24627 21235 24633
rect 30374 24624 30380 24676
rect 30432 24664 30438 24676
rect 30653 24667 30711 24673
rect 30653 24664 30665 24667
rect 30432 24636 30665 24664
rect 30432 24624 30438 24636
rect 30653 24633 30665 24636
rect 30699 24633 30711 24667
rect 30653 24627 30711 24633
rect 19334 24596 19340 24608
rect 19295 24568 19340 24596
rect 19334 24556 19340 24568
rect 19392 24556 19398 24608
rect 27614 24596 27620 24608
rect 27527 24568 27620 24596
rect 27614 24556 27620 24568
rect 27672 24596 27678 24608
rect 28074 24596 28080 24608
rect 27672 24568 28080 24596
rect 27672 24556 27678 24568
rect 28074 24556 28080 24568
rect 28132 24556 28138 24608
rect 1104 24506 54372 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 54372 24506
rect 1104 24432 54372 24454
rect 20073 24395 20131 24401
rect 20073 24361 20085 24395
rect 20119 24392 20131 24395
rect 20714 24392 20720 24404
rect 20119 24364 20720 24392
rect 20119 24361 20131 24364
rect 20073 24355 20131 24361
rect 20714 24352 20720 24364
rect 20772 24352 20778 24404
rect 21358 24392 21364 24404
rect 21319 24364 21364 24392
rect 21358 24352 21364 24364
rect 21416 24352 21422 24404
rect 26326 24352 26332 24404
rect 26384 24392 26390 24404
rect 26789 24395 26847 24401
rect 26789 24392 26801 24395
rect 26384 24364 26801 24392
rect 26384 24352 26390 24364
rect 26789 24361 26801 24364
rect 26835 24392 26847 24395
rect 27341 24395 27399 24401
rect 27341 24392 27353 24395
rect 26835 24364 27353 24392
rect 26835 24361 26847 24364
rect 26789 24355 26847 24361
rect 27341 24361 27353 24364
rect 27387 24361 27399 24395
rect 30466 24392 30472 24404
rect 30427 24364 30472 24392
rect 27341 24355 27399 24361
rect 30466 24352 30472 24364
rect 30524 24352 30530 24404
rect 20901 24327 20959 24333
rect 20901 24293 20913 24327
rect 20947 24324 20959 24327
rect 22002 24324 22008 24336
rect 20947 24296 22008 24324
rect 20947 24293 20959 24296
rect 20901 24287 20959 24293
rect 22002 24284 22008 24296
rect 22060 24284 22066 24336
rect 22097 24259 22155 24265
rect 22097 24225 22109 24259
rect 22143 24256 22155 24259
rect 22649 24259 22707 24265
rect 22649 24256 22661 24259
rect 22143 24228 22661 24256
rect 22143 24225 22155 24228
rect 22097 24219 22155 24225
rect 22649 24225 22661 24228
rect 22695 24256 22707 24259
rect 27614 24256 27620 24268
rect 22695 24228 27620 24256
rect 22695 24225 22707 24228
rect 22649 24219 22707 24225
rect 21361 24191 21419 24197
rect 21361 24188 21373 24191
rect 20548 24160 21373 24188
rect 20548 24132 20576 24160
rect 21361 24157 21373 24160
rect 21407 24157 21419 24191
rect 21361 24151 21419 24157
rect 21545 24191 21603 24197
rect 21545 24157 21557 24191
rect 21591 24188 21603 24191
rect 22112 24188 22140 24219
rect 27614 24216 27620 24228
rect 27672 24216 27678 24268
rect 30098 24256 30104 24268
rect 30059 24228 30104 24256
rect 30098 24216 30104 24228
rect 30156 24216 30162 24268
rect 21591 24160 22140 24188
rect 30193 24191 30251 24197
rect 21591 24157 21603 24160
rect 21545 24151 21603 24157
rect 30193 24157 30205 24191
rect 30239 24188 30251 24191
rect 30239 24160 30696 24188
rect 30239 24157 30251 24160
rect 30193 24151 30251 24157
rect 19521 24123 19579 24129
rect 19521 24089 19533 24123
rect 19567 24120 19579 24123
rect 20530 24120 20536 24132
rect 19567 24092 20536 24120
rect 19567 24089 19579 24092
rect 19521 24083 19579 24089
rect 20530 24080 20536 24092
rect 20588 24080 20594 24132
rect 20717 24123 20775 24129
rect 20717 24089 20729 24123
rect 20763 24120 20775 24123
rect 20806 24120 20812 24132
rect 20763 24092 20812 24120
rect 20763 24089 20775 24092
rect 20717 24083 20775 24089
rect 20806 24080 20812 24092
rect 20864 24120 20870 24132
rect 21560 24120 21588 24151
rect 20864 24092 21588 24120
rect 20864 24080 20870 24092
rect 30668 24064 30696 24160
rect 30650 24012 30656 24064
rect 30708 24052 30714 24064
rect 31021 24055 31079 24061
rect 31021 24052 31033 24055
rect 30708 24024 31033 24052
rect 30708 24012 30714 24024
rect 31021 24021 31033 24024
rect 31067 24021 31079 24055
rect 31021 24015 31079 24021
rect 1104 23962 54372 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 54372 23962
rect 1104 23888 54372 23910
rect 20809 23851 20867 23857
rect 20809 23817 20821 23851
rect 20855 23848 20867 23851
rect 21266 23848 21272 23860
rect 20855 23820 21272 23848
rect 20855 23817 20867 23820
rect 20809 23811 20867 23817
rect 21266 23808 21272 23820
rect 21324 23808 21330 23860
rect 29362 23808 29368 23860
rect 29420 23848 29426 23860
rect 30009 23851 30067 23857
rect 30009 23848 30021 23851
rect 29420 23820 30021 23848
rect 29420 23808 29426 23820
rect 30009 23817 30021 23820
rect 30055 23817 30067 23851
rect 30009 23811 30067 23817
rect 51718 23808 51724 23860
rect 51776 23848 51782 23860
rect 52825 23851 52883 23857
rect 52825 23848 52837 23851
rect 51776 23820 52837 23848
rect 51776 23808 51782 23820
rect 52825 23817 52837 23820
rect 52871 23817 52883 23851
rect 52825 23811 52883 23817
rect 20530 23712 20536 23724
rect 20088 23684 20536 23712
rect 19978 23468 19984 23520
rect 20036 23508 20042 23520
rect 20088 23517 20116 23684
rect 20530 23672 20536 23684
rect 20588 23712 20594 23724
rect 20625 23715 20683 23721
rect 20625 23712 20637 23715
rect 20588 23684 20637 23712
rect 20588 23672 20594 23684
rect 20625 23681 20637 23684
rect 20671 23681 20683 23715
rect 20806 23712 20812 23724
rect 20767 23684 20812 23712
rect 20625 23675 20683 23681
rect 20640 23644 20668 23675
rect 20806 23672 20812 23684
rect 20864 23672 20870 23724
rect 52840 23712 52868 23811
rect 53377 23715 53435 23721
rect 53377 23712 53389 23715
rect 52840 23684 53389 23712
rect 53377 23681 53389 23684
rect 53423 23681 53435 23715
rect 53377 23675 53435 23681
rect 21821 23647 21879 23653
rect 21821 23644 21833 23647
rect 20640 23616 21833 23644
rect 21821 23613 21833 23616
rect 21867 23613 21879 23647
rect 21821 23607 21879 23613
rect 20073 23511 20131 23517
rect 20073 23508 20085 23511
rect 20036 23480 20085 23508
rect 20036 23468 20042 23480
rect 20073 23477 20085 23480
rect 20119 23477 20131 23511
rect 53558 23508 53564 23520
rect 53519 23480 53564 23508
rect 20073 23471 20131 23477
rect 53558 23468 53564 23480
rect 53616 23468 53622 23520
rect 1104 23418 54372 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 54372 23418
rect 1104 23344 54372 23366
rect 20806 23264 20812 23316
rect 20864 23304 20870 23316
rect 20901 23307 20959 23313
rect 20901 23304 20913 23307
rect 20864 23276 20913 23304
rect 20864 23264 20870 23276
rect 20901 23273 20913 23276
rect 20947 23273 20959 23307
rect 20901 23267 20959 23273
rect 1104 22874 54372 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 54372 22874
rect 1104 22800 54372 22822
rect 1394 22624 1400 22636
rect 1355 22596 1400 22624
rect 1394 22584 1400 22596
rect 1452 22584 1458 22636
rect 1673 22559 1731 22565
rect 1673 22525 1685 22559
rect 1719 22556 1731 22559
rect 34790 22556 34796 22568
rect 1719 22528 34796 22556
rect 1719 22525 1731 22528
rect 1673 22519 1731 22525
rect 34790 22516 34796 22528
rect 34848 22516 34854 22568
rect 1104 22330 54372 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 54372 22330
rect 1104 22256 54372 22278
rect 1394 22216 1400 22228
rect 1355 22188 1400 22216
rect 1394 22176 1400 22188
rect 1452 22176 1458 22228
rect 1104 21786 54372 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 54372 21786
rect 1104 21712 54372 21734
rect 53377 21539 53435 21545
rect 53377 21536 53389 21539
rect 52840 21508 53389 21536
rect 39942 21360 39948 21412
rect 40000 21400 40006 21412
rect 52840 21409 52868 21508
rect 53377 21505 53389 21508
rect 53423 21505 53435 21539
rect 53377 21499 53435 21505
rect 52825 21403 52883 21409
rect 52825 21400 52837 21403
rect 40000 21372 52837 21400
rect 40000 21360 40006 21372
rect 52825 21369 52837 21372
rect 52871 21369 52883 21403
rect 52825 21363 52883 21369
rect 53558 21332 53564 21344
rect 53519 21304 53564 21332
rect 53558 21292 53564 21304
rect 53616 21292 53622 21344
rect 1104 21242 54372 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 54372 21242
rect 1104 21168 54372 21190
rect 1394 20924 1400 20936
rect 1355 20896 1400 20924
rect 1394 20884 1400 20896
rect 1452 20884 1458 20936
rect 1578 20788 1584 20800
rect 1539 20760 1584 20788
rect 1578 20748 1584 20760
rect 1636 20748 1642 20800
rect 1104 20698 54372 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 54372 20698
rect 1104 20624 54372 20646
rect 1394 20516 1400 20528
rect 1355 20488 1400 20516
rect 1394 20476 1400 20488
rect 1452 20476 1458 20528
rect 1104 20154 54372 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 54372 20154
rect 1104 20080 54372 20102
rect 1104 19610 54372 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 54372 19610
rect 1104 19536 54372 19558
rect 1104 19066 54372 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 54372 19066
rect 1104 18992 54372 19014
rect 36078 18640 36084 18692
rect 36136 18680 36142 18692
rect 53377 18683 53435 18689
rect 53377 18680 53389 18683
rect 36136 18652 53389 18680
rect 36136 18640 36142 18652
rect 53377 18649 53389 18652
rect 53423 18649 53435 18683
rect 53558 18680 53564 18692
rect 53519 18652 53564 18680
rect 53377 18643 53435 18649
rect 53558 18640 53564 18652
rect 53616 18640 53622 18692
rect 52917 18615 52975 18621
rect 52917 18581 52929 18615
rect 52963 18612 52975 18615
rect 53576 18612 53604 18640
rect 52963 18584 53604 18612
rect 52963 18581 52975 18584
rect 52917 18575 52975 18581
rect 1104 18522 54372 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 54372 18522
rect 1104 18448 54372 18470
rect 1578 18232 1584 18284
rect 1636 18272 1642 18284
rect 1857 18275 1915 18281
rect 1857 18272 1869 18275
rect 1636 18244 1869 18272
rect 1636 18232 1642 18244
rect 1857 18241 1869 18244
rect 1903 18241 1915 18275
rect 1857 18235 1915 18241
rect 2133 18071 2191 18077
rect 2133 18037 2145 18071
rect 2179 18068 2191 18071
rect 33134 18068 33140 18080
rect 2179 18040 33140 18068
rect 2179 18037 2191 18040
rect 2133 18031 2191 18037
rect 33134 18028 33140 18040
rect 33192 18028 33198 18080
rect 1104 17978 54372 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 54372 17978
rect 1104 17904 54372 17926
rect 1578 17796 1584 17808
rect 1539 17768 1584 17796
rect 1578 17756 1584 17768
rect 1636 17756 1642 17808
rect 1104 17434 54372 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 54372 17434
rect 1104 17360 54372 17382
rect 1104 16890 54372 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 54372 16890
rect 1104 16816 54372 16838
rect 30282 16600 30288 16652
rect 30340 16640 30346 16652
rect 52825 16643 52883 16649
rect 52825 16640 52837 16643
rect 30340 16612 52837 16640
rect 30340 16600 30346 16612
rect 52825 16609 52837 16612
rect 52871 16609 52883 16643
rect 52825 16603 52883 16609
rect 52840 16572 52868 16603
rect 53377 16575 53435 16581
rect 53377 16572 53389 16575
rect 52840 16544 53389 16572
rect 53377 16541 53389 16544
rect 53423 16541 53435 16575
rect 53377 16535 53435 16541
rect 53558 16436 53564 16448
rect 53519 16408 53564 16436
rect 53558 16396 53564 16408
rect 53616 16396 53622 16448
rect 1104 16346 54372 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 54372 16346
rect 1104 16272 54372 16294
rect 1394 16096 1400 16108
rect 1355 16068 1400 16096
rect 1394 16056 1400 16068
rect 1452 16056 1458 16108
rect 1581 15895 1639 15901
rect 1581 15861 1593 15895
rect 1627 15892 1639 15895
rect 34514 15892 34520 15904
rect 1627 15864 34520 15892
rect 1627 15861 1639 15864
rect 1581 15855 1639 15861
rect 34514 15852 34520 15864
rect 34572 15852 34578 15904
rect 1104 15802 54372 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 54372 15802
rect 1104 15728 54372 15750
rect 1394 15688 1400 15700
rect 1355 15660 1400 15688
rect 1394 15648 1400 15660
rect 1452 15648 1458 15700
rect 1104 15258 54372 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 54372 15258
rect 1104 15184 54372 15206
rect 1104 14714 54372 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 54372 14714
rect 1104 14640 54372 14662
rect 1104 14170 54372 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 54372 14170
rect 1104 14096 54372 14118
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13920 1731 13923
rect 2225 13923 2283 13929
rect 2225 13920 2237 13923
rect 1719 13892 2237 13920
rect 1719 13889 1731 13892
rect 1673 13883 1731 13889
rect 2225 13889 2237 13892
rect 2271 13920 2283 13923
rect 21082 13920 21088 13932
rect 2271 13892 21088 13920
rect 2271 13889 2283 13892
rect 2225 13883 2283 13889
rect 21082 13880 21088 13892
rect 21140 13880 21146 13932
rect 52917 13923 52975 13929
rect 52917 13889 52929 13923
rect 52963 13920 52975 13923
rect 53650 13920 53656 13932
rect 52963 13892 53656 13920
rect 52963 13889 52975 13892
rect 52917 13883 52975 13889
rect 53650 13880 53656 13892
rect 53708 13880 53714 13932
rect 42058 13812 42064 13864
rect 42116 13852 42122 13864
rect 42116 13824 53512 13852
rect 42116 13812 42122 13824
rect 53484 13793 53512 13824
rect 53469 13787 53527 13793
rect 53469 13753 53481 13787
rect 53515 13753 53527 13787
rect 53469 13747 53527 13753
rect 1486 13716 1492 13728
rect 1447 13688 1492 13716
rect 1486 13676 1492 13688
rect 1544 13676 1550 13728
rect 1104 13626 54372 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 54372 13626
rect 1104 13552 54372 13574
rect 1104 13082 54372 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 54372 13082
rect 1104 13008 54372 13030
rect 1104 12538 54372 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 54372 12538
rect 1104 12464 54372 12486
rect 1104 11994 54372 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 54372 11994
rect 1104 11920 54372 11942
rect 53377 11747 53435 11753
rect 53377 11744 53389 11747
rect 52840 11716 53389 11744
rect 27430 11568 27436 11620
rect 27488 11608 27494 11620
rect 52840 11617 52868 11716
rect 53377 11713 53389 11716
rect 53423 11713 53435 11747
rect 53377 11707 53435 11713
rect 52825 11611 52883 11617
rect 52825 11608 52837 11611
rect 27488 11580 52837 11608
rect 27488 11568 27494 11580
rect 52825 11577 52837 11580
rect 52871 11577 52883 11611
rect 53558 11608 53564 11620
rect 53519 11580 53564 11608
rect 52825 11571 52883 11577
rect 53558 11568 53564 11580
rect 53616 11568 53622 11620
rect 1104 11450 54372 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 54372 11450
rect 1104 11376 54372 11398
rect 1578 11024 1584 11076
rect 1636 11064 1642 11076
rect 1857 11067 1915 11073
rect 1857 11064 1869 11067
rect 1636 11036 1869 11064
rect 1636 11024 1642 11036
rect 1857 11033 1869 11036
rect 1903 11033 1915 11067
rect 1857 11027 1915 11033
rect 2225 11067 2283 11073
rect 2225 11033 2237 11067
rect 2271 11064 2283 11067
rect 33962 11064 33968 11076
rect 2271 11036 33968 11064
rect 2271 11033 2283 11036
rect 2225 11027 2283 11033
rect 33962 11024 33968 11036
rect 34020 11024 34026 11076
rect 1104 10906 54372 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 54372 10906
rect 1104 10832 54372 10854
rect 1578 10792 1584 10804
rect 1539 10764 1584 10792
rect 1578 10752 1584 10764
rect 1636 10752 1642 10804
rect 1104 10362 54372 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 54372 10362
rect 1104 10288 54372 10310
rect 53377 9979 53435 9985
rect 53377 9976 53389 9979
rect 45526 9948 53389 9976
rect 40402 9868 40408 9920
rect 40460 9908 40466 9920
rect 45526 9908 45554 9948
rect 53377 9945 53389 9948
rect 53423 9945 53435 9979
rect 53558 9976 53564 9988
rect 53519 9948 53564 9976
rect 53377 9939 53435 9945
rect 53558 9936 53564 9948
rect 53616 9936 53622 9988
rect 40460 9880 45554 9908
rect 52917 9911 52975 9917
rect 40460 9868 40466 9880
rect 52917 9877 52929 9911
rect 52963 9908 52975 9911
rect 53576 9908 53604 9936
rect 52963 9880 53604 9908
rect 52963 9877 52975 9880
rect 52917 9871 52975 9877
rect 1104 9818 54372 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 54372 9818
rect 1104 9744 54372 9766
rect 1104 9274 54372 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 54372 9274
rect 1104 9200 54372 9222
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8925 1731 8959
rect 1673 8919 1731 8925
rect 1688 8888 1716 8919
rect 2225 8891 2283 8897
rect 2225 8888 2237 8891
rect 1688 8860 2237 8888
rect 2225 8857 2237 8860
rect 2271 8888 2283 8891
rect 29454 8888 29460 8900
rect 2271 8860 29460 8888
rect 2271 8857 2283 8860
rect 2225 8851 2283 8857
rect 29454 8848 29460 8860
rect 29512 8848 29518 8900
rect 1486 8820 1492 8832
rect 1447 8792 1492 8820
rect 1486 8780 1492 8792
rect 1544 8780 1550 8832
rect 1104 8730 54372 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 54372 8730
rect 1104 8656 54372 8678
rect 1104 8186 54372 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 54372 8186
rect 1104 8112 54372 8134
rect 1104 7642 54372 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 54372 7642
rect 1104 7568 54372 7590
rect 1854 7392 1860 7404
rect 1815 7364 1860 7392
rect 1854 7352 1860 7364
rect 1912 7352 1918 7404
rect 52917 7395 52975 7401
rect 52917 7361 52929 7395
rect 52963 7392 52975 7395
rect 53650 7392 53656 7404
rect 52963 7364 53656 7392
rect 52963 7361 52975 7364
rect 52917 7355 52975 7361
rect 53650 7352 53656 7364
rect 53708 7352 53714 7404
rect 53469 7259 53527 7265
rect 53469 7256 53481 7259
rect 45526 7228 53481 7256
rect 1949 7191 2007 7197
rect 1949 7157 1961 7191
rect 1995 7188 2007 7191
rect 13630 7188 13636 7200
rect 1995 7160 13636 7188
rect 1995 7157 2007 7160
rect 1949 7151 2007 7157
rect 13630 7148 13636 7160
rect 13688 7148 13694 7200
rect 17954 7148 17960 7200
rect 18012 7188 18018 7200
rect 45526 7188 45554 7228
rect 53469 7225 53481 7228
rect 53515 7225 53527 7259
rect 53469 7219 53527 7225
rect 18012 7160 45554 7188
rect 18012 7148 18018 7160
rect 1104 7098 54372 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 54372 7098
rect 1104 7024 54372 7046
rect 1578 6944 1584 6996
rect 1636 6984 1642 6996
rect 1673 6987 1731 6993
rect 1673 6984 1685 6987
rect 1636 6956 1685 6984
rect 1636 6944 1642 6956
rect 1673 6953 1685 6956
rect 1719 6984 1731 6987
rect 1854 6984 1860 6996
rect 1719 6956 1860 6984
rect 1719 6953 1731 6956
rect 1673 6947 1731 6953
rect 1854 6944 1860 6956
rect 1912 6944 1918 6996
rect 1104 6554 54372 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 54372 6554
rect 1104 6480 54372 6502
rect 1104 6010 54372 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 54372 6010
rect 1104 5936 54372 5958
rect 1104 5466 54372 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 54372 5466
rect 1104 5392 54372 5414
rect 53377 5219 53435 5225
rect 53377 5216 53389 5219
rect 52840 5188 53389 5216
rect 38102 5040 38108 5092
rect 38160 5080 38166 5092
rect 52840 5089 52868 5188
rect 53377 5185 53389 5188
rect 53423 5185 53435 5219
rect 53377 5179 53435 5185
rect 52825 5083 52883 5089
rect 52825 5080 52837 5083
rect 38160 5052 52837 5080
rect 38160 5040 38166 5052
rect 52825 5049 52837 5052
rect 52871 5049 52883 5083
rect 52825 5043 52883 5049
rect 53558 5012 53564 5024
rect 53519 4984 53564 5012
rect 53558 4972 53564 4984
rect 53616 4972 53622 5024
rect 1104 4922 54372 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 54372 4922
rect 1104 4848 54372 4870
rect 1673 4607 1731 4613
rect 1673 4573 1685 4607
rect 1719 4604 1731 4607
rect 2225 4607 2283 4613
rect 2225 4604 2237 4607
rect 1719 4576 2237 4604
rect 1719 4573 1731 4576
rect 1673 4567 1731 4573
rect 2225 4573 2237 4576
rect 2271 4604 2283 4607
rect 15930 4604 15936 4616
rect 2271 4576 15936 4604
rect 2271 4573 2283 4576
rect 2225 4567 2283 4573
rect 15930 4564 15936 4576
rect 15988 4564 15994 4616
rect 1486 4468 1492 4480
rect 1447 4440 1492 4468
rect 1486 4428 1492 4440
rect 1544 4428 1550 4480
rect 1104 4378 54372 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 54372 4378
rect 1104 4304 54372 4326
rect 1104 3834 54372 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 54372 3834
rect 1104 3760 54372 3782
rect 53377 3519 53435 3525
rect 53377 3516 53389 3519
rect 52840 3488 53389 3516
rect 33502 3408 33508 3460
rect 33560 3448 33566 3460
rect 52840 3457 52868 3488
rect 53377 3485 53389 3488
rect 53423 3485 53435 3519
rect 53377 3479 53435 3485
rect 52825 3451 52883 3457
rect 52825 3448 52837 3451
rect 33560 3420 52837 3448
rect 33560 3408 33566 3420
rect 52825 3417 52837 3420
rect 52871 3417 52883 3451
rect 52825 3411 52883 3417
rect 1302 3340 1308 3392
rect 1360 3380 1366 3392
rect 1581 3383 1639 3389
rect 1581 3380 1593 3383
rect 1360 3352 1593 3380
rect 1360 3340 1366 3352
rect 1581 3349 1593 3352
rect 1627 3349 1639 3383
rect 1581 3343 1639 3349
rect 1854 3340 1860 3392
rect 1912 3380 1918 3392
rect 2133 3383 2191 3389
rect 2133 3380 2145 3383
rect 1912 3352 2145 3380
rect 1912 3340 1918 3352
rect 2133 3349 2145 3352
rect 2179 3349 2191 3383
rect 2133 3343 2191 3349
rect 53561 3383 53619 3389
rect 53561 3349 53573 3383
rect 53607 3380 53619 3383
rect 54110 3380 54116 3392
rect 53607 3352 54116 3380
rect 53607 3349 53619 3352
rect 53561 3343 53619 3349
rect 54110 3340 54116 3352
rect 54168 3340 54174 3392
rect 1104 3290 54372 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 54372 3290
rect 1104 3216 54372 3238
rect 51442 3176 51448 3188
rect 51403 3148 51448 3176
rect 51442 3136 51448 3148
rect 51500 3136 51506 3188
rect 14 3000 20 3052
rect 72 3040 78 3052
rect 1302 3040 1308 3052
rect 72 3012 1308 3040
rect 72 3000 78 3012
rect 1302 3000 1308 3012
rect 1360 3040 1366 3052
rect 1857 3043 1915 3049
rect 1857 3040 1869 3043
rect 1360 3012 1869 3040
rect 1360 3000 1366 3012
rect 1857 3009 1869 3012
rect 1903 3009 1915 3043
rect 53377 3043 53435 3049
rect 53377 3040 53389 3043
rect 1857 3003 1915 3009
rect 52840 3012 53389 3040
rect 2133 2975 2191 2981
rect 2133 2941 2145 2975
rect 2179 2972 2191 2975
rect 34422 2972 34428 2984
rect 2179 2944 34428 2972
rect 2179 2941 2191 2944
rect 2133 2935 2191 2941
rect 34422 2932 34428 2944
rect 34480 2932 34486 2984
rect 13262 2864 13268 2916
rect 13320 2904 13326 2916
rect 13449 2907 13507 2913
rect 13449 2904 13461 2907
rect 13320 2876 13461 2904
rect 13320 2864 13326 2876
rect 13449 2873 13461 2876
rect 13495 2904 13507 2907
rect 30558 2904 30564 2916
rect 13495 2876 30564 2904
rect 13495 2873 13507 2876
rect 13449 2867 13507 2873
rect 30558 2864 30564 2876
rect 30616 2864 30622 2916
rect 31110 2864 31116 2916
rect 31168 2904 31174 2916
rect 52840 2913 52868 3012
rect 53377 3009 53389 3012
rect 53423 3009 53435 3043
rect 53377 3003 53435 3009
rect 52825 2907 52883 2913
rect 52825 2904 52837 2907
rect 31168 2876 52837 2904
rect 31168 2864 31174 2876
rect 52825 2873 52837 2876
rect 52871 2873 52883 2907
rect 52825 2867 52883 2873
rect 1946 2796 1952 2848
rect 2004 2836 2010 2848
rect 2774 2836 2780 2848
rect 2004 2808 2780 2836
rect 2004 2796 2010 2808
rect 2774 2796 2780 2808
rect 2832 2796 2838 2848
rect 6454 2836 6460 2848
rect 6415 2808 6460 2836
rect 6454 2796 6460 2808
rect 6512 2796 6518 2848
rect 19334 2836 19340 2848
rect 19295 2808 19340 2836
rect 19334 2796 19340 2808
rect 19392 2796 19398 2848
rect 21266 2796 21272 2848
rect 21324 2836 21330 2848
rect 22097 2839 22155 2845
rect 22097 2836 22109 2839
rect 21324 2808 22109 2836
rect 21324 2796 21330 2808
rect 22097 2805 22109 2808
rect 22143 2836 22155 2839
rect 22278 2836 22284 2848
rect 22143 2808 22284 2836
rect 22143 2805 22155 2808
rect 22097 2799 22155 2805
rect 22278 2796 22284 2808
rect 22336 2796 22342 2848
rect 32214 2836 32220 2848
rect 32175 2808 32220 2836
rect 32214 2796 32220 2808
rect 32272 2796 32278 2848
rect 34514 2796 34520 2848
rect 34572 2836 34578 2848
rect 34885 2839 34943 2845
rect 34885 2836 34897 2839
rect 34572 2808 34897 2836
rect 34572 2796 34578 2808
rect 34885 2805 34897 2808
rect 34931 2805 34943 2839
rect 45094 2836 45100 2848
rect 45055 2808 45100 2836
rect 34885 2799 34943 2805
rect 45094 2796 45100 2808
rect 45152 2796 45158 2848
rect 47670 2796 47676 2848
rect 47728 2836 47734 2848
rect 47765 2839 47823 2845
rect 47765 2836 47777 2839
rect 47728 2808 47777 2836
rect 47728 2796 47734 2808
rect 47765 2805 47777 2808
rect 47811 2805 47823 2839
rect 50338 2836 50344 2848
rect 50299 2808 50344 2836
rect 47765 2799 47823 2805
rect 50338 2796 50344 2808
rect 50396 2796 50402 2848
rect 52181 2839 52239 2845
rect 52181 2805 52193 2839
rect 52227 2836 52239 2839
rect 52454 2836 52460 2848
rect 52227 2808 52460 2836
rect 52227 2805 52239 2808
rect 52181 2799 52239 2805
rect 52454 2796 52460 2808
rect 52512 2796 52518 2848
rect 53558 2836 53564 2848
rect 53519 2808 53564 2836
rect 53558 2796 53564 2808
rect 53616 2796 53622 2848
rect 1104 2746 54372 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 54372 2746
rect 1104 2672 54372 2694
rect 2133 2635 2191 2641
rect 2133 2601 2145 2635
rect 2179 2632 2191 2635
rect 21542 2632 21548 2644
rect 2179 2604 21548 2632
rect 2179 2601 2191 2604
rect 2133 2595 2191 2601
rect 21542 2592 21548 2604
rect 21600 2592 21606 2644
rect 22186 2592 22192 2644
rect 22244 2632 22250 2644
rect 22373 2635 22431 2641
rect 22373 2632 22385 2635
rect 22244 2604 22385 2632
rect 22244 2592 22250 2604
rect 22373 2601 22385 2604
rect 22419 2601 22431 2635
rect 25961 2635 26019 2641
rect 25961 2632 25973 2635
rect 22373 2595 22431 2601
rect 22480 2604 25973 2632
rect 6733 2567 6791 2573
rect 6733 2533 6745 2567
rect 6779 2564 6791 2567
rect 14274 2564 14280 2576
rect 6779 2536 14280 2564
rect 6779 2533 6791 2536
rect 6733 2527 6791 2533
rect 14274 2524 14280 2536
rect 14332 2524 14338 2576
rect 15010 2524 15016 2576
rect 15068 2564 15074 2576
rect 15105 2567 15163 2573
rect 15105 2564 15117 2567
rect 15068 2536 15117 2564
rect 15068 2524 15074 2536
rect 15105 2533 15117 2536
rect 15151 2533 15163 2567
rect 19426 2564 19432 2576
rect 15105 2527 15163 2533
rect 16546 2536 19432 2564
rect 2961 2499 3019 2505
rect 2961 2465 2973 2499
rect 3007 2496 3019 2499
rect 3007 2468 10272 2496
rect 3007 2465 3019 2468
rect 2961 2459 3019 2465
rect 2774 2428 2780 2440
rect 2735 2400 2780 2428
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2428 4307 2431
rect 4295 2400 4844 2428
rect 4295 2397 4307 2400
rect 4249 2391 4307 2397
rect 1854 2360 1860 2372
rect 1815 2332 1860 2360
rect 1854 2320 1860 2332
rect 1912 2320 1918 2372
rect 4816 2304 4844 2400
rect 6454 2388 6460 2440
rect 6512 2428 6518 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 6512 2400 6561 2428
rect 6512 2388 6518 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 8941 2431 8999 2437
rect 8941 2428 8953 2431
rect 6549 2391 6607 2397
rect 8404 2400 8953 2428
rect 8404 2304 8432 2400
rect 8941 2397 8953 2400
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 10244 2360 10272 2468
rect 10318 2456 10324 2508
rect 10376 2496 10382 2508
rect 10965 2499 11023 2505
rect 10965 2496 10977 2499
rect 10376 2468 10977 2496
rect 10376 2456 10382 2468
rect 10965 2465 10977 2468
rect 11011 2496 11023 2499
rect 11517 2499 11575 2505
rect 11517 2496 11529 2499
rect 11011 2468 11529 2496
rect 11011 2465 11023 2468
rect 10965 2459 11023 2465
rect 11517 2465 11529 2468
rect 11563 2465 11575 2499
rect 16546 2496 16574 2536
rect 19426 2524 19432 2536
rect 19484 2524 19490 2576
rect 22480 2564 22508 2604
rect 25961 2601 25973 2604
rect 26007 2601 26019 2635
rect 25961 2595 26019 2601
rect 28166 2592 28172 2644
rect 28224 2632 28230 2644
rect 50706 2632 50712 2644
rect 28224 2604 45554 2632
rect 50667 2604 50712 2632
rect 28224 2592 28230 2604
rect 24578 2564 24584 2576
rect 19628 2536 22508 2564
rect 24539 2536 24584 2564
rect 11517 2459 11575 2465
rect 13188 2468 16574 2496
rect 10689 2431 10747 2437
rect 10689 2397 10701 2431
rect 10735 2428 10747 2431
rect 13188 2428 13216 2468
rect 16850 2456 16856 2508
rect 16908 2496 16914 2508
rect 19628 2496 19656 2536
rect 24578 2524 24584 2536
rect 24636 2524 24642 2576
rect 32493 2567 32551 2573
rect 32493 2564 32505 2567
rect 26206 2536 32505 2564
rect 16908 2468 19656 2496
rect 19705 2499 19763 2505
rect 16908 2456 16914 2468
rect 19705 2465 19717 2499
rect 19751 2496 19763 2499
rect 19978 2496 19984 2508
rect 19751 2468 19984 2496
rect 19751 2465 19763 2468
rect 19705 2459 19763 2465
rect 19978 2456 19984 2468
rect 20036 2456 20042 2508
rect 23750 2456 23756 2508
rect 23808 2496 23814 2508
rect 26206 2496 26234 2536
rect 32493 2533 32505 2536
rect 32539 2533 32551 2567
rect 32493 2527 32551 2533
rect 35345 2567 35403 2573
rect 35345 2533 35357 2567
rect 35391 2564 35403 2567
rect 35894 2564 35900 2576
rect 35391 2536 35900 2564
rect 35391 2533 35403 2536
rect 35345 2527 35403 2533
rect 35894 2524 35900 2536
rect 35952 2524 35958 2576
rect 36906 2524 36912 2576
rect 36964 2564 36970 2576
rect 38933 2567 38991 2573
rect 38933 2564 38945 2567
rect 36964 2536 38945 2564
rect 36964 2524 36970 2536
rect 38933 2533 38945 2536
rect 38979 2533 38991 2567
rect 38933 2527 38991 2533
rect 41506 2524 41512 2576
rect 41564 2564 41570 2576
rect 41601 2567 41659 2573
rect 41601 2564 41613 2567
rect 41564 2536 41613 2564
rect 41564 2524 41570 2536
rect 41601 2533 41613 2536
rect 41647 2533 41659 2567
rect 45526 2564 45554 2604
rect 50706 2592 50712 2604
rect 50764 2592 50770 2644
rect 53285 2567 53343 2573
rect 53285 2564 53297 2567
rect 45526 2536 53297 2564
rect 41601 2527 41659 2533
rect 53285 2533 53297 2536
rect 53331 2533 53343 2567
rect 53285 2527 53343 2533
rect 30650 2496 30656 2508
rect 23808 2468 26234 2496
rect 30611 2468 30656 2496
rect 23808 2456 23814 2468
rect 30650 2456 30656 2468
rect 30708 2456 30714 2508
rect 10735 2400 13216 2428
rect 10735 2397 10747 2400
rect 10689 2391 10747 2397
rect 13262 2388 13268 2440
rect 13320 2428 13326 2440
rect 14461 2431 14519 2437
rect 13320 2400 13365 2428
rect 13320 2388 13326 2400
rect 14461 2397 14473 2431
rect 14507 2428 14519 2431
rect 14826 2428 14832 2440
rect 14507 2400 14832 2428
rect 14507 2397 14519 2400
rect 14461 2391 14519 2397
rect 14826 2388 14832 2400
rect 14884 2428 14890 2440
rect 14921 2431 14979 2437
rect 14921 2428 14933 2431
rect 14884 2400 14933 2428
rect 14884 2388 14890 2400
rect 14921 2397 14933 2400
rect 14967 2397 14979 2431
rect 14921 2391 14979 2397
rect 17129 2431 17187 2437
rect 17129 2397 17141 2431
rect 17175 2428 17187 2431
rect 17175 2400 17724 2428
rect 17175 2397 17187 2400
rect 17129 2391 17187 2397
rect 16298 2360 16304 2372
rect 10244 2332 16304 2360
rect 16298 2320 16304 2332
rect 16356 2320 16362 2372
rect 17696 2304 17724 2400
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 19392 2400 19441 2428
rect 19392 2388 19398 2400
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 22278 2428 22284 2440
rect 22239 2400 22284 2428
rect 19429 2391 19487 2397
rect 22278 2388 22284 2400
rect 22336 2388 22342 2440
rect 24397 2431 24455 2437
rect 24397 2428 24409 2431
rect 23860 2400 24409 2428
rect 23860 2304 23888 2400
rect 24397 2397 24409 2400
rect 24443 2397 24455 2431
rect 24397 2391 24455 2397
rect 29917 2431 29975 2437
rect 29917 2397 29929 2431
rect 29963 2428 29975 2431
rect 30282 2428 30288 2440
rect 29963 2400 30288 2428
rect 29963 2397 29975 2400
rect 29917 2391 29975 2397
rect 30282 2388 30288 2400
rect 30340 2428 30346 2440
rect 30377 2431 30435 2437
rect 30377 2428 30389 2431
rect 30340 2400 30389 2428
rect 30340 2388 30346 2400
rect 30377 2397 30389 2400
rect 30423 2397 30435 2431
rect 30377 2391 30435 2397
rect 32214 2388 32220 2440
rect 32272 2428 32278 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 32272 2400 32321 2428
rect 32272 2388 32278 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 35342 2428 35348 2440
rect 32309 2391 32367 2397
rect 32416 2400 35348 2428
rect 25409 2363 25467 2369
rect 25409 2329 25421 2363
rect 25455 2360 25467 2363
rect 25774 2360 25780 2372
rect 25455 2332 25780 2360
rect 25455 2329 25467 2332
rect 25409 2323 25467 2329
rect 25774 2320 25780 2332
rect 25832 2360 25838 2372
rect 26053 2363 26111 2369
rect 26053 2360 26065 2363
rect 25832 2332 26065 2360
rect 25832 2320 25838 2332
rect 26053 2329 26065 2332
rect 26099 2329 26111 2363
rect 26053 2323 26111 2329
rect 27341 2363 27399 2369
rect 27341 2329 27353 2363
rect 27387 2360 27399 2363
rect 27706 2360 27712 2372
rect 27387 2332 27712 2360
rect 27387 2329 27399 2332
rect 27341 2323 27399 2329
rect 27706 2320 27712 2332
rect 27764 2360 27770 2372
rect 27893 2363 27951 2369
rect 27893 2360 27905 2363
rect 27764 2332 27905 2360
rect 27764 2320 27770 2332
rect 27893 2329 27905 2332
rect 27939 2329 27951 2363
rect 27893 2323 27951 2329
rect 28077 2363 28135 2369
rect 28077 2329 28089 2363
rect 28123 2360 28135 2363
rect 32416 2360 32444 2400
rect 35342 2388 35348 2400
rect 35400 2388 35406 2440
rect 36725 2431 36783 2437
rect 36725 2397 36737 2431
rect 36771 2428 36783 2431
rect 37553 2431 37611 2437
rect 37553 2428 37565 2431
rect 36771 2400 37565 2428
rect 36771 2397 36783 2400
rect 36725 2391 36783 2397
rect 37553 2397 37565 2400
rect 37599 2428 37611 2431
rect 37734 2428 37740 2440
rect 37599 2400 37740 2428
rect 37599 2397 37611 2400
rect 37553 2391 37611 2397
rect 37734 2388 37740 2400
rect 37792 2388 37798 2440
rect 38289 2431 38347 2437
rect 38289 2397 38301 2431
rect 38335 2428 38347 2431
rect 38654 2428 38660 2440
rect 38335 2400 38660 2428
rect 38335 2397 38347 2400
rect 38289 2391 38347 2397
rect 38654 2388 38660 2400
rect 38712 2428 38718 2440
rect 38749 2431 38807 2437
rect 38749 2428 38761 2431
rect 38712 2400 38761 2428
rect 38712 2388 38718 2400
rect 38749 2397 38761 2400
rect 38795 2397 38807 2431
rect 43257 2431 43315 2437
rect 43257 2428 43269 2431
rect 38749 2391 38807 2397
rect 42812 2400 43269 2428
rect 28123 2332 32444 2360
rect 28123 2329 28135 2332
rect 28077 2323 28135 2329
rect 34514 2320 34520 2372
rect 34572 2360 34578 2372
rect 35161 2363 35219 2369
rect 35161 2360 35173 2363
rect 34572 2332 35173 2360
rect 34572 2320 34578 2332
rect 35161 2329 35173 2332
rect 35207 2329 35219 2363
rect 35161 2323 35219 2329
rect 40865 2363 40923 2369
rect 40865 2329 40877 2363
rect 40911 2360 40923 2363
rect 41230 2360 41236 2372
rect 40911 2332 41236 2360
rect 40911 2329 40923 2332
rect 40865 2323 40923 2329
rect 41230 2320 41236 2332
rect 41288 2360 41294 2372
rect 41417 2363 41475 2369
rect 41417 2360 41429 2363
rect 41288 2332 41429 2360
rect 41288 2320 41294 2332
rect 41417 2329 41429 2332
rect 41463 2329 41475 2363
rect 41417 2323 41475 2329
rect 42812 2304 42840 2400
rect 43257 2397 43269 2400
rect 43303 2397 43315 2431
rect 43257 2391 43315 2397
rect 45094 2388 45100 2440
rect 45152 2428 45158 2440
rect 45189 2431 45247 2437
rect 45189 2428 45201 2431
rect 45152 2400 45201 2428
rect 45152 2388 45158 2400
rect 45189 2397 45201 2400
rect 45235 2397 45247 2431
rect 45189 2391 45247 2397
rect 49694 2388 49700 2440
rect 49752 2428 49758 2440
rect 50338 2428 50344 2440
rect 49752 2400 50344 2428
rect 49752 2388 49758 2400
rect 50338 2388 50344 2400
rect 50396 2428 50402 2440
rect 50617 2431 50675 2437
rect 50617 2428 50629 2431
rect 50396 2400 50629 2428
rect 50396 2388 50402 2400
rect 50617 2397 50629 2400
rect 50663 2397 50675 2431
rect 50617 2391 50675 2397
rect 51442 2388 51448 2440
rect 51500 2428 51506 2440
rect 51629 2431 51687 2437
rect 51629 2428 51641 2431
rect 51500 2400 51641 2428
rect 51500 2388 51506 2400
rect 51629 2397 51641 2400
rect 51675 2397 51687 2431
rect 51629 2391 51687 2397
rect 47670 2320 47676 2372
rect 47728 2360 47734 2372
rect 48041 2363 48099 2369
rect 48041 2360 48053 2363
rect 47728 2332 48053 2360
rect 47728 2320 47734 2332
rect 48041 2329 48053 2332
rect 48087 2329 48099 2363
rect 48041 2323 48099 2329
rect 52454 2320 52460 2372
rect 52512 2360 52518 2372
rect 53558 2360 53564 2372
rect 52512 2332 53564 2360
rect 52512 2320 52518 2332
rect 53558 2320 53564 2332
rect 53616 2320 53622 2372
rect 3878 2252 3884 2304
rect 3936 2292 3942 2304
rect 4065 2295 4123 2301
rect 4065 2292 4077 2295
rect 3936 2264 4077 2292
rect 3936 2252 3942 2264
rect 4065 2261 4077 2264
rect 4111 2261 4123 2295
rect 4798 2292 4804 2304
rect 4759 2264 4804 2292
rect 4065 2255 4123 2261
rect 4798 2252 4804 2264
rect 4856 2252 4862 2304
rect 8386 2292 8392 2304
rect 8347 2264 8392 2292
rect 8386 2252 8392 2264
rect 8444 2252 8450 2304
rect 9122 2292 9128 2304
rect 9083 2264 9128 2292
rect 9122 2252 9128 2264
rect 9180 2252 9186 2304
rect 12894 2252 12900 2304
rect 12952 2292 12958 2304
rect 13081 2295 13139 2301
rect 13081 2292 13093 2295
rect 12952 2264 13093 2292
rect 12952 2252 12958 2264
rect 13081 2261 13093 2264
rect 13127 2261 13139 2295
rect 13081 2255 13139 2261
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 16945 2295 17003 2301
rect 16945 2292 16957 2295
rect 16816 2264 16957 2292
rect 16816 2252 16822 2264
rect 16945 2261 16957 2264
rect 16991 2261 17003 2295
rect 17678 2292 17684 2304
rect 17639 2264 17684 2292
rect 16945 2255 17003 2261
rect 17678 2252 17684 2264
rect 17736 2252 17742 2304
rect 23842 2292 23848 2304
rect 23803 2264 23848 2292
rect 23842 2252 23848 2264
rect 23900 2252 23906 2304
rect 36722 2252 36728 2304
rect 36780 2292 36786 2304
rect 37369 2295 37427 2301
rect 37369 2292 37381 2295
rect 36780 2264 37381 2292
rect 36780 2252 36786 2264
rect 37369 2261 37381 2264
rect 37415 2261 37427 2295
rect 42794 2292 42800 2304
rect 42755 2264 42800 2292
rect 37369 2255 37427 2261
rect 42794 2252 42800 2264
rect 42852 2252 42858 2304
rect 43162 2252 43168 2304
rect 43220 2292 43226 2304
rect 43441 2295 43499 2301
rect 43441 2292 43453 2295
rect 43220 2264 43453 2292
rect 43220 2252 43226 2264
rect 43441 2261 43453 2264
rect 43487 2261 43499 2295
rect 45370 2292 45376 2304
rect 45331 2264 45376 2292
rect 43441 2255 43499 2261
rect 45370 2252 45376 2264
rect 45428 2252 45434 2304
rect 48130 2292 48136 2304
rect 48091 2264 48136 2292
rect 48130 2252 48136 2264
rect 48188 2252 48194 2304
rect 51534 2252 51540 2304
rect 51592 2292 51598 2304
rect 51813 2295 51871 2301
rect 51813 2292 51825 2295
rect 51592 2264 51825 2292
rect 51592 2252 51598 2264
rect 51813 2261 51825 2264
rect 51859 2261 51871 2295
rect 51813 2255 51871 2261
rect 1104 2202 54372 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 54372 2202
rect 1104 2128 54372 2150
rect 4798 1980 4804 2032
rect 4856 2020 4862 2032
rect 22462 2020 22468 2032
rect 4856 1992 22468 2020
rect 4856 1980 4862 1992
rect 22462 1980 22468 1992
rect 22520 1980 22526 2032
rect 28350 1980 28356 2032
rect 28408 2020 28414 2032
rect 42794 2020 42800 2032
rect 28408 1992 42800 2020
rect 28408 1980 28414 1992
rect 42794 1980 42800 1992
rect 42852 1980 42858 2032
rect 17678 1912 17684 1964
rect 17736 1952 17742 1964
rect 26786 1952 26792 1964
rect 17736 1924 26792 1952
rect 17736 1912 17742 1924
rect 26786 1912 26792 1924
rect 26844 1912 26850 1964
rect 24946 1844 24952 1896
rect 25004 1884 25010 1896
rect 48130 1884 48136 1896
rect 25004 1856 48136 1884
rect 25004 1844 25010 1856
rect 48130 1844 48136 1856
rect 48188 1844 48194 1896
<< via1 >>
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 5816 54816 5868 54868
rect 14188 54816 14240 54868
rect 24676 54816 24728 54868
rect 25136 54816 25188 54868
rect 29644 54816 29696 54868
rect 36084 54816 36136 54868
rect 38660 54816 38712 54868
rect 40592 54816 40644 54868
rect 47032 54816 47084 54868
rect 48964 54816 49016 54868
rect 51540 54816 51592 54868
rect 3884 54680 3936 54732
rect 1400 54655 1452 54664
rect 1400 54621 1409 54655
rect 1409 54621 1443 54655
rect 1443 54621 1452 54655
rect 1400 54612 1452 54621
rect 1676 54655 1728 54664
rect 1676 54621 1685 54655
rect 1685 54621 1719 54655
rect 1719 54621 1728 54655
rect 1676 54612 1728 54621
rect 6644 54655 6696 54664
rect 2780 54587 2832 54596
rect 2780 54553 2789 54587
rect 2789 54553 2823 54587
rect 2823 54553 2832 54587
rect 2780 54544 2832 54553
rect 6644 54621 6653 54655
rect 6653 54621 6687 54655
rect 6687 54621 6696 54655
rect 14648 54748 14700 54800
rect 22192 54748 22244 54800
rect 22376 54748 22428 54800
rect 10324 54680 10376 54732
rect 10968 54723 11020 54732
rect 10968 54689 10977 54723
rect 10977 54689 11011 54723
rect 11011 54689 11020 54723
rect 10968 54680 11020 54689
rect 27712 54680 27764 54732
rect 6644 54612 6696 54621
rect 7748 54612 7800 54664
rect 10692 54655 10744 54664
rect 10692 54621 10701 54655
rect 10701 54621 10735 54655
rect 10735 54621 10744 54655
rect 10692 54612 10744 54621
rect 12256 54612 12308 54664
rect 14648 54544 14700 54596
rect 18696 54655 18748 54664
rect 2872 54519 2924 54528
rect 2872 54485 2881 54519
rect 2881 54485 2915 54519
rect 2915 54485 2924 54519
rect 2872 54476 2924 54485
rect 8024 54519 8076 54528
rect 8024 54485 8033 54519
rect 8033 54485 8067 54519
rect 8067 54485 8076 54519
rect 8024 54476 8076 54485
rect 15108 54519 15160 54528
rect 15108 54485 15117 54519
rect 15117 54485 15151 54519
rect 15151 54485 15160 54519
rect 15108 54476 15160 54485
rect 16764 54476 16816 54528
rect 18696 54621 18705 54655
rect 18705 54621 18739 54655
rect 18739 54621 18748 54655
rect 18696 54612 18748 54621
rect 21272 54612 21324 54664
rect 23204 54612 23256 54664
rect 22284 54587 22336 54596
rect 18880 54476 18932 54528
rect 22284 54553 22293 54587
rect 22293 54553 22327 54587
rect 22327 54553 22336 54587
rect 22284 54544 22336 54553
rect 24860 54544 24912 54596
rect 25228 54612 25280 54664
rect 27896 54612 27948 54664
rect 28172 54612 28224 54664
rect 30472 54612 30524 54664
rect 33876 54680 33928 54732
rect 45100 54680 45152 54732
rect 32680 54655 32732 54664
rect 32404 54544 32456 54596
rect 32680 54621 32689 54655
rect 32689 54621 32723 54655
rect 32723 54621 32732 54655
rect 32680 54612 32732 54621
rect 36084 54612 36136 54664
rect 38660 54612 38712 54664
rect 34520 54544 34572 54596
rect 42800 54655 42852 54664
rect 42800 54621 42809 54655
rect 42809 54621 42843 54655
rect 42843 54621 42852 54655
rect 42800 54612 42852 54621
rect 45468 54655 45520 54664
rect 45468 54621 45477 54655
rect 45477 54621 45511 54655
rect 45511 54621 45520 54655
rect 45468 54612 45520 54621
rect 47584 54655 47636 54664
rect 47584 54621 47593 54655
rect 47593 54621 47627 54655
rect 47627 54621 47636 54655
rect 47584 54612 47636 54621
rect 48964 54612 49016 54664
rect 51632 54655 51684 54664
rect 51632 54621 51641 54655
rect 51641 54621 51675 54655
rect 51675 54621 51684 54655
rect 51632 54612 51684 54621
rect 53472 54612 53524 54664
rect 24032 54476 24084 54528
rect 30104 54476 30156 54528
rect 30748 54476 30800 54528
rect 33048 54476 33100 54528
rect 34796 54476 34848 54528
rect 38844 54519 38896 54528
rect 38844 54485 38853 54519
rect 38853 54485 38887 54519
rect 38887 54485 38896 54519
rect 38844 54476 38896 54485
rect 40132 54519 40184 54528
rect 40132 54485 40141 54519
rect 40141 54485 40175 54519
rect 40175 54485 40184 54519
rect 40132 54476 40184 54485
rect 42616 54519 42668 54528
rect 42616 54485 42625 54519
rect 42625 54485 42659 54519
rect 42659 54485 42668 54519
rect 42616 54476 42668 54485
rect 49148 54519 49200 54528
rect 49148 54485 49157 54519
rect 49157 54485 49191 54519
rect 49191 54485 49200 54519
rect 49148 54476 49200 54485
rect 53656 54476 53708 54528
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 2780 54272 2832 54324
rect 3884 54315 3936 54324
rect 3884 54281 3893 54315
rect 3893 54281 3927 54315
rect 3927 54281 3936 54315
rect 3884 54272 3936 54281
rect 6644 54272 6696 54324
rect 10968 54272 11020 54324
rect 22284 54272 22336 54324
rect 23204 54315 23256 54324
rect 23204 54281 23213 54315
rect 23213 54281 23247 54315
rect 23247 54281 23256 54315
rect 23204 54272 23256 54281
rect 24676 54272 24728 54324
rect 31392 54272 31444 54324
rect 34520 54272 34572 54324
rect 1308 54204 1360 54256
rect 22192 54204 22244 54256
rect 30564 54204 30616 54256
rect 31208 54204 31260 54256
rect 40132 54272 40184 54324
rect 45100 54315 45152 54324
rect 45100 54281 45109 54315
rect 45109 54281 45143 54315
rect 45143 54281 45152 54315
rect 45100 54272 45152 54281
rect 53564 54247 53616 54256
rect 53564 54213 53573 54247
rect 53573 54213 53607 54247
rect 53607 54213 53616 54247
rect 53564 54204 53616 54213
rect 28264 54136 28316 54188
rect 15108 54068 15160 54120
rect 2136 54000 2188 54052
rect 29460 54136 29512 54188
rect 24860 53932 24912 53984
rect 25964 53932 26016 53984
rect 26976 53975 27028 53984
rect 26976 53941 26985 53975
rect 26985 53941 27019 53975
rect 27019 53941 27028 53975
rect 26976 53932 27028 53941
rect 28080 53932 28132 53984
rect 30104 54068 30156 54120
rect 31944 54068 31996 54120
rect 32404 54111 32456 54120
rect 32404 54077 32413 54111
rect 32413 54077 32447 54111
rect 32447 54077 32456 54111
rect 32404 54068 32456 54077
rect 32680 54136 32732 54188
rect 33048 54136 33100 54188
rect 33324 54136 33376 54188
rect 42616 54000 42668 54052
rect 53380 54043 53432 54052
rect 53380 54009 53389 54043
rect 53389 54009 53423 54043
rect 53423 54009 53432 54043
rect 53380 54000 53432 54009
rect 28908 53975 28960 53984
rect 28908 53941 28917 53975
rect 28917 53941 28951 53975
rect 28951 53941 28960 53975
rect 28908 53932 28960 53941
rect 29552 53932 29604 53984
rect 30748 53932 30800 53984
rect 32220 53932 32272 53984
rect 33232 53932 33284 53984
rect 33416 53975 33468 53984
rect 33416 53941 33425 53975
rect 33425 53941 33459 53975
rect 33459 53941 33468 53975
rect 33416 53932 33468 53941
rect 36084 53975 36136 53984
rect 36084 53941 36093 53975
rect 36093 53941 36127 53975
rect 36127 53941 36136 53975
rect 36084 53932 36136 53941
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 1308 53728 1360 53780
rect 29460 53592 29512 53644
rect 28080 53524 28132 53576
rect 31300 53728 31352 53780
rect 31392 53703 31444 53712
rect 31392 53669 31401 53703
rect 31401 53669 31435 53703
rect 31435 53669 31444 53703
rect 31392 53660 31444 53669
rect 33416 53728 33468 53780
rect 34428 53728 34480 53780
rect 33324 53660 33376 53712
rect 36176 53728 36228 53780
rect 30012 53635 30064 53644
rect 30012 53601 30021 53635
rect 30021 53601 30055 53635
rect 30055 53601 30064 53635
rect 30012 53592 30064 53601
rect 27160 53499 27212 53508
rect 27160 53465 27194 53499
rect 27194 53465 27212 53499
rect 30564 53567 30616 53576
rect 30564 53533 30573 53567
rect 30573 53533 30607 53567
rect 30607 53533 30616 53567
rect 30564 53524 30616 53533
rect 30748 53567 30800 53576
rect 30748 53533 30757 53567
rect 30757 53533 30791 53567
rect 30791 53533 30800 53567
rect 30748 53524 30800 53533
rect 32128 53524 32180 53576
rect 27160 53456 27212 53465
rect 29368 53456 29420 53508
rect 29552 53456 29604 53508
rect 32036 53456 32088 53508
rect 32956 53456 33008 53508
rect 34520 53456 34572 53508
rect 53564 53499 53616 53508
rect 53564 53465 53573 53499
rect 53573 53465 53607 53499
rect 53607 53465 53616 53499
rect 53564 53456 53616 53465
rect 24492 53431 24544 53440
rect 24492 53397 24501 53431
rect 24501 53397 24535 53431
rect 24535 53397 24544 53431
rect 24492 53388 24544 53397
rect 28172 53388 28224 53440
rect 28816 53431 28868 53440
rect 28816 53397 28825 53431
rect 28825 53397 28859 53431
rect 28859 53397 28868 53431
rect 28816 53388 28868 53397
rect 31668 53388 31720 53440
rect 33508 53431 33560 53440
rect 33508 53397 33517 53431
rect 33517 53397 33551 53431
rect 33551 53397 33560 53431
rect 33784 53431 33836 53440
rect 33508 53388 33560 53397
rect 33784 53397 33793 53431
rect 33793 53397 33827 53431
rect 33827 53397 33836 53431
rect 33784 53388 33836 53397
rect 52460 53388 52512 53440
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 1400 53227 1452 53236
rect 1400 53193 1409 53227
rect 1409 53193 1443 53227
rect 1443 53193 1452 53227
rect 1400 53184 1452 53193
rect 24492 53184 24544 53236
rect 31392 53184 31444 53236
rect 33324 53184 33376 53236
rect 33508 53184 33560 53236
rect 34152 53184 34204 53236
rect 34428 53227 34480 53236
rect 34428 53193 34437 53227
rect 34437 53193 34471 53227
rect 34471 53193 34480 53227
rect 34428 53184 34480 53193
rect 45468 53116 45520 53168
rect 24032 53091 24084 53100
rect 24032 53057 24041 53091
rect 24041 53057 24075 53091
rect 24075 53057 24084 53091
rect 24032 53048 24084 53057
rect 28816 53048 28868 53100
rect 31668 53048 31720 53100
rect 32036 53048 32088 53100
rect 34244 53048 34296 53100
rect 34336 53091 34388 53100
rect 34336 53057 34345 53091
rect 34345 53057 34379 53091
rect 34379 53057 34388 53091
rect 34336 53048 34388 53057
rect 27988 53023 28040 53032
rect 27988 52989 27997 53023
rect 27997 52989 28031 53023
rect 28031 52989 28040 53023
rect 27988 52980 28040 52989
rect 28080 52980 28132 53032
rect 29000 53023 29052 53032
rect 29000 52989 29009 53023
rect 29009 52989 29043 53023
rect 29043 52989 29052 53023
rect 29000 52980 29052 52989
rect 31484 52980 31536 53032
rect 33508 53023 33560 53032
rect 33508 52989 33517 53023
rect 33517 52989 33551 53023
rect 33551 52989 33560 53023
rect 33508 52980 33560 52989
rect 30840 52955 30892 52964
rect 30840 52921 30849 52955
rect 30849 52921 30883 52955
rect 30883 52921 30892 52955
rect 30840 52912 30892 52921
rect 34520 52980 34572 53032
rect 55404 53048 55456 53100
rect 23848 52887 23900 52896
rect 23848 52853 23857 52887
rect 23857 52853 23891 52887
rect 23891 52853 23900 52887
rect 23848 52844 23900 52853
rect 26240 52887 26292 52896
rect 26240 52853 26249 52887
rect 26249 52853 26283 52887
rect 26283 52853 26292 52887
rect 26240 52844 26292 52853
rect 28724 52844 28776 52896
rect 30104 52887 30156 52896
rect 30104 52853 30113 52887
rect 30113 52853 30147 52887
rect 30147 52853 30156 52887
rect 30104 52844 30156 52853
rect 32220 52887 32272 52896
rect 32220 52853 32229 52887
rect 32229 52853 32263 52887
rect 32263 52853 32272 52887
rect 32220 52844 32272 52853
rect 33508 52844 33560 52896
rect 33692 52844 33744 52896
rect 35624 52844 35676 52896
rect 53288 52844 53340 52896
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 29000 52683 29052 52692
rect 29000 52649 29009 52683
rect 29009 52649 29043 52683
rect 29043 52649 29052 52683
rect 29000 52640 29052 52649
rect 31668 52640 31720 52692
rect 34244 52640 34296 52692
rect 35348 52640 35400 52692
rect 1952 52572 2004 52624
rect 24032 52572 24084 52624
rect 27988 52615 28040 52624
rect 1400 52479 1452 52488
rect 1400 52445 1409 52479
rect 1409 52445 1443 52479
rect 1443 52445 1452 52479
rect 1400 52436 1452 52445
rect 23480 52436 23532 52488
rect 25596 52547 25648 52556
rect 25596 52513 25605 52547
rect 25605 52513 25639 52547
rect 25639 52513 25648 52547
rect 25596 52504 25648 52513
rect 23848 52479 23900 52488
rect 23848 52445 23857 52479
rect 23857 52445 23891 52479
rect 23891 52445 23900 52479
rect 23848 52436 23900 52445
rect 24492 52436 24544 52488
rect 26148 52504 26200 52556
rect 27988 52581 27997 52615
rect 27997 52581 28031 52615
rect 28031 52581 28040 52615
rect 27988 52572 28040 52581
rect 29552 52547 29604 52556
rect 29552 52513 29561 52547
rect 29561 52513 29595 52547
rect 29595 52513 29604 52547
rect 29552 52504 29604 52513
rect 32036 52504 32088 52556
rect 26240 52368 26292 52420
rect 27712 52436 27764 52488
rect 28724 52479 28776 52488
rect 28724 52445 28733 52479
rect 28733 52445 28767 52479
rect 28767 52445 28776 52479
rect 28724 52436 28776 52445
rect 28816 52479 28868 52488
rect 28816 52445 28825 52479
rect 28825 52445 28859 52479
rect 28859 52445 28868 52479
rect 28816 52436 28868 52445
rect 29368 52436 29420 52488
rect 29828 52436 29880 52488
rect 30288 52436 30340 52488
rect 30564 52436 30616 52488
rect 33048 52504 33100 52556
rect 33600 52504 33652 52556
rect 29000 52411 29052 52420
rect 29000 52377 29009 52411
rect 29009 52377 29043 52411
rect 29043 52377 29052 52411
rect 29000 52368 29052 52377
rect 30748 52368 30800 52420
rect 33876 52436 33928 52488
rect 34152 52479 34204 52488
rect 23848 52300 23900 52352
rect 27344 52300 27396 52352
rect 33324 52368 33376 52420
rect 34152 52445 34161 52479
rect 34161 52445 34195 52479
rect 34195 52445 34204 52479
rect 34152 52436 34204 52445
rect 35716 52411 35768 52420
rect 35716 52377 35725 52411
rect 35725 52377 35759 52411
rect 35759 52377 35768 52411
rect 35716 52368 35768 52377
rect 33692 52300 33744 52352
rect 34612 52300 34664 52352
rect 35900 52300 35952 52352
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 1400 52139 1452 52148
rect 1400 52105 1409 52139
rect 1409 52105 1443 52139
rect 1443 52105 1452 52139
rect 1400 52096 1452 52105
rect 25596 52096 25648 52148
rect 27712 52096 27764 52148
rect 29828 52139 29880 52148
rect 29828 52105 29837 52139
rect 29837 52105 29871 52139
rect 29871 52105 29880 52139
rect 29828 52096 29880 52105
rect 31300 52139 31352 52148
rect 31300 52105 31309 52139
rect 31309 52105 31343 52139
rect 31343 52105 31352 52139
rect 31300 52096 31352 52105
rect 33416 52096 33468 52148
rect 35348 52139 35400 52148
rect 23480 52028 23532 52080
rect 23756 52071 23808 52080
rect 23756 52037 23765 52071
rect 23765 52037 23799 52071
rect 23799 52037 23808 52071
rect 23756 52028 23808 52037
rect 23572 52003 23624 52012
rect 23572 51969 23581 52003
rect 23581 51969 23615 52003
rect 23615 51969 23624 52003
rect 23572 51960 23624 51969
rect 23664 52003 23716 52012
rect 23664 51969 23673 52003
rect 23673 51969 23707 52003
rect 23707 51969 23716 52003
rect 23664 51960 23716 51969
rect 23848 52003 23900 52012
rect 23848 51969 23857 52003
rect 23857 51969 23891 52003
rect 23891 51969 23900 52003
rect 23848 51960 23900 51969
rect 29460 52071 29512 52080
rect 29460 52037 29469 52071
rect 29469 52037 29503 52071
rect 29503 52037 29512 52071
rect 29460 52028 29512 52037
rect 30104 52028 30156 52080
rect 27988 51960 28040 52012
rect 23204 51892 23256 51944
rect 27620 51935 27672 51944
rect 27620 51901 27629 51935
rect 27629 51901 27663 51935
rect 27663 51901 27672 51935
rect 27620 51892 27672 51901
rect 26240 51824 26292 51876
rect 22836 51799 22888 51808
rect 22836 51765 22845 51799
rect 22845 51765 22879 51799
rect 22879 51765 22888 51799
rect 22836 51756 22888 51765
rect 30012 51960 30064 52012
rect 32220 52028 32272 52080
rect 35348 52105 35357 52139
rect 35357 52105 35391 52139
rect 35391 52105 35400 52139
rect 35348 52096 35400 52105
rect 35716 52096 35768 52148
rect 34152 52028 34204 52080
rect 31760 51960 31812 52012
rect 33324 51960 33376 52012
rect 33692 52003 33744 52012
rect 33692 51969 33701 52003
rect 33701 51969 33735 52003
rect 33735 51969 33744 52003
rect 34520 52003 34572 52012
rect 33692 51960 33744 51969
rect 34520 51969 34529 52003
rect 34529 51969 34563 52003
rect 34563 51969 34572 52003
rect 34520 51960 34572 51969
rect 35532 52003 35584 52012
rect 35532 51969 35541 52003
rect 35541 51969 35575 52003
rect 35575 51969 35584 52003
rect 35532 51960 35584 51969
rect 33140 51892 33192 51944
rect 31484 51867 31536 51876
rect 31484 51833 31493 51867
rect 31493 51833 31527 51867
rect 31527 51833 31536 51867
rect 31484 51824 31536 51833
rect 35348 51892 35400 51944
rect 35900 51892 35952 51944
rect 33600 51824 33652 51876
rect 35624 51824 35676 51876
rect 28724 51799 28776 51808
rect 28724 51765 28733 51799
rect 28733 51765 28767 51799
rect 28767 51765 28776 51799
rect 28724 51756 28776 51765
rect 30748 51756 30800 51808
rect 35440 51756 35492 51808
rect 37280 51799 37332 51808
rect 37280 51765 37289 51799
rect 37289 51765 37323 51799
rect 37323 51765 37332 51799
rect 37280 51756 37332 51765
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 22652 51552 22704 51604
rect 22836 51552 22888 51604
rect 23204 51595 23256 51604
rect 23204 51561 23213 51595
rect 23213 51561 23247 51595
rect 23247 51561 23256 51595
rect 23204 51552 23256 51561
rect 26240 51595 26292 51604
rect 26240 51561 26249 51595
rect 26249 51561 26283 51595
rect 26283 51561 26292 51595
rect 26240 51552 26292 51561
rect 27620 51595 27672 51604
rect 27620 51561 27629 51595
rect 27629 51561 27663 51595
rect 27663 51561 27672 51595
rect 27620 51552 27672 51561
rect 28816 51552 28868 51604
rect 32588 51552 32640 51604
rect 35532 51552 35584 51604
rect 23572 51484 23624 51536
rect 23848 51484 23900 51536
rect 24860 51527 24912 51536
rect 24860 51493 24869 51527
rect 24869 51493 24903 51527
rect 24903 51493 24912 51527
rect 24860 51484 24912 51493
rect 26976 51484 27028 51536
rect 35624 51484 35676 51536
rect 24492 51416 24544 51468
rect 23756 51348 23808 51400
rect 24952 51348 25004 51400
rect 25596 51348 25648 51400
rect 27344 51391 27396 51400
rect 27344 51357 27353 51391
rect 27353 51357 27387 51391
rect 27387 51357 27396 51391
rect 27344 51348 27396 51357
rect 28816 51348 28868 51400
rect 30748 51416 30800 51468
rect 36452 51416 36504 51468
rect 30840 51391 30892 51400
rect 30840 51357 30849 51391
rect 30849 51357 30883 51391
rect 30883 51357 30892 51391
rect 30840 51348 30892 51357
rect 31300 51391 31352 51400
rect 31300 51357 31309 51391
rect 31309 51357 31343 51391
rect 31343 51357 31352 51391
rect 31300 51348 31352 51357
rect 33508 51391 33560 51400
rect 22560 51280 22612 51332
rect 23664 51280 23716 51332
rect 27252 51280 27304 51332
rect 26148 51212 26200 51264
rect 27528 51212 27580 51264
rect 30012 51280 30064 51332
rect 33508 51357 33517 51391
rect 33517 51357 33551 51391
rect 33551 51357 33560 51391
rect 33508 51348 33560 51357
rect 33784 51391 33836 51400
rect 33784 51357 33793 51391
rect 33793 51357 33827 51391
rect 33827 51357 33836 51391
rect 33784 51348 33836 51357
rect 34704 51391 34756 51400
rect 34704 51357 34713 51391
rect 34713 51357 34747 51391
rect 34747 51357 34756 51391
rect 34704 51348 34756 51357
rect 35716 51348 35768 51400
rect 33140 51280 33192 51332
rect 34336 51280 34388 51332
rect 34888 51323 34940 51332
rect 34888 51289 34897 51323
rect 34897 51289 34931 51323
rect 34931 51289 34940 51323
rect 34888 51280 34940 51289
rect 29828 51212 29880 51264
rect 31392 51255 31444 51264
rect 31392 51221 31401 51255
rect 31401 51221 31435 51255
rect 31435 51221 31444 51255
rect 31392 51212 31444 51221
rect 31944 51255 31996 51264
rect 31944 51221 31953 51255
rect 31953 51221 31987 51255
rect 31987 51221 31996 51255
rect 31944 51212 31996 51221
rect 32588 51255 32640 51264
rect 32588 51221 32597 51255
rect 32597 51221 32631 51255
rect 32631 51221 32640 51255
rect 32588 51212 32640 51221
rect 35532 51212 35584 51264
rect 37188 51212 37240 51264
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 23848 51051 23900 51060
rect 23848 51017 23857 51051
rect 23857 51017 23891 51051
rect 23891 51017 23900 51051
rect 23848 51008 23900 51017
rect 26056 51008 26108 51060
rect 31300 51008 31352 51060
rect 31760 51008 31812 51060
rect 35716 51008 35768 51060
rect 1400 50915 1452 50924
rect 1400 50881 1409 50915
rect 1409 50881 1443 50915
rect 1443 50881 1452 50915
rect 1400 50872 1452 50881
rect 22560 50915 22612 50924
rect 22560 50881 22569 50915
rect 22569 50881 22603 50915
rect 22603 50881 22612 50915
rect 22560 50872 22612 50881
rect 22744 50915 22796 50924
rect 22744 50881 22753 50915
rect 22753 50881 22787 50915
rect 22787 50881 22796 50915
rect 22744 50872 22796 50881
rect 23204 50915 23256 50924
rect 23204 50881 23213 50915
rect 23213 50881 23247 50915
rect 23247 50881 23256 50915
rect 23204 50872 23256 50881
rect 24492 50940 24544 50992
rect 30012 50983 30064 50992
rect 30012 50949 30021 50983
rect 30021 50949 30055 50983
rect 30055 50949 30064 50983
rect 30012 50940 30064 50949
rect 30380 50940 30432 50992
rect 23940 50872 23992 50924
rect 25136 50872 25188 50924
rect 25596 50872 25648 50924
rect 25872 50915 25924 50924
rect 25872 50881 25881 50915
rect 25881 50881 25915 50915
rect 25915 50881 25924 50915
rect 25872 50872 25924 50881
rect 30288 50915 30340 50924
rect 30288 50881 30297 50915
rect 30297 50881 30331 50915
rect 30331 50881 30340 50915
rect 30288 50872 30340 50881
rect 30840 50872 30892 50924
rect 32404 50915 32456 50924
rect 32404 50881 32413 50915
rect 32413 50881 32447 50915
rect 32447 50881 32456 50915
rect 32404 50872 32456 50881
rect 34888 50915 34940 50924
rect 34888 50881 34897 50915
rect 34897 50881 34931 50915
rect 34931 50881 34940 50915
rect 34888 50872 34940 50881
rect 35900 50872 35952 50924
rect 53564 50915 53616 50924
rect 53564 50881 53573 50915
rect 53573 50881 53607 50915
rect 53607 50881 53616 50915
rect 53564 50872 53616 50881
rect 24952 50847 25004 50856
rect 24952 50813 24961 50847
rect 24961 50813 24995 50847
rect 24995 50813 25004 50847
rect 24952 50804 25004 50813
rect 26148 50847 26200 50856
rect 26148 50813 26157 50847
rect 26157 50813 26191 50847
rect 26191 50813 26200 50847
rect 26148 50804 26200 50813
rect 30748 50847 30800 50856
rect 30748 50813 30757 50847
rect 30757 50813 30791 50847
rect 30791 50813 30800 50847
rect 30748 50804 30800 50813
rect 32496 50804 32548 50856
rect 34520 50847 34572 50856
rect 34520 50813 34529 50847
rect 34529 50813 34563 50847
rect 34563 50813 34572 50847
rect 34520 50804 34572 50813
rect 34704 50804 34756 50856
rect 35348 50804 35400 50856
rect 1768 50668 1820 50720
rect 22008 50711 22060 50720
rect 22008 50677 22017 50711
rect 22017 50677 22051 50711
rect 22051 50677 22060 50711
rect 25780 50736 25832 50788
rect 22008 50668 22060 50677
rect 23480 50668 23532 50720
rect 23756 50668 23808 50720
rect 24032 50668 24084 50720
rect 26240 50668 26292 50720
rect 26884 50668 26936 50720
rect 28724 50736 28776 50788
rect 35900 50736 35952 50788
rect 37188 50736 37240 50788
rect 28908 50668 28960 50720
rect 29276 50668 29328 50720
rect 30104 50668 30156 50720
rect 32220 50711 32272 50720
rect 32220 50677 32229 50711
rect 32229 50677 32263 50711
rect 32263 50677 32272 50711
rect 32220 50668 32272 50677
rect 32312 50711 32364 50720
rect 32312 50677 32321 50711
rect 32321 50677 32355 50711
rect 32355 50677 32364 50711
rect 32312 50668 32364 50677
rect 33784 50668 33836 50720
rect 37280 50668 37332 50720
rect 53472 50711 53524 50720
rect 53472 50677 53481 50711
rect 53481 50677 53515 50711
rect 53515 50677 53524 50711
rect 53472 50668 53524 50677
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 22560 50464 22612 50516
rect 24952 50464 25004 50516
rect 27160 50507 27212 50516
rect 27160 50473 27169 50507
rect 27169 50473 27203 50507
rect 27203 50473 27212 50507
rect 27160 50464 27212 50473
rect 30288 50507 30340 50516
rect 30288 50473 30297 50507
rect 30297 50473 30331 50507
rect 30331 50473 30340 50507
rect 30288 50464 30340 50473
rect 1400 50439 1452 50448
rect 1400 50405 1409 50439
rect 1409 50405 1443 50439
rect 1443 50405 1452 50439
rect 1400 50396 1452 50405
rect 23480 50396 23532 50448
rect 25780 50371 25832 50380
rect 25780 50337 25789 50371
rect 25789 50337 25823 50371
rect 25823 50337 25832 50371
rect 25780 50328 25832 50337
rect 26516 50328 26568 50380
rect 27528 50328 27580 50380
rect 29276 50328 29328 50380
rect 30380 50371 30432 50380
rect 30380 50337 30389 50371
rect 30389 50337 30423 50371
rect 30423 50337 30432 50371
rect 30380 50328 30432 50337
rect 31024 50328 31076 50380
rect 22008 50260 22060 50312
rect 22652 50303 22704 50312
rect 22652 50269 22661 50303
rect 22661 50269 22695 50303
rect 22695 50269 22704 50303
rect 22652 50260 22704 50269
rect 23204 50260 23256 50312
rect 25872 50303 25924 50312
rect 25872 50269 25881 50303
rect 25881 50269 25915 50303
rect 25915 50269 25924 50303
rect 25872 50260 25924 50269
rect 26700 50303 26752 50312
rect 26700 50269 26709 50303
rect 26709 50269 26743 50303
rect 26743 50269 26752 50303
rect 26700 50260 26752 50269
rect 26792 50303 26844 50312
rect 26792 50269 26801 50303
rect 26801 50269 26835 50303
rect 26835 50269 26844 50303
rect 26792 50260 26844 50269
rect 26976 50303 27028 50312
rect 26976 50269 26985 50303
rect 26985 50269 27019 50303
rect 27019 50269 27028 50303
rect 30104 50303 30156 50312
rect 26976 50260 27028 50269
rect 30104 50269 30113 50303
rect 30113 50269 30147 50303
rect 30147 50269 30156 50303
rect 30104 50260 30156 50269
rect 31300 50328 31352 50380
rect 31392 50303 31444 50312
rect 23572 50192 23624 50244
rect 24860 50235 24912 50244
rect 24860 50201 24869 50235
rect 24869 50201 24903 50235
rect 24903 50201 24912 50235
rect 24860 50192 24912 50201
rect 21640 50124 21692 50176
rect 24032 50124 24084 50176
rect 24676 50124 24728 50176
rect 25504 50192 25556 50244
rect 28172 50192 28224 50244
rect 31392 50269 31401 50303
rect 31401 50269 31435 50303
rect 31435 50269 31444 50303
rect 31392 50260 31444 50269
rect 32404 50464 32456 50516
rect 37188 50464 37240 50516
rect 53472 50464 53524 50516
rect 33324 50396 33376 50448
rect 32312 50260 32364 50312
rect 32496 50303 32548 50312
rect 32496 50269 32505 50303
rect 32505 50269 32539 50303
rect 32539 50269 32548 50303
rect 32496 50260 32548 50269
rect 34612 50328 34664 50380
rect 33784 50260 33836 50312
rect 34152 50303 34204 50312
rect 34152 50269 34161 50303
rect 34161 50269 34195 50303
rect 34195 50269 34204 50303
rect 34152 50260 34204 50269
rect 34336 50192 34388 50244
rect 53380 50192 53432 50244
rect 26240 50124 26292 50176
rect 28908 50167 28960 50176
rect 28908 50133 28917 50167
rect 28917 50133 28951 50167
rect 28951 50133 28960 50167
rect 28908 50124 28960 50133
rect 29920 50167 29972 50176
rect 29920 50133 29929 50167
rect 29929 50133 29963 50167
rect 29963 50133 29972 50167
rect 29920 50124 29972 50133
rect 31024 50124 31076 50176
rect 31392 50124 31444 50176
rect 32404 50124 32456 50176
rect 34428 50124 34480 50176
rect 35348 50124 35400 50176
rect 37280 50124 37332 50176
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 22744 49963 22796 49972
rect 22744 49929 22753 49963
rect 22753 49929 22787 49963
rect 22787 49929 22796 49963
rect 22744 49920 22796 49929
rect 24492 49920 24544 49972
rect 21640 49784 21692 49836
rect 22652 49827 22704 49836
rect 22652 49793 22661 49827
rect 22661 49793 22695 49827
rect 22695 49793 22704 49827
rect 22652 49784 22704 49793
rect 24768 49852 24820 49904
rect 26792 49920 26844 49972
rect 31024 49895 31076 49904
rect 31024 49861 31033 49895
rect 31033 49861 31067 49895
rect 31067 49861 31076 49895
rect 31024 49852 31076 49861
rect 32496 49920 32548 49972
rect 34152 49920 34204 49972
rect 22008 49716 22060 49768
rect 24032 49784 24084 49836
rect 24308 49827 24360 49836
rect 24308 49793 24317 49827
rect 24317 49793 24351 49827
rect 24351 49793 24360 49827
rect 24308 49784 24360 49793
rect 24492 49827 24544 49836
rect 24492 49793 24501 49827
rect 24501 49793 24535 49827
rect 24535 49793 24544 49827
rect 24492 49784 24544 49793
rect 24860 49784 24912 49836
rect 25504 49827 25556 49836
rect 25504 49793 25513 49827
rect 25513 49793 25547 49827
rect 25547 49793 25556 49827
rect 25504 49784 25556 49793
rect 26240 49827 26292 49836
rect 26240 49793 26249 49827
rect 26249 49793 26283 49827
rect 26283 49793 26292 49827
rect 26240 49784 26292 49793
rect 29736 49827 29788 49836
rect 29736 49793 29754 49827
rect 29754 49793 29788 49827
rect 29736 49784 29788 49793
rect 30288 49784 30340 49836
rect 31300 49784 31352 49836
rect 32128 49827 32180 49836
rect 32128 49793 32137 49827
rect 32137 49793 32171 49827
rect 32171 49793 32180 49827
rect 32128 49784 32180 49793
rect 33784 49852 33836 49904
rect 34428 49895 34480 49904
rect 34428 49861 34437 49895
rect 34437 49861 34471 49895
rect 34471 49861 34480 49895
rect 34428 49852 34480 49861
rect 34612 49895 34664 49904
rect 34612 49861 34621 49895
rect 34621 49861 34655 49895
rect 34655 49861 34664 49895
rect 34612 49852 34664 49861
rect 34336 49784 34388 49836
rect 25872 49716 25924 49768
rect 27620 49716 27672 49768
rect 28080 49759 28132 49768
rect 28080 49725 28089 49759
rect 28089 49725 28123 49759
rect 28123 49725 28132 49759
rect 28080 49716 28132 49725
rect 30012 49759 30064 49768
rect 30012 49725 30021 49759
rect 30021 49725 30055 49759
rect 30055 49725 30064 49759
rect 30012 49716 30064 49725
rect 32588 49716 32640 49768
rect 33048 49716 33100 49768
rect 52460 49920 52512 49972
rect 36912 49716 36964 49768
rect 37280 49716 37332 49768
rect 23848 49648 23900 49700
rect 23480 49580 23532 49632
rect 24492 49580 24544 49632
rect 29368 49580 29420 49632
rect 30748 49580 30800 49632
rect 33784 49580 33836 49632
rect 35532 49580 35584 49632
rect 35900 49580 35952 49632
rect 36176 49623 36228 49632
rect 36176 49589 36185 49623
rect 36185 49589 36219 49623
rect 36219 49589 36228 49623
rect 36176 49580 36228 49589
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 25412 49376 25464 49428
rect 29736 49376 29788 49428
rect 32588 49376 32640 49428
rect 24860 49308 24912 49360
rect 29920 49308 29972 49360
rect 23664 49240 23716 49292
rect 23940 49240 23992 49292
rect 23480 49215 23532 49224
rect 23480 49181 23489 49215
rect 23489 49181 23523 49215
rect 23523 49181 23532 49215
rect 23480 49172 23532 49181
rect 24400 49215 24452 49224
rect 24400 49181 24409 49215
rect 24409 49181 24443 49215
rect 24443 49181 24452 49215
rect 24400 49172 24452 49181
rect 24492 49215 24544 49224
rect 24492 49181 24501 49215
rect 24501 49181 24535 49215
rect 24535 49181 24544 49215
rect 24492 49172 24544 49181
rect 25504 49215 25556 49224
rect 23756 49104 23808 49156
rect 25504 49181 25513 49215
rect 25513 49181 25547 49215
rect 25547 49181 25556 49215
rect 25504 49172 25556 49181
rect 31944 49308 31996 49360
rect 33048 49308 33100 49360
rect 32496 49283 32548 49292
rect 22008 49036 22060 49088
rect 25044 49104 25096 49156
rect 27896 49172 27948 49224
rect 25320 49036 25372 49088
rect 26056 49036 26108 49088
rect 26240 49036 26292 49088
rect 26884 49104 26936 49156
rect 28540 49172 28592 49224
rect 29552 49172 29604 49224
rect 29736 49215 29788 49224
rect 29736 49181 29745 49215
rect 29745 49181 29779 49215
rect 29779 49181 29788 49215
rect 29736 49172 29788 49181
rect 29828 49172 29880 49224
rect 32496 49249 32505 49283
rect 32505 49249 32539 49283
rect 32539 49249 32548 49283
rect 32496 49240 32548 49249
rect 32588 49240 32640 49292
rect 31760 49172 31812 49224
rect 32220 49172 32272 49224
rect 32404 49215 32456 49224
rect 32404 49181 32413 49215
rect 32413 49181 32447 49215
rect 32447 49181 32456 49215
rect 32680 49215 32732 49224
rect 32404 49172 32456 49181
rect 32680 49181 32689 49215
rect 32689 49181 32723 49215
rect 32723 49181 32732 49215
rect 32680 49172 32732 49181
rect 33232 49172 33284 49224
rect 33508 49215 33560 49224
rect 33508 49181 33517 49215
rect 33517 49181 33551 49215
rect 33551 49181 33560 49215
rect 33508 49172 33560 49181
rect 33600 49215 33652 49224
rect 33600 49181 33609 49215
rect 33609 49181 33643 49215
rect 33643 49181 33652 49215
rect 35256 49240 35308 49292
rect 33600 49172 33652 49181
rect 32496 49104 32548 49156
rect 34336 49104 34388 49156
rect 35900 49172 35952 49224
rect 37188 49376 37240 49428
rect 26792 49036 26844 49088
rect 28080 49036 28132 49088
rect 28448 49036 28500 49088
rect 28816 49079 28868 49088
rect 28816 49045 28825 49079
rect 28825 49045 28859 49079
rect 28859 49045 28868 49079
rect 28816 49036 28868 49045
rect 29552 49036 29604 49088
rect 31116 49036 31168 49088
rect 33416 49036 33468 49088
rect 34612 49036 34664 49088
rect 35900 49036 35952 49088
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 23572 48832 23624 48884
rect 28264 48832 28316 48884
rect 33600 48832 33652 48884
rect 24492 48764 24544 48816
rect 23848 48739 23900 48748
rect 23848 48705 23857 48739
rect 23857 48705 23891 48739
rect 23891 48705 23900 48739
rect 23848 48696 23900 48705
rect 24860 48739 24912 48748
rect 23664 48671 23716 48680
rect 23664 48637 23673 48671
rect 23673 48637 23707 48671
rect 23707 48637 23716 48671
rect 23664 48628 23716 48637
rect 22928 48603 22980 48612
rect 22928 48569 22937 48603
rect 22937 48569 22971 48603
rect 22971 48569 22980 48603
rect 22928 48560 22980 48569
rect 23572 48560 23624 48612
rect 23940 48671 23992 48680
rect 23940 48637 23949 48671
rect 23949 48637 23983 48671
rect 23983 48637 23992 48671
rect 23940 48628 23992 48637
rect 24032 48560 24084 48612
rect 24860 48705 24869 48739
rect 24869 48705 24903 48739
rect 24903 48705 24912 48739
rect 24860 48696 24912 48705
rect 25136 48764 25188 48816
rect 26240 48739 26292 48748
rect 26240 48705 26249 48739
rect 26249 48705 26283 48739
rect 26283 48705 26292 48739
rect 26240 48696 26292 48705
rect 26884 48696 26936 48748
rect 29276 48764 29328 48816
rect 28356 48696 28408 48748
rect 28816 48696 28868 48748
rect 29552 48696 29604 48748
rect 30196 48739 30248 48748
rect 30196 48705 30205 48739
rect 30205 48705 30239 48739
rect 30239 48705 30248 48739
rect 30196 48696 30248 48705
rect 30840 48739 30892 48748
rect 25412 48628 25464 48680
rect 26608 48628 26660 48680
rect 26792 48628 26844 48680
rect 27712 48628 27764 48680
rect 28448 48671 28500 48680
rect 28448 48637 28457 48671
rect 28457 48637 28491 48671
rect 28491 48637 28500 48671
rect 28448 48628 28500 48637
rect 25044 48560 25096 48612
rect 27528 48603 27580 48612
rect 26332 48535 26384 48544
rect 26332 48501 26341 48535
rect 26341 48501 26375 48535
rect 26375 48501 26384 48535
rect 26332 48492 26384 48501
rect 27528 48569 27537 48603
rect 27537 48569 27571 48603
rect 27571 48569 27580 48603
rect 27528 48560 27580 48569
rect 29736 48628 29788 48680
rect 30840 48705 30849 48739
rect 30849 48705 30883 48739
rect 30883 48705 30892 48739
rect 30840 48696 30892 48705
rect 31024 48739 31076 48748
rect 31024 48705 31033 48739
rect 31033 48705 31067 48739
rect 31067 48705 31076 48739
rect 31024 48696 31076 48705
rect 29184 48560 29236 48612
rect 31300 48560 31352 48612
rect 29368 48535 29420 48544
rect 29368 48501 29377 48535
rect 29377 48501 29411 48535
rect 29411 48501 29420 48535
rect 29368 48492 29420 48501
rect 29920 48492 29972 48544
rect 30932 48535 30984 48544
rect 30932 48501 30941 48535
rect 30941 48501 30975 48535
rect 30975 48501 30984 48535
rect 30932 48492 30984 48501
rect 31484 48535 31536 48544
rect 31484 48501 31493 48535
rect 31493 48501 31527 48535
rect 31527 48501 31536 48535
rect 31484 48492 31536 48501
rect 33784 48764 33836 48816
rect 34244 48764 34296 48816
rect 34612 48807 34664 48816
rect 34612 48773 34621 48807
rect 34621 48773 34655 48807
rect 34655 48773 34664 48807
rect 34612 48764 34664 48773
rect 35256 48739 35308 48748
rect 35256 48705 35265 48739
rect 35265 48705 35299 48739
rect 35299 48705 35308 48739
rect 35256 48696 35308 48705
rect 53564 48739 53616 48748
rect 53564 48705 53573 48739
rect 53573 48705 53607 48739
rect 53607 48705 53616 48739
rect 53564 48696 53616 48705
rect 35532 48628 35584 48680
rect 33508 48560 33560 48612
rect 53104 48560 53156 48612
rect 33600 48492 33652 48544
rect 34796 48492 34848 48544
rect 35532 48492 35584 48544
rect 35808 48492 35860 48544
rect 36544 48492 36596 48544
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 24860 48288 24912 48340
rect 29828 48288 29880 48340
rect 30104 48288 30156 48340
rect 31484 48288 31536 48340
rect 24032 48220 24084 48272
rect 25044 48220 25096 48272
rect 24308 48152 24360 48204
rect 26424 48195 26476 48204
rect 20168 48084 20220 48136
rect 22928 48084 22980 48136
rect 26424 48161 26433 48195
rect 26433 48161 26467 48195
rect 26467 48161 26476 48195
rect 26424 48152 26476 48161
rect 2228 48059 2280 48068
rect 2228 48025 2237 48059
rect 2237 48025 2271 48059
rect 2271 48025 2280 48059
rect 2228 48016 2280 48025
rect 23848 48016 23900 48068
rect 24860 48084 24912 48136
rect 26332 48127 26384 48136
rect 26332 48093 26341 48127
rect 26341 48093 26375 48127
rect 26375 48093 26384 48127
rect 26332 48084 26384 48093
rect 27252 48220 27304 48272
rect 30196 48220 30248 48272
rect 27528 48127 27580 48136
rect 27528 48093 27537 48127
rect 27537 48093 27571 48127
rect 27571 48093 27580 48127
rect 27528 48084 27580 48093
rect 28908 48152 28960 48204
rect 29920 48195 29972 48204
rect 29920 48161 29929 48195
rect 29929 48161 29963 48195
rect 29963 48161 29972 48195
rect 29920 48152 29972 48161
rect 28172 48084 28224 48136
rect 28356 48127 28408 48136
rect 28356 48093 28365 48127
rect 28365 48093 28399 48127
rect 28399 48093 28408 48127
rect 28356 48084 28408 48093
rect 28540 48127 28592 48136
rect 28540 48093 28549 48127
rect 28549 48093 28583 48127
rect 28583 48093 28592 48127
rect 28540 48084 28592 48093
rect 28632 48127 28684 48136
rect 28632 48093 28641 48127
rect 28641 48093 28675 48127
rect 28675 48093 28684 48127
rect 28632 48084 28684 48093
rect 29276 48084 29328 48136
rect 30288 48084 30340 48136
rect 30932 48127 30984 48136
rect 30932 48093 30941 48127
rect 30941 48093 30975 48127
rect 30975 48093 30984 48127
rect 30932 48084 30984 48093
rect 31116 48127 31168 48136
rect 31116 48093 31125 48127
rect 31125 48093 31159 48127
rect 31159 48093 31168 48127
rect 31116 48084 31168 48093
rect 32220 48220 32272 48272
rect 32404 48152 32456 48204
rect 35348 48152 35400 48204
rect 35808 48152 35860 48204
rect 32588 48084 32640 48136
rect 33232 48084 33284 48136
rect 34428 48084 34480 48136
rect 33048 48016 33100 48068
rect 34244 48016 34296 48068
rect 1492 47991 1544 48000
rect 1492 47957 1501 47991
rect 1501 47957 1535 47991
rect 1535 47957 1544 47991
rect 1492 47948 1544 47957
rect 20720 47991 20772 48000
rect 20720 47957 20729 47991
rect 20729 47957 20763 47991
rect 20763 47957 20772 47991
rect 20720 47948 20772 47957
rect 22008 47948 22060 48000
rect 23112 47948 23164 48000
rect 26240 47948 26292 48000
rect 29920 47948 29972 48000
rect 31760 47948 31812 48000
rect 33140 47991 33192 48000
rect 33140 47957 33149 47991
rect 33149 47957 33183 47991
rect 33183 47957 33192 47991
rect 33140 47948 33192 47957
rect 34612 47948 34664 48000
rect 35532 48016 35584 48068
rect 36544 48084 36596 48136
rect 36544 47948 36596 48000
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 23940 47744 23992 47796
rect 24032 47787 24084 47796
rect 24032 47753 24041 47787
rect 24041 47753 24075 47787
rect 24075 47753 24084 47787
rect 24032 47744 24084 47753
rect 25688 47744 25740 47796
rect 26424 47787 26476 47796
rect 21548 47676 21600 47728
rect 22008 47676 22060 47728
rect 20168 47608 20220 47660
rect 22284 47651 22336 47660
rect 22284 47617 22293 47651
rect 22293 47617 22327 47651
rect 22327 47617 22336 47651
rect 22284 47608 22336 47617
rect 25504 47719 25556 47728
rect 25504 47685 25513 47719
rect 25513 47685 25547 47719
rect 25547 47685 25556 47719
rect 25504 47676 25556 47685
rect 26424 47753 26433 47787
rect 26433 47753 26467 47787
rect 26467 47753 26476 47787
rect 26424 47744 26476 47753
rect 29000 47787 29052 47796
rect 29000 47753 29009 47787
rect 29009 47753 29043 47787
rect 29043 47753 29052 47787
rect 29000 47744 29052 47753
rect 30840 47744 30892 47796
rect 32588 47744 32640 47796
rect 34428 47744 34480 47796
rect 20720 47540 20772 47592
rect 25136 47651 25188 47660
rect 25136 47617 25145 47651
rect 25145 47617 25179 47651
rect 25179 47617 25188 47651
rect 25136 47608 25188 47617
rect 26056 47651 26108 47660
rect 26056 47617 26065 47651
rect 26065 47617 26099 47651
rect 26099 47617 26108 47651
rect 26056 47608 26108 47617
rect 22284 47472 22336 47524
rect 23388 47540 23440 47592
rect 25320 47540 25372 47592
rect 25872 47540 25924 47592
rect 23664 47472 23716 47524
rect 27160 47608 27212 47660
rect 27436 47608 27488 47660
rect 27896 47676 27948 47728
rect 28632 47676 28684 47728
rect 29276 47719 29328 47728
rect 29276 47685 29285 47719
rect 29285 47685 29319 47719
rect 29319 47685 29328 47719
rect 29276 47676 29328 47685
rect 31300 47676 31352 47728
rect 29184 47651 29236 47660
rect 29184 47617 29188 47651
rect 29188 47617 29222 47651
rect 29222 47617 29236 47651
rect 29184 47608 29236 47617
rect 29368 47651 29420 47660
rect 29368 47617 29377 47651
rect 29377 47617 29411 47651
rect 29411 47617 29420 47651
rect 29368 47608 29420 47617
rect 20168 47447 20220 47456
rect 20168 47413 20177 47447
rect 20177 47413 20211 47447
rect 20211 47413 20220 47447
rect 20168 47404 20220 47413
rect 20720 47447 20772 47456
rect 20720 47413 20729 47447
rect 20729 47413 20763 47447
rect 20763 47413 20772 47447
rect 20720 47404 20772 47413
rect 21548 47404 21600 47456
rect 26056 47404 26108 47456
rect 28908 47540 28960 47592
rect 30564 47608 30616 47660
rect 31024 47651 31076 47660
rect 31024 47617 31033 47651
rect 31033 47617 31067 47651
rect 31067 47617 31076 47651
rect 31024 47608 31076 47617
rect 31116 47540 31168 47592
rect 32036 47608 32088 47660
rect 33784 47676 33836 47728
rect 32404 47608 32456 47660
rect 33048 47608 33100 47660
rect 33232 47651 33284 47660
rect 33232 47617 33241 47651
rect 33241 47617 33275 47651
rect 33275 47617 33284 47651
rect 33416 47651 33468 47660
rect 33232 47608 33284 47617
rect 33416 47617 33425 47651
rect 33425 47617 33459 47651
rect 33459 47617 33468 47651
rect 33416 47608 33468 47617
rect 34796 47608 34848 47660
rect 35348 47651 35400 47660
rect 35348 47617 35357 47651
rect 35357 47617 35391 47651
rect 35391 47617 35400 47651
rect 35348 47608 35400 47617
rect 33508 47540 33560 47592
rect 34612 47583 34664 47592
rect 34612 47549 34621 47583
rect 34621 47549 34655 47583
rect 34655 47549 34664 47583
rect 34612 47540 34664 47549
rect 26608 47472 26660 47524
rect 33232 47472 33284 47524
rect 35348 47472 35400 47524
rect 28540 47447 28592 47456
rect 28540 47413 28549 47447
rect 28549 47413 28583 47447
rect 28583 47413 28592 47447
rect 28540 47404 28592 47413
rect 33692 47447 33744 47456
rect 33692 47413 33701 47447
rect 33701 47413 33735 47447
rect 33735 47413 33744 47447
rect 33692 47404 33744 47413
rect 35808 47447 35860 47456
rect 35808 47413 35817 47447
rect 35817 47413 35851 47447
rect 35851 47413 35860 47447
rect 35808 47404 35860 47413
rect 37464 47404 37516 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 24676 47200 24728 47252
rect 26424 47200 26476 47252
rect 26976 47200 27028 47252
rect 24400 47132 24452 47184
rect 25228 47132 25280 47184
rect 25504 47132 25556 47184
rect 23388 47064 23440 47116
rect 24584 47064 24636 47116
rect 20168 46996 20220 47048
rect 23572 46996 23624 47048
rect 24676 46996 24728 47048
rect 24952 47039 25004 47048
rect 24952 47005 24961 47039
rect 24961 47005 24995 47039
rect 24995 47005 25004 47039
rect 24952 46996 25004 47005
rect 25044 46996 25096 47048
rect 20628 46928 20680 46980
rect 22468 46928 22520 46980
rect 25780 46996 25832 47048
rect 26240 47039 26292 47048
rect 26240 47005 26249 47039
rect 26249 47005 26283 47039
rect 26283 47005 26292 47039
rect 26240 46996 26292 47005
rect 19340 46860 19392 46912
rect 21824 46903 21876 46912
rect 21824 46869 21833 46903
rect 21833 46869 21867 46903
rect 21867 46869 21876 46903
rect 21824 46860 21876 46869
rect 22376 46903 22428 46912
rect 22376 46869 22385 46903
rect 22385 46869 22419 46903
rect 22419 46869 22428 46903
rect 22376 46860 22428 46869
rect 26240 46860 26292 46912
rect 26424 47039 26476 47048
rect 26424 47005 26433 47039
rect 26433 47005 26467 47039
rect 26467 47005 26476 47039
rect 27160 47039 27212 47048
rect 26424 46996 26476 47005
rect 27160 47005 27169 47039
rect 27169 47005 27203 47039
rect 27203 47005 27212 47039
rect 27160 46996 27212 47005
rect 29368 47200 29420 47252
rect 30288 47243 30340 47252
rect 30288 47209 30297 47243
rect 30297 47209 30331 47243
rect 30331 47209 30340 47243
rect 30288 47200 30340 47209
rect 30840 47200 30892 47252
rect 32680 47200 32732 47252
rect 28908 47132 28960 47184
rect 33784 47200 33836 47252
rect 35808 47200 35860 47252
rect 35348 47175 35400 47184
rect 27712 47064 27764 47116
rect 28540 47064 28592 47116
rect 29000 47064 29052 47116
rect 29460 47064 29512 47116
rect 30196 47064 30248 47116
rect 32496 47107 32548 47116
rect 27436 47039 27488 47048
rect 27436 47005 27445 47039
rect 27445 47005 27479 47039
rect 27479 47005 27488 47039
rect 27436 46996 27488 47005
rect 29552 46996 29604 47048
rect 27620 46928 27672 46980
rect 28448 46928 28500 46980
rect 29184 46928 29236 46980
rect 30748 46996 30800 47048
rect 32496 47073 32505 47107
rect 32505 47073 32539 47107
rect 32539 47073 32548 47107
rect 32496 47064 32548 47073
rect 31300 46996 31352 47048
rect 32220 47039 32272 47048
rect 32220 47005 32229 47039
rect 32229 47005 32263 47039
rect 32263 47005 32272 47039
rect 32220 46996 32272 47005
rect 33232 47064 33284 47116
rect 35348 47141 35357 47175
rect 35357 47141 35391 47175
rect 35391 47141 35400 47175
rect 35348 47132 35400 47141
rect 33140 47039 33192 47048
rect 33140 47005 33144 47039
rect 33144 47005 33178 47039
rect 33178 47005 33192 47039
rect 37188 47064 37240 47116
rect 33140 46996 33192 47005
rect 33968 46996 34020 47048
rect 30656 46928 30708 46980
rect 30932 46971 30984 46980
rect 30932 46937 30941 46971
rect 30941 46937 30975 46971
rect 30975 46937 30984 46971
rect 30932 46928 30984 46937
rect 31668 46971 31720 46980
rect 31668 46937 31677 46971
rect 31677 46937 31711 46971
rect 31711 46937 31720 46971
rect 31668 46928 31720 46937
rect 33232 46971 33284 46980
rect 33232 46937 33241 46971
rect 33241 46937 33275 46971
rect 33275 46937 33284 46971
rect 33232 46928 33284 46937
rect 33324 46971 33376 46980
rect 33324 46937 33333 46971
rect 33333 46937 33367 46971
rect 33367 46937 33376 46971
rect 33324 46928 33376 46937
rect 34060 46928 34112 46980
rect 30840 46860 30892 46912
rect 33140 46860 33192 46912
rect 34612 46860 34664 46912
rect 36544 46860 36596 46912
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 22100 46656 22152 46708
rect 22376 46656 22428 46708
rect 23756 46656 23808 46708
rect 24860 46656 24912 46708
rect 25228 46656 25280 46708
rect 29184 46699 29236 46708
rect 29184 46665 29193 46699
rect 29193 46665 29227 46699
rect 29227 46665 29236 46699
rect 29184 46656 29236 46665
rect 30196 46656 30248 46708
rect 30748 46699 30800 46708
rect 30748 46665 30757 46699
rect 30757 46665 30791 46699
rect 30791 46665 30800 46699
rect 30748 46656 30800 46665
rect 31208 46656 31260 46708
rect 33324 46656 33376 46708
rect 34060 46699 34112 46708
rect 34060 46665 34069 46699
rect 34069 46665 34103 46699
rect 34103 46665 34112 46699
rect 34060 46656 34112 46665
rect 26240 46588 26292 46640
rect 23388 46563 23440 46572
rect 23388 46529 23397 46563
rect 23397 46529 23431 46563
rect 23431 46529 23440 46563
rect 23388 46520 23440 46529
rect 23572 46563 23624 46572
rect 23572 46529 23581 46563
rect 23581 46529 23615 46563
rect 23615 46529 23624 46563
rect 23572 46520 23624 46529
rect 24400 46520 24452 46572
rect 25688 46563 25740 46572
rect 25688 46529 25697 46563
rect 25697 46529 25731 46563
rect 25731 46529 25740 46563
rect 25688 46520 25740 46529
rect 25872 46563 25924 46572
rect 25872 46529 25881 46563
rect 25881 46529 25915 46563
rect 25915 46529 25924 46563
rect 25872 46520 25924 46529
rect 26516 46520 26568 46572
rect 27528 46588 27580 46640
rect 29460 46588 29512 46640
rect 29920 46631 29972 46640
rect 29920 46597 29929 46631
rect 29929 46597 29963 46631
rect 29963 46597 29972 46631
rect 29920 46588 29972 46597
rect 32956 46588 33008 46640
rect 35440 46588 35492 46640
rect 29736 46520 29788 46572
rect 29828 46563 29880 46572
rect 29828 46529 29837 46563
rect 29837 46529 29871 46563
rect 29871 46529 29880 46563
rect 29828 46520 29880 46529
rect 30104 46520 30156 46572
rect 30840 46563 30892 46572
rect 21824 46452 21876 46504
rect 22284 46452 22336 46504
rect 24492 46452 24544 46504
rect 25504 46452 25556 46504
rect 30840 46529 30849 46563
rect 30849 46529 30883 46563
rect 30883 46529 30892 46563
rect 30840 46520 30892 46529
rect 32128 46520 32180 46572
rect 32588 46520 32640 46572
rect 33600 46563 33652 46572
rect 33600 46529 33609 46563
rect 33609 46529 33643 46563
rect 33643 46529 33652 46563
rect 33600 46520 33652 46529
rect 34796 46563 34848 46572
rect 34796 46529 34805 46563
rect 34805 46529 34839 46563
rect 34839 46529 34848 46563
rect 34796 46520 34848 46529
rect 35808 46520 35860 46572
rect 32220 46495 32272 46504
rect 18880 46359 18932 46368
rect 18880 46325 18889 46359
rect 18889 46325 18923 46359
rect 18923 46325 18932 46359
rect 18880 46316 18932 46325
rect 19340 46359 19392 46368
rect 19340 46325 19349 46359
rect 19349 46325 19383 46359
rect 19383 46325 19392 46359
rect 19340 46316 19392 46325
rect 20996 46316 21048 46368
rect 23204 46384 23256 46436
rect 25412 46384 25464 46436
rect 32220 46461 32229 46495
rect 32229 46461 32263 46495
rect 32263 46461 32272 46495
rect 32220 46452 32272 46461
rect 33140 46452 33192 46504
rect 33876 46452 33928 46504
rect 36636 46452 36688 46504
rect 30932 46384 30984 46436
rect 31668 46384 31720 46436
rect 22376 46359 22428 46368
rect 22376 46325 22385 46359
rect 22385 46325 22419 46359
rect 22419 46325 22428 46359
rect 22376 46316 22428 46325
rect 26424 46316 26476 46368
rect 26700 46316 26752 46368
rect 27436 46359 27488 46368
rect 27436 46325 27445 46359
rect 27445 46325 27479 46359
rect 27479 46325 27488 46359
rect 27436 46316 27488 46325
rect 28264 46359 28316 46368
rect 28264 46325 28273 46359
rect 28273 46325 28307 46359
rect 28307 46325 28316 46359
rect 28264 46316 28316 46325
rect 29000 46359 29052 46368
rect 29000 46325 29009 46359
rect 29009 46325 29043 46359
rect 29043 46325 29052 46359
rect 29000 46316 29052 46325
rect 29828 46316 29880 46368
rect 32404 46316 32456 46368
rect 34796 46316 34848 46368
rect 35348 46316 35400 46368
rect 36636 46359 36688 46368
rect 36636 46325 36645 46359
rect 36645 46325 36679 46359
rect 36679 46325 36688 46359
rect 36636 46316 36688 46325
rect 37280 46359 37332 46368
rect 37280 46325 37289 46359
rect 37289 46325 37323 46359
rect 37323 46325 37332 46359
rect 37280 46316 37332 46325
rect 37832 46359 37884 46368
rect 37832 46325 37841 46359
rect 37841 46325 37875 46359
rect 37875 46325 37884 46359
rect 37832 46316 37884 46325
rect 53564 46359 53616 46368
rect 53564 46325 53573 46359
rect 53573 46325 53607 46359
rect 53607 46325 53616 46359
rect 53564 46316 53616 46325
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 19340 46112 19392 46164
rect 20996 46155 21048 46164
rect 20996 46121 21005 46155
rect 21005 46121 21039 46155
rect 21039 46121 21048 46155
rect 20996 46112 21048 46121
rect 23204 46155 23256 46164
rect 23204 46121 23213 46155
rect 23213 46121 23247 46155
rect 23247 46121 23256 46155
rect 23204 46112 23256 46121
rect 25044 46112 25096 46164
rect 29552 46155 29604 46164
rect 29552 46121 29561 46155
rect 29561 46121 29595 46155
rect 29595 46121 29604 46155
rect 29552 46112 29604 46121
rect 32404 46112 32456 46164
rect 32496 46112 32548 46164
rect 33140 46155 33192 46164
rect 33140 46121 33149 46155
rect 33149 46121 33183 46155
rect 33183 46121 33192 46155
rect 33140 46112 33192 46121
rect 32128 46044 32180 46096
rect 34244 46044 34296 46096
rect 34520 46044 34572 46096
rect 18880 45976 18932 46028
rect 19248 45976 19300 46028
rect 19984 45908 20036 45960
rect 20996 45908 21048 45960
rect 27988 46019 28040 46028
rect 22836 45908 22888 45960
rect 25136 45908 25188 45960
rect 27988 45985 27997 46019
rect 27997 45985 28031 46019
rect 28031 45985 28040 46019
rect 27988 45976 28040 45985
rect 30840 45976 30892 46028
rect 33232 46019 33284 46028
rect 33232 45985 33241 46019
rect 33241 45985 33275 46019
rect 33275 45985 33284 46019
rect 33232 45976 33284 45985
rect 33876 45976 33928 46028
rect 26332 45908 26384 45960
rect 27436 45908 27488 45960
rect 29736 45951 29788 45960
rect 29736 45917 29745 45951
rect 29745 45917 29779 45951
rect 29779 45917 29788 45951
rect 29736 45908 29788 45917
rect 29828 45951 29880 45960
rect 29828 45917 29837 45951
rect 29837 45917 29871 45951
rect 29871 45917 29880 45951
rect 29828 45908 29880 45917
rect 30196 45908 30248 45960
rect 1584 45840 1636 45892
rect 2136 45840 2188 45892
rect 21824 45840 21876 45892
rect 24400 45840 24452 45892
rect 29460 45840 29512 45892
rect 17500 45815 17552 45824
rect 17500 45781 17509 45815
rect 17509 45781 17543 45815
rect 17543 45781 17552 45815
rect 17500 45772 17552 45781
rect 20076 45772 20128 45824
rect 23020 45772 23072 45824
rect 24492 45815 24544 45824
rect 24492 45781 24501 45815
rect 24501 45781 24535 45815
rect 24535 45781 24544 45815
rect 24492 45772 24544 45781
rect 26700 45772 26752 45824
rect 28356 45772 28408 45824
rect 30932 45840 30984 45892
rect 32128 45883 32180 45892
rect 32128 45849 32137 45883
rect 32137 45849 32171 45883
rect 32171 45849 32180 45883
rect 32128 45840 32180 45849
rect 32220 45840 32272 45892
rect 34152 45951 34204 45960
rect 34152 45917 34161 45951
rect 34161 45917 34195 45951
rect 34195 45917 34204 45951
rect 34152 45908 34204 45917
rect 33416 45840 33468 45892
rect 33876 45883 33928 45892
rect 33876 45849 33885 45883
rect 33885 45849 33919 45883
rect 33919 45849 33928 45883
rect 33876 45840 33928 45849
rect 30380 45772 30432 45824
rect 31484 45815 31536 45824
rect 31484 45781 31493 45815
rect 31493 45781 31527 45815
rect 31527 45781 31536 45815
rect 31484 45772 31536 45781
rect 33324 45772 33376 45824
rect 33600 45772 33652 45824
rect 34428 45772 34480 45824
rect 34612 45908 34664 45960
rect 34980 45951 35032 45960
rect 34980 45917 34989 45951
rect 34989 45917 35023 45951
rect 35023 45917 35032 45951
rect 34980 45908 35032 45917
rect 35440 45908 35492 45960
rect 35808 45951 35860 45960
rect 35808 45917 35817 45951
rect 35817 45917 35851 45951
rect 35851 45917 35860 45951
rect 35808 45908 35860 45917
rect 37832 45908 37884 45960
rect 34612 45772 34664 45824
rect 35808 45815 35860 45824
rect 35808 45781 35817 45815
rect 35817 45781 35851 45815
rect 35851 45781 35860 45815
rect 35808 45772 35860 45781
rect 36544 45772 36596 45824
rect 37740 45772 37792 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 1584 45611 1636 45620
rect 1584 45577 1593 45611
rect 1593 45577 1627 45611
rect 1627 45577 1636 45611
rect 1584 45568 1636 45577
rect 20996 45568 21048 45620
rect 22376 45568 22428 45620
rect 24400 45568 24452 45620
rect 25136 45568 25188 45620
rect 27528 45568 27580 45620
rect 31208 45611 31260 45620
rect 31208 45577 31217 45611
rect 31217 45577 31251 45611
rect 31251 45577 31260 45611
rect 31208 45568 31260 45577
rect 32128 45568 32180 45620
rect 33600 45611 33652 45620
rect 33600 45577 33625 45611
rect 33625 45577 33652 45611
rect 33600 45568 33652 45577
rect 33876 45568 33928 45620
rect 34980 45568 35032 45620
rect 18696 45432 18748 45484
rect 19984 45475 20036 45484
rect 17776 45407 17828 45416
rect 17776 45373 17785 45407
rect 17785 45373 17819 45407
rect 17819 45373 17828 45407
rect 17776 45364 17828 45373
rect 19432 45364 19484 45416
rect 19984 45441 19993 45475
rect 19993 45441 20027 45475
rect 20027 45441 20036 45475
rect 19984 45432 20036 45441
rect 21364 45500 21416 45552
rect 25780 45543 25832 45552
rect 21456 45432 21508 45484
rect 22744 45432 22796 45484
rect 21180 45364 21232 45416
rect 22100 45364 22152 45416
rect 22376 45364 22428 45416
rect 23756 45432 23808 45484
rect 25780 45509 25789 45543
rect 25789 45509 25823 45543
rect 25823 45509 25832 45543
rect 25780 45500 25832 45509
rect 26332 45543 26384 45552
rect 26332 45509 26341 45543
rect 26341 45509 26375 45543
rect 26375 45509 26384 45543
rect 26332 45500 26384 45509
rect 28080 45500 28132 45552
rect 28908 45500 28960 45552
rect 32404 45500 32456 45552
rect 34060 45500 34112 45552
rect 34336 45500 34388 45552
rect 26700 45432 26752 45484
rect 32220 45475 32272 45484
rect 32220 45441 32229 45475
rect 32229 45441 32263 45475
rect 32263 45441 32272 45475
rect 32220 45432 32272 45441
rect 32588 45432 32640 45484
rect 37280 45500 37332 45552
rect 34612 45432 34664 45484
rect 35348 45432 35400 45484
rect 23940 45364 23992 45416
rect 26884 45364 26936 45416
rect 34336 45407 34388 45416
rect 34336 45373 34345 45407
rect 34345 45373 34379 45407
rect 34379 45373 34388 45407
rect 34336 45364 34388 45373
rect 34796 45407 34848 45416
rect 34796 45373 34805 45407
rect 34805 45373 34839 45407
rect 34839 45373 34848 45407
rect 35808 45407 35860 45416
rect 34796 45364 34848 45373
rect 35808 45373 35817 45407
rect 35817 45373 35851 45407
rect 35851 45373 35860 45407
rect 35808 45364 35860 45373
rect 19248 45296 19300 45348
rect 20720 45296 20772 45348
rect 21640 45296 21692 45348
rect 22560 45296 22612 45348
rect 27804 45296 27856 45348
rect 33140 45296 33192 45348
rect 33508 45296 33560 45348
rect 35348 45296 35400 45348
rect 18052 45228 18104 45280
rect 18880 45271 18932 45280
rect 18880 45237 18889 45271
rect 18889 45237 18923 45271
rect 18923 45237 18932 45271
rect 18880 45228 18932 45237
rect 21088 45228 21140 45280
rect 22100 45228 22152 45280
rect 23388 45228 23440 45280
rect 24216 45228 24268 45280
rect 24400 45228 24452 45280
rect 25412 45228 25464 45280
rect 27528 45228 27580 45280
rect 28356 45228 28408 45280
rect 28448 45228 28500 45280
rect 29000 45228 29052 45280
rect 30380 45228 30432 45280
rect 34520 45228 34572 45280
rect 34704 45228 34756 45280
rect 37740 45228 37792 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 16948 45024 17000 45076
rect 17316 45024 17368 45076
rect 17776 45024 17828 45076
rect 19248 45067 19300 45076
rect 19248 45033 19257 45067
rect 19257 45033 19291 45067
rect 19291 45033 19300 45067
rect 19248 45024 19300 45033
rect 19432 45024 19484 45076
rect 22560 45024 22612 45076
rect 22744 45067 22796 45076
rect 22744 45033 22753 45067
rect 22753 45033 22787 45067
rect 22787 45033 22796 45067
rect 22744 45024 22796 45033
rect 23112 45024 23164 45076
rect 27528 45024 27580 45076
rect 28264 45024 28316 45076
rect 30932 45067 30984 45076
rect 17224 44999 17276 45008
rect 17224 44965 17233 44999
rect 17233 44965 17267 44999
rect 17267 44965 17276 44999
rect 17224 44956 17276 44965
rect 19340 44956 19392 45008
rect 22928 44956 22980 45008
rect 15292 44727 15344 44736
rect 15292 44693 15301 44727
rect 15301 44693 15335 44727
rect 15335 44693 15344 44727
rect 16856 44820 16908 44872
rect 16304 44752 16356 44804
rect 17500 44820 17552 44872
rect 20904 44931 20956 44940
rect 20904 44897 20913 44931
rect 20913 44897 20947 44931
rect 20947 44897 20956 44931
rect 20904 44888 20956 44897
rect 20996 44888 21048 44940
rect 30932 45033 30941 45067
rect 30941 45033 30975 45067
rect 30975 45033 30984 45067
rect 30932 45024 30984 45033
rect 24676 44956 24728 45008
rect 23388 44931 23440 44940
rect 17132 44752 17184 44804
rect 19984 44863 20036 44872
rect 19984 44829 19993 44863
rect 19993 44829 20027 44863
rect 20027 44829 20036 44863
rect 19984 44820 20036 44829
rect 20812 44863 20864 44872
rect 20812 44829 20821 44863
rect 20821 44829 20855 44863
rect 20855 44829 20864 44863
rect 20812 44820 20864 44829
rect 21640 44863 21692 44872
rect 21640 44829 21649 44863
rect 21649 44829 21683 44863
rect 21683 44829 21692 44863
rect 21640 44820 21692 44829
rect 18328 44752 18380 44804
rect 20076 44752 20128 44804
rect 22008 44820 22060 44872
rect 23388 44897 23397 44931
rect 23397 44897 23431 44931
rect 23431 44897 23440 44931
rect 23388 44888 23440 44897
rect 22468 44820 22520 44872
rect 23756 44820 23808 44872
rect 24400 44863 24452 44872
rect 24400 44829 24409 44863
rect 24409 44829 24443 44863
rect 24443 44829 24452 44863
rect 24400 44820 24452 44829
rect 24676 44863 24728 44872
rect 24676 44829 24685 44863
rect 24685 44829 24719 44863
rect 24719 44829 24728 44863
rect 24676 44820 24728 44829
rect 25320 44956 25372 45008
rect 28908 44956 28960 45008
rect 25688 44863 25740 44872
rect 22928 44752 22980 44804
rect 25412 44795 25464 44804
rect 25412 44761 25421 44795
rect 25421 44761 25455 44795
rect 25455 44761 25464 44795
rect 25412 44752 25464 44761
rect 25688 44829 25697 44863
rect 25697 44829 25731 44863
rect 25731 44829 25740 44863
rect 25688 44820 25740 44829
rect 27712 44820 27764 44872
rect 30564 44956 30616 45008
rect 33968 45024 34020 45076
rect 34796 45024 34848 45076
rect 37280 45024 37332 45076
rect 38108 45024 38160 45076
rect 34428 44956 34480 45008
rect 30012 44888 30064 44940
rect 35348 44888 35400 44940
rect 35624 44888 35676 44940
rect 32496 44820 32548 44872
rect 32772 44863 32824 44872
rect 26424 44795 26476 44804
rect 26424 44761 26433 44795
rect 26433 44761 26467 44795
rect 26467 44761 26476 44795
rect 26424 44752 26476 44761
rect 26884 44752 26936 44804
rect 28264 44752 28316 44804
rect 32772 44829 32781 44863
rect 32781 44829 32815 44863
rect 32815 44829 32824 44863
rect 32772 44820 32824 44829
rect 33508 44820 33560 44872
rect 34152 44820 34204 44872
rect 34336 44820 34388 44872
rect 34888 44863 34940 44872
rect 34888 44829 34897 44863
rect 34897 44829 34931 44863
rect 34931 44829 34940 44863
rect 34888 44820 34940 44829
rect 35716 44863 35768 44872
rect 33324 44752 33376 44804
rect 33600 44752 33652 44804
rect 34796 44752 34848 44804
rect 35716 44829 35725 44863
rect 35725 44829 35759 44863
rect 35759 44829 35768 44863
rect 35716 44820 35768 44829
rect 36176 44863 36228 44872
rect 36176 44829 36185 44863
rect 36185 44829 36219 44863
rect 36219 44829 36228 44863
rect 36176 44820 36228 44829
rect 36544 44820 36596 44872
rect 35808 44795 35860 44804
rect 35808 44761 35817 44795
rect 35817 44761 35851 44795
rect 35851 44761 35860 44795
rect 35808 44752 35860 44761
rect 36268 44752 36320 44804
rect 15292 44684 15344 44693
rect 17592 44684 17644 44736
rect 17868 44727 17920 44736
rect 17868 44693 17877 44727
rect 17877 44693 17911 44727
rect 17911 44693 17920 44727
rect 17868 44684 17920 44693
rect 20260 44684 20312 44736
rect 20996 44684 21048 44736
rect 23020 44684 23072 44736
rect 24676 44684 24728 44736
rect 25044 44684 25096 44736
rect 27160 44727 27212 44736
rect 27160 44693 27169 44727
rect 27169 44693 27203 44727
rect 27203 44693 27212 44727
rect 27160 44684 27212 44693
rect 28172 44727 28224 44736
rect 28172 44693 28181 44727
rect 28181 44693 28215 44727
rect 28215 44693 28224 44727
rect 28172 44684 28224 44693
rect 30840 44684 30892 44736
rect 32312 44684 32364 44736
rect 33232 44727 33284 44736
rect 33232 44693 33241 44727
rect 33241 44693 33275 44727
rect 33275 44693 33284 44727
rect 33232 44684 33284 44693
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 21088 44480 21140 44532
rect 23388 44480 23440 44532
rect 27160 44480 27212 44532
rect 30840 44523 30892 44532
rect 30840 44489 30849 44523
rect 30849 44489 30883 44523
rect 30883 44489 30892 44523
rect 30840 44480 30892 44489
rect 33508 44523 33560 44532
rect 33508 44489 33517 44523
rect 33517 44489 33551 44523
rect 33551 44489 33560 44523
rect 33508 44480 33560 44489
rect 34796 44480 34848 44532
rect 34888 44480 34940 44532
rect 36176 44523 36228 44532
rect 36176 44489 36185 44523
rect 36185 44489 36219 44523
rect 36219 44489 36228 44523
rect 36176 44480 36228 44489
rect 36636 44480 36688 44532
rect 19248 44412 19300 44464
rect 20076 44455 20128 44464
rect 20076 44421 20085 44455
rect 20085 44421 20119 44455
rect 20119 44421 20128 44455
rect 20076 44412 20128 44421
rect 20260 44455 20312 44464
rect 20260 44421 20269 44455
rect 20269 44421 20303 44455
rect 20303 44421 20312 44455
rect 20260 44412 20312 44421
rect 21456 44412 21508 44464
rect 21824 44455 21876 44464
rect 21824 44421 21833 44455
rect 21833 44421 21867 44455
rect 21867 44421 21876 44455
rect 21824 44412 21876 44421
rect 23572 44412 23624 44464
rect 15108 44344 15160 44396
rect 15752 44387 15804 44396
rect 15752 44353 15761 44387
rect 15761 44353 15795 44387
rect 15795 44353 15804 44387
rect 15752 44344 15804 44353
rect 16948 44344 17000 44396
rect 17132 44344 17184 44396
rect 17500 44387 17552 44396
rect 17500 44353 17509 44387
rect 17509 44353 17543 44387
rect 17543 44353 17552 44387
rect 17500 44344 17552 44353
rect 18420 44387 18472 44396
rect 18420 44353 18429 44387
rect 18429 44353 18463 44387
rect 18463 44353 18472 44387
rect 18420 44344 18472 44353
rect 18512 44387 18564 44396
rect 18512 44353 18521 44387
rect 18521 44353 18555 44387
rect 18555 44353 18564 44387
rect 18512 44344 18564 44353
rect 21364 44344 21416 44396
rect 22284 44344 22336 44396
rect 22836 44387 22888 44396
rect 22836 44353 22845 44387
rect 22845 44353 22879 44387
rect 22879 44353 22888 44387
rect 22836 44344 22888 44353
rect 23480 44387 23532 44396
rect 23480 44353 23489 44387
rect 23489 44353 23523 44387
rect 23523 44353 23532 44387
rect 23480 44344 23532 44353
rect 23848 44344 23900 44396
rect 25412 44412 25464 44464
rect 25504 44387 25556 44396
rect 25504 44353 25513 44387
rect 25513 44353 25547 44387
rect 25547 44353 25556 44387
rect 25504 44344 25556 44353
rect 25596 44387 25648 44396
rect 25596 44353 25605 44387
rect 25605 44353 25639 44387
rect 25639 44353 25648 44387
rect 27988 44412 28040 44464
rect 28632 44455 28684 44464
rect 28632 44421 28641 44455
rect 28641 44421 28675 44455
rect 28675 44421 28684 44455
rect 28632 44412 28684 44421
rect 30932 44412 30984 44464
rect 32404 44412 32456 44464
rect 25596 44344 25648 44353
rect 18052 44276 18104 44328
rect 18604 44276 18656 44328
rect 18880 44276 18932 44328
rect 22100 44276 22152 44328
rect 22468 44276 22520 44328
rect 24216 44319 24268 44328
rect 24216 44285 24225 44319
rect 24225 44285 24259 44319
rect 24259 44285 24268 44319
rect 24216 44276 24268 44285
rect 26792 44344 26844 44396
rect 27528 44344 27580 44396
rect 30380 44387 30432 44396
rect 30380 44353 30389 44387
rect 30389 44353 30423 44387
rect 30423 44353 30432 44387
rect 30380 44344 30432 44353
rect 28080 44276 28132 44328
rect 17040 44208 17092 44260
rect 18696 44251 18748 44260
rect 18696 44217 18705 44251
rect 18705 44217 18739 44251
rect 18739 44217 18748 44251
rect 18696 44208 18748 44217
rect 21180 44208 21232 44260
rect 26148 44208 26200 44260
rect 31300 44387 31352 44396
rect 31300 44353 31309 44387
rect 31309 44353 31343 44387
rect 31343 44353 31352 44387
rect 31300 44344 31352 44353
rect 32312 44387 32364 44396
rect 32312 44353 32321 44387
rect 32321 44353 32355 44387
rect 32355 44353 32364 44387
rect 32312 44344 32364 44353
rect 32588 44344 32640 44396
rect 33048 44387 33100 44396
rect 33048 44353 33057 44387
rect 33057 44353 33091 44387
rect 33091 44353 33100 44387
rect 33048 44344 33100 44353
rect 33140 44319 33192 44328
rect 33140 44285 33149 44319
rect 33149 44285 33183 44319
rect 33183 44285 33192 44319
rect 34428 44387 34480 44396
rect 34428 44353 34437 44387
rect 34437 44353 34471 44387
rect 34471 44353 34480 44387
rect 34428 44344 34480 44353
rect 36268 44344 36320 44396
rect 36544 44387 36596 44396
rect 36544 44353 36553 44387
rect 36553 44353 36587 44387
rect 36587 44353 36596 44387
rect 36544 44344 36596 44353
rect 35716 44319 35768 44328
rect 33140 44276 33192 44285
rect 32956 44208 33008 44260
rect 33416 44208 33468 44260
rect 34152 44251 34204 44260
rect 34152 44217 34161 44251
rect 34161 44217 34195 44251
rect 34195 44217 34204 44251
rect 34152 44208 34204 44217
rect 35716 44285 35725 44319
rect 35725 44285 35759 44319
rect 35759 44285 35768 44319
rect 35716 44276 35768 44285
rect 1676 44140 1728 44192
rect 14096 44140 14148 44192
rect 14464 44183 14516 44192
rect 14464 44149 14473 44183
rect 14473 44149 14507 44183
rect 14507 44149 14516 44183
rect 14464 44140 14516 44149
rect 15016 44183 15068 44192
rect 15016 44149 15025 44183
rect 15025 44149 15059 44183
rect 15059 44149 15068 44183
rect 15016 44140 15068 44149
rect 17132 44140 17184 44192
rect 17684 44183 17736 44192
rect 17684 44149 17693 44183
rect 17693 44149 17727 44183
rect 17727 44149 17736 44183
rect 17684 44140 17736 44149
rect 18512 44140 18564 44192
rect 20812 44140 20864 44192
rect 25044 44140 25096 44192
rect 26240 44140 26292 44192
rect 31300 44140 31352 44192
rect 31576 44140 31628 44192
rect 34796 44140 34848 44192
rect 36728 44208 36780 44260
rect 38384 44251 38436 44260
rect 38384 44217 38393 44251
rect 38393 44217 38427 44251
rect 38427 44217 38436 44251
rect 38384 44208 38436 44217
rect 35716 44140 35768 44192
rect 39120 44140 39172 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 10692 43936 10744 43988
rect 15292 43936 15344 43988
rect 18420 43979 18472 43988
rect 16856 43868 16908 43920
rect 1584 43664 1636 43716
rect 14464 43800 14516 43852
rect 14740 43775 14792 43784
rect 14740 43741 14749 43775
rect 14749 43741 14783 43775
rect 14783 43741 14792 43775
rect 14740 43732 14792 43741
rect 14924 43775 14976 43784
rect 14924 43741 14933 43775
rect 14933 43741 14967 43775
rect 14967 43741 14976 43775
rect 14924 43732 14976 43741
rect 15292 43732 15344 43784
rect 16304 43800 16356 43852
rect 17500 43868 17552 43920
rect 18420 43945 18429 43979
rect 18429 43945 18463 43979
rect 18463 43945 18472 43979
rect 18420 43936 18472 43945
rect 18604 43936 18656 43988
rect 19984 43868 20036 43920
rect 20352 43868 20404 43920
rect 20904 43936 20956 43988
rect 23756 43936 23808 43988
rect 24584 43936 24636 43988
rect 25688 43936 25740 43988
rect 17224 43843 17276 43852
rect 17224 43809 17233 43843
rect 17233 43809 17267 43843
rect 17267 43809 17276 43843
rect 17224 43800 17276 43809
rect 17684 43800 17736 43852
rect 23940 43868 23992 43920
rect 29000 43936 29052 43988
rect 32772 43936 32824 43988
rect 33416 43979 33468 43988
rect 17040 43732 17092 43784
rect 17592 43732 17644 43784
rect 22284 43800 22336 43852
rect 16304 43707 16356 43716
rect 16304 43673 16313 43707
rect 16313 43673 16347 43707
rect 16347 43673 16356 43707
rect 16304 43664 16356 43673
rect 17868 43664 17920 43716
rect 19432 43732 19484 43784
rect 20076 43732 20128 43784
rect 20720 43775 20772 43784
rect 20720 43741 20729 43775
rect 20729 43741 20763 43775
rect 20763 43741 20772 43775
rect 20720 43732 20772 43741
rect 21180 43775 21232 43784
rect 21180 43741 21189 43775
rect 21189 43741 21223 43775
rect 21223 43741 21232 43775
rect 21180 43732 21232 43741
rect 21456 43775 21508 43784
rect 21456 43741 21465 43775
rect 21465 43741 21499 43775
rect 21499 43741 21508 43775
rect 21456 43732 21508 43741
rect 22008 43732 22060 43784
rect 22100 43775 22152 43784
rect 22100 43741 22109 43775
rect 22109 43741 22143 43775
rect 22143 43741 22152 43775
rect 22100 43732 22152 43741
rect 22836 43732 22888 43784
rect 23572 43775 23624 43784
rect 23572 43741 23581 43775
rect 23581 43741 23615 43775
rect 23615 43741 23624 43775
rect 23572 43732 23624 43741
rect 24032 43800 24084 43852
rect 25044 43843 25096 43852
rect 25044 43809 25053 43843
rect 25053 43809 25087 43843
rect 25087 43809 25096 43843
rect 25044 43800 25096 43809
rect 26148 43868 26200 43920
rect 25320 43775 25372 43784
rect 25320 43741 25329 43775
rect 25329 43741 25363 43775
rect 25363 43741 25372 43775
rect 25320 43732 25372 43741
rect 25780 43732 25832 43784
rect 28632 43800 28684 43852
rect 33416 43945 33425 43979
rect 33425 43945 33459 43979
rect 33459 43945 33468 43979
rect 33416 43936 33468 43945
rect 34796 43936 34848 43988
rect 36544 43936 36596 43988
rect 36268 43868 36320 43920
rect 37832 43868 37884 43920
rect 33048 43800 33100 43852
rect 34796 43800 34848 43852
rect 35900 43843 35952 43852
rect 35900 43809 35909 43843
rect 35909 43809 35943 43843
rect 35943 43809 35952 43843
rect 35900 43800 35952 43809
rect 18604 43664 18656 43716
rect 14464 43596 14516 43648
rect 15384 43596 15436 43648
rect 17408 43596 17460 43648
rect 17776 43596 17828 43648
rect 19340 43596 19392 43648
rect 19984 43664 20036 43716
rect 21088 43664 21140 43716
rect 23480 43664 23532 43716
rect 23848 43707 23900 43716
rect 23848 43673 23857 43707
rect 23857 43673 23891 43707
rect 23891 43673 23900 43707
rect 23848 43664 23900 43673
rect 24032 43664 24084 43716
rect 25596 43664 25648 43716
rect 20076 43596 20128 43648
rect 21364 43639 21416 43648
rect 21364 43605 21373 43639
rect 21373 43605 21407 43639
rect 21407 43605 21416 43639
rect 21364 43596 21416 43605
rect 23572 43596 23624 43648
rect 24400 43639 24452 43648
rect 24400 43605 24409 43639
rect 24409 43605 24443 43639
rect 24443 43605 24452 43639
rect 24400 43596 24452 43605
rect 28908 43732 28960 43784
rect 30104 43732 30156 43784
rect 30932 43732 30984 43784
rect 33232 43732 33284 43784
rect 33600 43775 33652 43784
rect 33600 43741 33609 43775
rect 33609 43741 33643 43775
rect 33643 43741 33652 43775
rect 33600 43732 33652 43741
rect 36268 43732 36320 43784
rect 36452 43732 36504 43784
rect 28264 43596 28316 43648
rect 30748 43596 30800 43648
rect 32680 43664 32732 43716
rect 31484 43596 31536 43648
rect 36728 43596 36780 43648
rect 38660 43596 38712 43648
rect 39120 43639 39172 43648
rect 39120 43605 39129 43639
rect 39129 43605 39163 43639
rect 39163 43605 39172 43639
rect 39120 43596 39172 43605
rect 52368 43596 52420 43648
rect 53564 43639 53616 43648
rect 53564 43605 53573 43639
rect 53573 43605 53607 43639
rect 53607 43605 53616 43639
rect 53564 43596 53616 43605
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 1584 43435 1636 43444
rect 1584 43401 1593 43435
rect 1593 43401 1627 43435
rect 1627 43401 1636 43435
rect 1584 43392 1636 43401
rect 14924 43435 14976 43444
rect 14924 43401 14933 43435
rect 14933 43401 14967 43435
rect 14967 43401 14976 43435
rect 14924 43392 14976 43401
rect 16948 43392 17000 43444
rect 17592 43392 17644 43444
rect 18512 43435 18564 43444
rect 18512 43401 18521 43435
rect 18521 43401 18555 43435
rect 18555 43401 18564 43435
rect 18512 43392 18564 43401
rect 19340 43392 19392 43444
rect 14096 43367 14148 43376
rect 14096 43333 14105 43367
rect 14105 43333 14139 43367
rect 14139 43333 14148 43367
rect 14096 43324 14148 43333
rect 14280 43299 14332 43308
rect 14280 43265 14289 43299
rect 14289 43265 14323 43299
rect 14323 43265 14332 43299
rect 14280 43256 14332 43265
rect 14740 43256 14792 43308
rect 16856 43299 16908 43308
rect 16856 43265 16865 43299
rect 16865 43265 16899 43299
rect 16899 43265 16908 43299
rect 16856 43256 16908 43265
rect 17316 43324 17368 43376
rect 17040 43256 17092 43308
rect 17224 43299 17276 43308
rect 17224 43265 17233 43299
rect 17233 43265 17267 43299
rect 17267 43265 17276 43299
rect 17684 43324 17736 43376
rect 17224 43256 17276 43265
rect 17960 43256 18012 43308
rect 18604 43299 18656 43308
rect 18604 43265 18613 43299
rect 18613 43265 18647 43299
rect 18647 43265 18656 43299
rect 19984 43324 20036 43376
rect 20812 43367 20864 43376
rect 20812 43333 20821 43367
rect 20821 43333 20855 43367
rect 20855 43333 20864 43367
rect 20812 43324 20864 43333
rect 18604 43256 18656 43265
rect 15752 43188 15804 43240
rect 16764 43120 16816 43172
rect 16672 43095 16724 43104
rect 16672 43061 16681 43095
rect 16681 43061 16715 43095
rect 16715 43061 16724 43095
rect 16672 43052 16724 43061
rect 17500 43188 17552 43240
rect 18052 43231 18104 43240
rect 18052 43197 18061 43231
rect 18061 43197 18095 43231
rect 18095 43197 18104 43231
rect 18052 43188 18104 43197
rect 17592 43120 17644 43172
rect 19432 43052 19484 43104
rect 22100 43299 22152 43308
rect 22100 43265 22109 43299
rect 22109 43265 22143 43299
rect 22143 43265 22152 43299
rect 22100 43256 22152 43265
rect 22376 43256 22428 43308
rect 23204 43392 23256 43444
rect 25688 43392 25740 43444
rect 27712 43435 27764 43444
rect 27712 43401 27721 43435
rect 27721 43401 27755 43435
rect 27755 43401 27764 43435
rect 27712 43392 27764 43401
rect 30104 43435 30156 43444
rect 30104 43401 30113 43435
rect 30113 43401 30147 43435
rect 30147 43401 30156 43435
rect 30104 43392 30156 43401
rect 31116 43392 31168 43444
rect 31208 43392 31260 43444
rect 32680 43392 32732 43444
rect 51632 43392 51684 43444
rect 23848 43324 23900 43376
rect 29000 43324 29052 43376
rect 30012 43324 30064 43376
rect 30840 43367 30892 43376
rect 23388 43299 23440 43308
rect 23388 43265 23397 43299
rect 23397 43265 23431 43299
rect 23431 43265 23440 43299
rect 23388 43256 23440 43265
rect 23572 43299 23624 43308
rect 23572 43265 23581 43299
rect 23581 43265 23615 43299
rect 23615 43265 23624 43299
rect 23572 43256 23624 43265
rect 23940 43256 23992 43308
rect 25320 43256 25372 43308
rect 25504 43256 25556 43308
rect 27068 43299 27120 43308
rect 27068 43265 27077 43299
rect 27077 43265 27111 43299
rect 27111 43265 27120 43299
rect 27068 43256 27120 43265
rect 24584 43231 24636 43240
rect 24584 43197 24593 43231
rect 24593 43197 24627 43231
rect 24627 43197 24636 43231
rect 24584 43188 24636 43197
rect 25044 43188 25096 43240
rect 25412 43231 25464 43240
rect 25412 43197 25421 43231
rect 25421 43197 25455 43231
rect 25455 43197 25464 43231
rect 25412 43188 25464 43197
rect 26424 43188 26476 43240
rect 28448 43256 28500 43308
rect 30380 43256 30432 43308
rect 30840 43333 30849 43367
rect 30849 43333 30883 43367
rect 30883 43333 30892 43367
rect 30840 43324 30892 43333
rect 31300 43324 31352 43376
rect 31392 43367 31444 43376
rect 31392 43333 31401 43367
rect 31401 43333 31435 43367
rect 31435 43333 31444 43367
rect 31392 43324 31444 43333
rect 32588 43324 32640 43376
rect 22376 43120 22428 43172
rect 23664 43120 23716 43172
rect 19984 43052 20036 43104
rect 21088 43052 21140 43104
rect 23204 43052 23256 43104
rect 24308 43052 24360 43104
rect 26516 43120 26568 43172
rect 28540 43188 28592 43240
rect 31208 43299 31260 43308
rect 31208 43265 31217 43299
rect 31217 43265 31251 43299
rect 31251 43265 31260 43299
rect 31208 43256 31260 43265
rect 31484 43256 31536 43308
rect 32128 43256 32180 43308
rect 33784 43299 33836 43308
rect 33784 43265 33793 43299
rect 33793 43265 33827 43299
rect 33827 43265 33836 43299
rect 33784 43256 33836 43265
rect 34244 43299 34296 43308
rect 34244 43265 34253 43299
rect 34253 43265 34287 43299
rect 34287 43265 34296 43299
rect 34244 43256 34296 43265
rect 34336 43256 34388 43308
rect 35532 43299 35584 43308
rect 35532 43265 35541 43299
rect 35541 43265 35575 43299
rect 35575 43265 35584 43299
rect 35532 43256 35584 43265
rect 35992 43324 36044 43376
rect 37188 43324 37240 43376
rect 37832 43367 37884 43376
rect 37832 43333 37841 43367
rect 37841 43333 37875 43367
rect 37875 43333 37884 43367
rect 37832 43324 37884 43333
rect 31300 43188 31352 43240
rect 33140 43188 33192 43240
rect 33968 43188 34020 43240
rect 35900 43188 35952 43240
rect 36268 43299 36320 43308
rect 36268 43265 36277 43299
rect 36277 43265 36311 43299
rect 36311 43265 36320 43299
rect 36268 43256 36320 43265
rect 37372 43256 37424 43308
rect 37188 43188 37240 43240
rect 33692 43163 33744 43172
rect 25044 43052 25096 43104
rect 27252 43052 27304 43104
rect 27344 43052 27396 43104
rect 33692 43129 33701 43163
rect 33701 43129 33735 43163
rect 33735 43129 33744 43163
rect 33692 43120 33744 43129
rect 33876 43120 33928 43172
rect 39948 43120 40000 43172
rect 29828 43052 29880 43104
rect 32404 43052 32456 43104
rect 33232 43052 33284 43104
rect 36176 43052 36228 43104
rect 36360 43052 36412 43104
rect 38384 43052 38436 43104
rect 39488 43095 39540 43104
rect 39488 43061 39497 43095
rect 39497 43061 39531 43095
rect 39531 43061 39540 43095
rect 39488 43052 39540 43061
rect 40500 43052 40552 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 14096 42848 14148 42900
rect 14740 42848 14792 42900
rect 16856 42848 16908 42900
rect 17684 42891 17736 42900
rect 17684 42857 17693 42891
rect 17693 42857 17727 42891
rect 17727 42857 17736 42891
rect 17684 42848 17736 42857
rect 18328 42848 18380 42900
rect 27068 42848 27120 42900
rect 28264 42848 28316 42900
rect 15108 42755 15160 42764
rect 15108 42721 15117 42755
rect 15117 42721 15151 42755
rect 15151 42721 15160 42755
rect 15108 42712 15160 42721
rect 14096 42687 14148 42696
rect 14096 42653 14105 42687
rect 14105 42653 14139 42687
rect 14139 42653 14148 42687
rect 14096 42644 14148 42653
rect 14280 42687 14332 42696
rect 14280 42653 14289 42687
rect 14289 42653 14323 42687
rect 14323 42653 14332 42687
rect 16672 42712 16724 42764
rect 17132 42712 17184 42764
rect 14280 42644 14332 42653
rect 16764 42687 16816 42696
rect 13636 42576 13688 42628
rect 14924 42619 14976 42628
rect 14924 42585 14933 42619
rect 14933 42585 14967 42619
rect 14967 42585 14976 42619
rect 14924 42576 14976 42585
rect 15384 42576 15436 42628
rect 16764 42653 16773 42687
rect 16773 42653 16807 42687
rect 16807 42653 16816 42687
rect 16764 42644 16816 42653
rect 17224 42644 17276 42696
rect 18972 42712 19024 42764
rect 24032 42780 24084 42832
rect 27252 42823 27304 42832
rect 27252 42789 27261 42823
rect 27261 42789 27295 42823
rect 27295 42789 27304 42823
rect 27252 42780 27304 42789
rect 27528 42780 27580 42832
rect 28080 42780 28132 42832
rect 17776 42687 17828 42696
rect 17776 42653 17785 42687
rect 17785 42653 17819 42687
rect 17819 42653 17828 42687
rect 17776 42644 17828 42653
rect 20076 42644 20128 42696
rect 20352 42687 20404 42696
rect 20352 42653 20361 42687
rect 20361 42653 20395 42687
rect 20395 42653 20404 42687
rect 20352 42644 20404 42653
rect 17592 42576 17644 42628
rect 20260 42619 20312 42628
rect 20260 42585 20269 42619
rect 20269 42585 20303 42619
rect 20303 42585 20312 42619
rect 20260 42576 20312 42585
rect 2872 42508 2924 42560
rect 15752 42508 15804 42560
rect 17316 42508 17368 42560
rect 18052 42551 18104 42560
rect 18052 42517 18061 42551
rect 18061 42517 18095 42551
rect 18095 42517 18104 42551
rect 18052 42508 18104 42517
rect 20168 42551 20220 42560
rect 20168 42517 20177 42551
rect 20177 42517 20211 42551
rect 20211 42517 20220 42551
rect 20168 42508 20220 42517
rect 22008 42712 22060 42764
rect 22100 42712 22152 42764
rect 23664 42712 23716 42764
rect 25320 42755 25372 42764
rect 25320 42721 25329 42755
rect 25329 42721 25363 42755
rect 25363 42721 25372 42755
rect 25320 42712 25372 42721
rect 23112 42687 23164 42696
rect 23112 42653 23121 42687
rect 23121 42653 23155 42687
rect 23155 42653 23164 42687
rect 23112 42644 23164 42653
rect 23480 42644 23532 42696
rect 24492 42644 24544 42696
rect 25412 42687 25464 42696
rect 25412 42653 25421 42687
rect 25421 42653 25455 42687
rect 25455 42653 25464 42687
rect 25412 42644 25464 42653
rect 26792 42687 26844 42696
rect 26792 42653 26801 42687
rect 26801 42653 26835 42687
rect 26835 42653 26844 42687
rect 26792 42644 26844 42653
rect 27252 42644 27304 42696
rect 29552 42712 29604 42764
rect 31116 42848 31168 42900
rect 32128 42891 32180 42900
rect 32128 42857 32137 42891
rect 32137 42857 32171 42891
rect 32171 42857 32180 42891
rect 32128 42848 32180 42857
rect 35532 42891 35584 42900
rect 30472 42780 30524 42832
rect 34060 42823 34112 42832
rect 31392 42712 31444 42764
rect 27436 42644 27488 42696
rect 24216 42508 24268 42560
rect 28908 42576 28960 42628
rect 30012 42687 30064 42696
rect 30012 42653 30021 42687
rect 30021 42653 30055 42687
rect 30055 42653 30064 42687
rect 34060 42789 34069 42823
rect 34069 42789 34103 42823
rect 34103 42789 34112 42823
rect 34060 42780 34112 42789
rect 33600 42712 33652 42764
rect 34336 42712 34388 42764
rect 35532 42857 35541 42891
rect 35541 42857 35575 42891
rect 35575 42857 35584 42891
rect 35532 42848 35584 42857
rect 35992 42891 36044 42900
rect 35992 42857 36001 42891
rect 36001 42857 36035 42891
rect 36035 42857 36044 42891
rect 35992 42848 36044 42857
rect 36452 42848 36504 42900
rect 36268 42780 36320 42832
rect 37464 42780 37516 42832
rect 39488 42780 39540 42832
rect 30012 42644 30064 42653
rect 30840 42576 30892 42628
rect 31024 42576 31076 42628
rect 33048 42687 33100 42696
rect 33048 42653 33057 42687
rect 33057 42653 33091 42687
rect 33091 42653 33100 42687
rect 33048 42644 33100 42653
rect 33692 42644 33744 42696
rect 34244 42644 34296 42696
rect 36728 42712 36780 42764
rect 36820 42712 36872 42764
rect 34796 42644 34848 42696
rect 35348 42687 35400 42696
rect 35348 42653 35357 42687
rect 35357 42653 35391 42687
rect 35391 42653 35400 42687
rect 35348 42644 35400 42653
rect 35532 42687 35584 42696
rect 35532 42653 35541 42687
rect 35541 42653 35575 42687
rect 35575 42653 35584 42687
rect 35532 42644 35584 42653
rect 36452 42644 36504 42696
rect 37004 42689 37056 42696
rect 37004 42655 37013 42689
rect 37013 42655 37047 42689
rect 37047 42655 37056 42689
rect 37004 42644 37056 42655
rect 34980 42576 35032 42628
rect 38660 42712 38712 42764
rect 40040 42712 40092 42764
rect 38936 42644 38988 42696
rect 39120 42576 39172 42628
rect 26240 42551 26292 42560
rect 26240 42517 26249 42551
rect 26249 42517 26283 42551
rect 26283 42517 26292 42551
rect 26240 42508 26292 42517
rect 27712 42508 27764 42560
rect 28172 42508 28224 42560
rect 29644 42508 29696 42560
rect 30564 42551 30616 42560
rect 30564 42517 30573 42551
rect 30573 42517 30607 42551
rect 30607 42517 30616 42551
rect 30564 42508 30616 42517
rect 33600 42508 33652 42560
rect 33968 42508 34020 42560
rect 37464 42508 37516 42560
rect 38384 42508 38436 42560
rect 39948 42551 40000 42560
rect 39948 42517 39957 42551
rect 39957 42517 39991 42551
rect 39991 42517 40000 42551
rect 39948 42508 40000 42517
rect 40960 42551 41012 42560
rect 40960 42517 40969 42551
rect 40969 42517 41003 42551
rect 41003 42517 41012 42551
rect 40960 42508 41012 42517
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 15752 42304 15804 42356
rect 15384 42236 15436 42288
rect 13636 42168 13688 42220
rect 14924 42211 14976 42220
rect 14924 42177 14933 42211
rect 14933 42177 14967 42211
rect 14967 42177 14976 42211
rect 14924 42168 14976 42177
rect 16672 42304 16724 42356
rect 17132 42304 17184 42356
rect 17776 42304 17828 42356
rect 20260 42304 20312 42356
rect 20444 42304 20496 42356
rect 22376 42347 22428 42356
rect 22376 42313 22385 42347
rect 22385 42313 22419 42347
rect 22419 42313 22428 42347
rect 22376 42304 22428 42313
rect 23848 42304 23900 42356
rect 25412 42304 25464 42356
rect 25780 42304 25832 42356
rect 26332 42347 26384 42356
rect 26332 42313 26341 42347
rect 26341 42313 26375 42347
rect 26375 42313 26384 42347
rect 26332 42304 26384 42313
rect 27344 42304 27396 42356
rect 28908 42304 28960 42356
rect 29552 42347 29604 42356
rect 29552 42313 29561 42347
rect 29561 42313 29595 42347
rect 29595 42313 29604 42347
rect 29552 42304 29604 42313
rect 30564 42304 30616 42356
rect 30840 42304 30892 42356
rect 31208 42304 31260 42356
rect 31484 42304 31536 42356
rect 34980 42347 35032 42356
rect 34980 42313 34989 42347
rect 34989 42313 35023 42347
rect 35023 42313 35032 42347
rect 34980 42304 35032 42313
rect 35808 42304 35860 42356
rect 16212 42236 16264 42288
rect 18880 42236 18932 42288
rect 19432 42236 19484 42288
rect 17040 42168 17092 42220
rect 17408 42168 17460 42220
rect 17868 42168 17920 42220
rect 20076 42168 20128 42220
rect 20444 42211 20496 42220
rect 20444 42177 20453 42211
rect 20453 42177 20487 42211
rect 20487 42177 20496 42211
rect 20444 42168 20496 42177
rect 20720 42211 20772 42220
rect 20720 42177 20729 42211
rect 20729 42177 20763 42211
rect 20763 42177 20772 42211
rect 20720 42168 20772 42177
rect 21824 42236 21876 42288
rect 23296 42236 23348 42288
rect 23204 42211 23256 42220
rect 19984 42100 20036 42152
rect 23204 42177 23213 42211
rect 23213 42177 23247 42211
rect 23247 42177 23256 42211
rect 23204 42168 23256 42177
rect 23388 42211 23440 42220
rect 23388 42177 23397 42211
rect 23397 42177 23431 42211
rect 23431 42177 23440 42211
rect 23388 42168 23440 42177
rect 24216 42168 24268 42220
rect 24492 42168 24544 42220
rect 27712 42236 27764 42288
rect 27344 42211 27396 42220
rect 27344 42177 27353 42211
rect 27353 42177 27387 42211
rect 27387 42177 27396 42211
rect 27344 42168 27396 42177
rect 27528 42168 27580 42220
rect 23112 42100 23164 42152
rect 26240 42100 26292 42152
rect 28908 42211 28960 42220
rect 28908 42177 28917 42211
rect 28917 42177 28951 42211
rect 28951 42177 28960 42211
rect 28908 42168 28960 42177
rect 30748 42236 30800 42288
rect 33784 42236 33836 42288
rect 35348 42279 35400 42288
rect 30656 42211 30708 42220
rect 30656 42177 30674 42211
rect 30674 42177 30708 42211
rect 30656 42168 30708 42177
rect 30932 42211 30984 42220
rect 30932 42177 30941 42211
rect 30941 42177 30975 42211
rect 30975 42177 30984 42211
rect 30932 42168 30984 42177
rect 32128 42211 32180 42220
rect 32128 42177 32137 42211
rect 32137 42177 32171 42211
rect 32171 42177 32180 42211
rect 32128 42168 32180 42177
rect 34060 42211 34112 42220
rect 33232 42143 33284 42152
rect 16028 42032 16080 42084
rect 17684 42032 17736 42084
rect 13636 42007 13688 42016
rect 13636 41973 13645 42007
rect 13645 41973 13679 42007
rect 13679 41973 13688 42007
rect 13636 41964 13688 41973
rect 14280 41964 14332 42016
rect 18512 41964 18564 42016
rect 20444 41964 20496 42016
rect 21364 42032 21416 42084
rect 26792 42032 26844 42084
rect 22008 41964 22060 42016
rect 27896 41964 27948 42016
rect 33232 42109 33241 42143
rect 33241 42109 33275 42143
rect 33275 42109 33284 42143
rect 33232 42100 33284 42109
rect 34060 42177 34069 42211
rect 34069 42177 34103 42211
rect 34103 42177 34112 42211
rect 34060 42168 34112 42177
rect 35348 42245 35357 42279
rect 35357 42245 35391 42279
rect 35391 42245 35400 42279
rect 35348 42236 35400 42245
rect 34612 42100 34664 42152
rect 35900 42211 35952 42220
rect 35900 42177 35909 42211
rect 35909 42177 35943 42211
rect 35943 42177 35952 42211
rect 35900 42168 35952 42177
rect 35992 42168 36044 42220
rect 36820 42236 36872 42288
rect 37372 42279 37424 42288
rect 37372 42245 37381 42279
rect 37381 42245 37415 42279
rect 37415 42245 37424 42279
rect 37372 42236 37424 42245
rect 38384 42304 38436 42356
rect 40500 42347 40552 42356
rect 28540 42032 28592 42084
rect 33600 42032 33652 42084
rect 33876 42032 33928 42084
rect 35532 42032 35584 42084
rect 37188 42168 37240 42220
rect 38016 42236 38068 42288
rect 40500 42313 40509 42347
rect 40509 42313 40543 42347
rect 40543 42313 40552 42347
rect 40500 42304 40552 42313
rect 37832 42168 37884 42220
rect 38108 42100 38160 42152
rect 37372 42032 37424 42084
rect 32404 41964 32456 42016
rect 34336 41964 34388 42016
rect 34796 41964 34848 42016
rect 37556 41964 37608 42016
rect 39028 41964 39080 42016
rect 40960 41964 41012 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 13636 41760 13688 41812
rect 16948 41760 17000 41812
rect 17592 41803 17644 41812
rect 17592 41769 17601 41803
rect 17601 41769 17635 41803
rect 17635 41769 17644 41803
rect 17592 41760 17644 41769
rect 18328 41760 18380 41812
rect 24492 41760 24544 41812
rect 21640 41692 21692 41744
rect 20168 41624 20220 41676
rect 28448 41760 28500 41812
rect 30380 41803 30432 41812
rect 30380 41769 30389 41803
rect 30389 41769 30423 41803
rect 30423 41769 30432 41803
rect 30380 41760 30432 41769
rect 33692 41760 33744 41812
rect 34152 41760 34204 41812
rect 35716 41760 35768 41812
rect 38936 41803 38988 41812
rect 38936 41769 38945 41803
rect 38945 41769 38979 41803
rect 38979 41769 38988 41803
rect 38936 41760 38988 41769
rect 40040 41760 40092 41812
rect 40408 41760 40460 41812
rect 40960 41760 41012 41812
rect 27436 41692 27488 41744
rect 17776 41599 17828 41608
rect 17776 41565 17785 41599
rect 17785 41565 17819 41599
rect 17819 41565 17828 41599
rect 17776 41556 17828 41565
rect 17960 41599 18012 41608
rect 17960 41565 17969 41599
rect 17969 41565 18003 41599
rect 18003 41565 18012 41599
rect 17960 41556 18012 41565
rect 18236 41556 18288 41608
rect 20260 41599 20312 41608
rect 20260 41565 20269 41599
rect 20269 41565 20303 41599
rect 20303 41565 20312 41599
rect 20260 41556 20312 41565
rect 20444 41599 20496 41608
rect 20444 41565 20453 41599
rect 20453 41565 20487 41599
rect 20487 41565 20496 41599
rect 20444 41556 20496 41565
rect 20996 41599 21048 41608
rect 17132 41531 17184 41540
rect 17132 41497 17141 41531
rect 17141 41497 17175 41531
rect 17175 41497 17184 41531
rect 17132 41488 17184 41497
rect 19432 41488 19484 41540
rect 20352 41488 20404 41540
rect 20996 41565 21005 41599
rect 21005 41565 21039 41599
rect 21039 41565 21048 41599
rect 20996 41556 21048 41565
rect 21180 41599 21232 41608
rect 21180 41565 21189 41599
rect 21189 41565 21223 41599
rect 21223 41565 21232 41599
rect 21824 41599 21876 41608
rect 21180 41556 21232 41565
rect 21824 41565 21833 41599
rect 21833 41565 21867 41599
rect 21867 41565 21876 41599
rect 21824 41556 21876 41565
rect 22744 41556 22796 41608
rect 23296 41556 23348 41608
rect 25320 41556 25372 41608
rect 25504 41599 25556 41608
rect 25504 41565 25513 41599
rect 25513 41565 25547 41599
rect 25547 41565 25556 41599
rect 25504 41556 25556 41565
rect 25596 41556 25648 41608
rect 23848 41488 23900 41540
rect 24676 41531 24728 41540
rect 24676 41497 24685 41531
rect 24685 41497 24719 41531
rect 24719 41497 24728 41531
rect 24676 41488 24728 41497
rect 27712 41556 27764 41608
rect 37188 41692 37240 41744
rect 27896 41624 27948 41676
rect 30932 41624 30984 41676
rect 34428 41624 34480 41676
rect 36360 41667 36412 41676
rect 31576 41556 31628 41608
rect 32404 41599 32456 41608
rect 32404 41565 32438 41599
rect 32438 41565 32456 41599
rect 32404 41556 32456 41565
rect 34152 41556 34204 41608
rect 36360 41633 36369 41667
rect 36369 41633 36403 41667
rect 36403 41633 36412 41667
rect 36360 41624 36412 41633
rect 37004 41624 37056 41676
rect 35992 41556 36044 41608
rect 29000 41531 29052 41540
rect 29000 41497 29009 41531
rect 29009 41497 29043 41531
rect 29043 41497 29052 41531
rect 29000 41488 29052 41497
rect 30288 41488 30340 41540
rect 32220 41488 32272 41540
rect 34244 41488 34296 41540
rect 36268 41488 36320 41540
rect 38108 41556 38160 41608
rect 40040 41624 40092 41676
rect 39028 41556 39080 41608
rect 39120 41599 39172 41608
rect 39120 41565 39129 41599
rect 39129 41565 39163 41599
rect 39163 41565 39172 41599
rect 39120 41556 39172 41565
rect 37464 41531 37516 41540
rect 37464 41497 37473 41531
rect 37473 41497 37507 41531
rect 37507 41497 37516 41531
rect 37464 41488 37516 41497
rect 16028 41463 16080 41472
rect 16028 41429 16037 41463
rect 16037 41429 16071 41463
rect 16071 41429 16080 41463
rect 16028 41420 16080 41429
rect 19340 41420 19392 41472
rect 20628 41420 20680 41472
rect 26608 41420 26660 41472
rect 26884 41420 26936 41472
rect 27068 41420 27120 41472
rect 33876 41420 33928 41472
rect 33968 41420 34020 41472
rect 34428 41420 34480 41472
rect 35348 41420 35400 41472
rect 35808 41420 35860 41472
rect 36360 41420 36412 41472
rect 36728 41420 36780 41472
rect 37372 41463 37424 41472
rect 37372 41429 37381 41463
rect 37381 41429 37415 41463
rect 37415 41429 37424 41463
rect 37372 41420 37424 41429
rect 38200 41420 38252 41472
rect 53380 41531 53432 41540
rect 53380 41497 53389 41531
rect 53389 41497 53423 41531
rect 53423 41497 53432 41531
rect 53380 41488 53432 41497
rect 53564 41531 53616 41540
rect 53564 41497 53573 41531
rect 53573 41497 53607 41531
rect 53607 41497 53616 41531
rect 53564 41488 53616 41497
rect 42064 41463 42116 41472
rect 42064 41429 42073 41463
rect 42073 41429 42107 41463
rect 42107 41429 42116 41463
rect 42064 41420 42116 41429
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 16028 41259 16080 41268
rect 16028 41225 16037 41259
rect 16037 41225 16071 41259
rect 16071 41225 16080 41259
rect 16028 41216 16080 41225
rect 17960 41216 18012 41268
rect 18144 41216 18196 41268
rect 25504 41216 25556 41268
rect 26884 41216 26936 41268
rect 18052 41148 18104 41200
rect 26056 41148 26108 41200
rect 26332 41148 26384 41200
rect 26516 41148 26568 41200
rect 28172 41216 28224 41268
rect 30656 41216 30708 41268
rect 32128 41216 32180 41268
rect 34428 41216 34480 41268
rect 36636 41259 36688 41268
rect 36636 41225 36645 41259
rect 36645 41225 36679 41259
rect 36679 41225 36688 41259
rect 36636 41216 36688 41225
rect 37188 41216 37240 41268
rect 38016 41259 38068 41268
rect 38016 41225 38025 41259
rect 38025 41225 38059 41259
rect 38059 41225 38068 41259
rect 38016 41216 38068 41225
rect 29920 41148 29972 41200
rect 32680 41148 32732 41200
rect 33600 41191 33652 41200
rect 33600 41157 33635 41191
rect 33635 41157 33652 41191
rect 33600 41148 33652 41157
rect 33784 41148 33836 41200
rect 38660 41216 38712 41268
rect 41052 41216 41104 41268
rect 18236 41080 18288 41132
rect 18604 41123 18656 41132
rect 18604 41089 18613 41123
rect 18613 41089 18647 41123
rect 18647 41089 18656 41123
rect 18604 41080 18656 41089
rect 19432 41080 19484 41132
rect 17592 41012 17644 41064
rect 16948 40944 17000 40996
rect 1492 40919 1544 40928
rect 1492 40885 1501 40919
rect 1501 40885 1535 40919
rect 1535 40885 1544 40919
rect 1492 40876 1544 40885
rect 16672 40876 16724 40928
rect 17960 40944 18012 40996
rect 18788 40987 18840 40996
rect 18788 40953 18797 40987
rect 18797 40953 18831 40987
rect 18831 40953 18840 40987
rect 18788 40944 18840 40953
rect 20720 41080 20772 41132
rect 21272 41123 21324 41132
rect 21272 41089 21281 41123
rect 21281 41089 21315 41123
rect 21315 41089 21324 41123
rect 21272 41080 21324 41089
rect 23664 41123 23716 41132
rect 23664 41089 23673 41123
rect 23673 41089 23707 41123
rect 23707 41089 23716 41123
rect 23664 41080 23716 41089
rect 23848 41123 23900 41132
rect 23848 41089 23857 41123
rect 23857 41089 23891 41123
rect 23891 41089 23900 41123
rect 23848 41080 23900 41089
rect 24032 41080 24084 41132
rect 24676 41080 24728 41132
rect 25320 41080 25372 41132
rect 26792 41080 26844 41132
rect 29000 41080 29052 41132
rect 29552 41123 29604 41132
rect 29552 41089 29561 41123
rect 29561 41089 29595 41123
rect 29595 41089 29604 41123
rect 29552 41080 29604 41089
rect 30288 41080 30340 41132
rect 30932 41123 30984 41132
rect 30932 41089 30941 41123
rect 30941 41089 30975 41123
rect 30975 41089 30984 41123
rect 30932 41080 30984 41089
rect 32404 41123 32456 41132
rect 21180 41012 21232 41064
rect 23388 41012 23440 41064
rect 24308 41055 24360 41064
rect 24308 41021 24317 41055
rect 24317 41021 24351 41055
rect 24351 41021 24360 41055
rect 24308 41012 24360 41021
rect 26976 41055 27028 41064
rect 26976 41021 26985 41055
rect 26985 41021 27019 41055
rect 27019 41021 27028 41055
rect 26976 41012 27028 41021
rect 27252 41055 27304 41064
rect 27252 41021 27261 41055
rect 27261 41021 27295 41055
rect 27295 41021 27304 41055
rect 27252 41012 27304 41021
rect 29828 41055 29880 41064
rect 20904 40944 20956 40996
rect 22744 40944 22796 40996
rect 26240 40944 26292 40996
rect 26884 40944 26936 40996
rect 17500 40919 17552 40928
rect 17500 40885 17509 40919
rect 17509 40885 17543 40919
rect 17543 40885 17552 40919
rect 17500 40876 17552 40885
rect 23112 40919 23164 40928
rect 23112 40885 23121 40919
rect 23121 40885 23155 40919
rect 23155 40885 23164 40919
rect 23112 40876 23164 40885
rect 23756 40919 23808 40928
rect 23756 40885 23765 40919
rect 23765 40885 23799 40919
rect 23799 40885 23808 40919
rect 23756 40876 23808 40885
rect 24400 40919 24452 40928
rect 24400 40885 24409 40919
rect 24409 40885 24443 40919
rect 24443 40885 24452 40919
rect 24400 40876 24452 40885
rect 25044 40876 25096 40928
rect 26332 40919 26384 40928
rect 26332 40885 26341 40919
rect 26341 40885 26375 40919
rect 26375 40885 26384 40919
rect 26332 40876 26384 40885
rect 26516 40876 26568 40928
rect 27160 40876 27212 40928
rect 29828 41021 29837 41055
rect 29837 41021 29871 41055
rect 29871 41021 29880 41055
rect 29828 41012 29880 41021
rect 29920 41055 29972 41064
rect 29920 41021 29929 41055
rect 29929 41021 29963 41055
rect 29963 41021 29972 41055
rect 29920 41012 29972 41021
rect 28448 40944 28500 40996
rect 29736 40944 29788 40996
rect 32404 41089 32413 41123
rect 32413 41089 32447 41123
rect 32447 41089 32456 41123
rect 32404 41080 32456 41089
rect 32588 41123 32640 41132
rect 32588 41089 32597 41123
rect 32597 41089 32631 41123
rect 32631 41089 32640 41123
rect 32588 41080 32640 41089
rect 33416 41123 33468 41132
rect 33416 41089 33425 41123
rect 33425 41089 33459 41123
rect 33459 41089 33468 41123
rect 33416 41080 33468 41089
rect 34152 41080 34204 41132
rect 34704 41080 34756 41132
rect 35900 41080 35952 41132
rect 28540 40876 28592 40928
rect 29644 40876 29696 40928
rect 31208 40919 31260 40928
rect 31208 40885 31217 40919
rect 31217 40885 31251 40919
rect 31251 40885 31260 40919
rect 31208 40876 31260 40885
rect 33232 40876 33284 40928
rect 34244 41012 34296 41064
rect 36728 41123 36780 41132
rect 36728 41089 36737 41123
rect 36737 41089 36771 41123
rect 36771 41089 36780 41123
rect 36728 41080 36780 41089
rect 37832 41080 37884 41132
rect 38108 41123 38160 41132
rect 38108 41089 38117 41123
rect 38117 41089 38151 41123
rect 38151 41089 38160 41123
rect 38108 41080 38160 41089
rect 38200 41055 38252 41064
rect 38200 41021 38234 41055
rect 38234 41021 38252 41055
rect 38660 41080 38712 41132
rect 39212 41080 39264 41132
rect 39396 41123 39448 41132
rect 39396 41089 39405 41123
rect 39405 41089 39439 41123
rect 39439 41089 39448 41123
rect 39396 41080 39448 41089
rect 38200 41012 38252 41021
rect 35808 40919 35860 40928
rect 35808 40885 35817 40919
rect 35817 40885 35851 40919
rect 35851 40885 35860 40919
rect 35808 40876 35860 40885
rect 37648 40876 37700 40928
rect 40408 40919 40460 40928
rect 40408 40885 40417 40919
rect 40417 40885 40451 40919
rect 40451 40885 40460 40919
rect 40408 40876 40460 40885
rect 41512 40876 41564 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 16028 40715 16080 40724
rect 16028 40681 16037 40715
rect 16037 40681 16071 40715
rect 16071 40681 16080 40715
rect 16028 40672 16080 40681
rect 16580 40672 16632 40724
rect 17132 40715 17184 40724
rect 17132 40681 17141 40715
rect 17141 40681 17175 40715
rect 17175 40681 17184 40715
rect 17132 40672 17184 40681
rect 18604 40672 18656 40724
rect 20260 40672 20312 40724
rect 27252 40672 27304 40724
rect 30932 40672 30984 40724
rect 32404 40672 32456 40724
rect 34612 40672 34664 40724
rect 16672 40647 16724 40656
rect 16672 40613 16681 40647
rect 16681 40613 16715 40647
rect 16715 40613 16724 40647
rect 16672 40604 16724 40613
rect 16948 40604 17000 40656
rect 18972 40604 19024 40656
rect 18144 40536 18196 40588
rect 18512 40536 18564 40588
rect 19432 40536 19484 40588
rect 16028 40332 16080 40384
rect 17684 40443 17736 40452
rect 17684 40409 17693 40443
rect 17693 40409 17727 40443
rect 17727 40409 17736 40443
rect 17684 40400 17736 40409
rect 18052 40468 18104 40520
rect 18788 40468 18840 40520
rect 20720 40511 20772 40520
rect 20720 40477 20729 40511
rect 20729 40477 20763 40511
rect 20763 40477 20772 40511
rect 20720 40468 20772 40477
rect 20904 40511 20956 40520
rect 20904 40477 20913 40511
rect 20913 40477 20947 40511
rect 20947 40477 20956 40511
rect 20904 40468 20956 40477
rect 23664 40604 23716 40656
rect 27712 40604 27764 40656
rect 23296 40536 23348 40588
rect 24400 40536 24452 40588
rect 18236 40400 18288 40452
rect 18880 40400 18932 40452
rect 19340 40400 19392 40452
rect 20812 40400 20864 40452
rect 23388 40468 23440 40520
rect 23664 40511 23716 40520
rect 23664 40477 23673 40511
rect 23673 40477 23707 40511
rect 23707 40477 23716 40511
rect 24584 40511 24636 40520
rect 23664 40468 23716 40477
rect 18696 40332 18748 40384
rect 21916 40332 21968 40384
rect 22468 40332 22520 40384
rect 24124 40400 24176 40452
rect 24584 40477 24593 40511
rect 24593 40477 24627 40511
rect 24627 40477 24636 40511
rect 24584 40468 24636 40477
rect 26332 40536 26384 40588
rect 26608 40579 26660 40588
rect 26608 40545 26617 40579
rect 26617 40545 26651 40579
rect 26651 40545 26660 40579
rect 26608 40536 26660 40545
rect 26056 40468 26108 40520
rect 26792 40511 26844 40520
rect 26792 40477 26801 40511
rect 26801 40477 26835 40511
rect 26835 40477 26844 40511
rect 26792 40468 26844 40477
rect 27528 40468 27580 40520
rect 28540 40604 28592 40656
rect 31484 40604 31536 40656
rect 28908 40579 28960 40588
rect 28908 40545 28917 40579
rect 28917 40545 28951 40579
rect 28951 40545 28960 40579
rect 28908 40536 28960 40545
rect 29828 40579 29880 40588
rect 29828 40545 29837 40579
rect 29837 40545 29871 40579
rect 29871 40545 29880 40579
rect 29828 40536 29880 40545
rect 30748 40511 30800 40520
rect 24216 40332 24268 40384
rect 26884 40400 26936 40452
rect 27344 40400 27396 40452
rect 30748 40477 30757 40511
rect 30757 40477 30791 40511
rect 30791 40477 30800 40511
rect 30748 40468 30800 40477
rect 30840 40511 30892 40520
rect 30840 40477 30849 40511
rect 30849 40477 30883 40511
rect 30883 40477 30892 40511
rect 30840 40468 30892 40477
rect 31024 40468 31076 40520
rect 33416 40604 33468 40656
rect 33232 40579 33284 40588
rect 33232 40545 33241 40579
rect 33241 40545 33275 40579
rect 33275 40545 33284 40579
rect 33232 40536 33284 40545
rect 33784 40536 33836 40588
rect 34152 40536 34204 40588
rect 33416 40511 33468 40520
rect 31392 40400 31444 40452
rect 33416 40477 33425 40511
rect 33425 40477 33459 40511
rect 33459 40477 33468 40511
rect 33416 40468 33468 40477
rect 33508 40511 33560 40520
rect 33508 40477 33517 40511
rect 33517 40477 33551 40511
rect 33551 40477 33560 40511
rect 34704 40511 34756 40520
rect 33508 40468 33560 40477
rect 32956 40400 33008 40452
rect 34704 40477 34713 40511
rect 34713 40477 34747 40511
rect 34747 40477 34756 40511
rect 34704 40468 34756 40477
rect 35348 40511 35400 40520
rect 35348 40477 35357 40511
rect 35357 40477 35391 40511
rect 35391 40477 35400 40511
rect 35348 40468 35400 40477
rect 36176 40672 36228 40724
rect 41052 40715 41104 40724
rect 41052 40681 41061 40715
rect 41061 40681 41095 40715
rect 41095 40681 41104 40715
rect 41052 40672 41104 40681
rect 35900 40604 35952 40656
rect 35808 40536 35860 40588
rect 37832 40604 37884 40656
rect 38384 40604 38436 40656
rect 36636 40511 36688 40520
rect 36636 40477 36645 40511
rect 36645 40477 36679 40511
rect 36679 40477 36688 40511
rect 36636 40468 36688 40477
rect 36728 40468 36780 40520
rect 37096 40468 37148 40520
rect 38108 40468 38160 40520
rect 38660 40468 38712 40520
rect 39212 40511 39264 40520
rect 39212 40477 39221 40511
rect 39221 40477 39255 40511
rect 39255 40477 39264 40511
rect 39212 40468 39264 40477
rect 40040 40511 40092 40520
rect 40040 40477 40049 40511
rect 40049 40477 40083 40511
rect 40083 40477 40092 40511
rect 40040 40468 40092 40477
rect 33876 40400 33928 40452
rect 38476 40443 38528 40452
rect 38476 40409 38485 40443
rect 38485 40409 38519 40443
rect 38519 40409 38528 40443
rect 38476 40400 38528 40409
rect 39672 40400 39724 40452
rect 41512 40400 41564 40452
rect 25780 40375 25832 40384
rect 25780 40341 25789 40375
rect 25789 40341 25823 40375
rect 25823 40341 25832 40375
rect 25780 40332 25832 40341
rect 26240 40332 26292 40384
rect 26516 40332 26568 40384
rect 30564 40375 30616 40384
rect 30564 40341 30573 40375
rect 30573 40341 30607 40375
rect 30607 40341 30616 40375
rect 30564 40332 30616 40341
rect 31576 40332 31628 40384
rect 31760 40332 31812 40384
rect 35348 40332 35400 40384
rect 35624 40332 35676 40384
rect 38108 40332 38160 40384
rect 40408 40332 40460 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 16764 40128 16816 40180
rect 20720 40128 20772 40180
rect 23940 40128 23992 40180
rect 16948 40060 17000 40112
rect 17500 40060 17552 40112
rect 17960 40060 18012 40112
rect 19432 39992 19484 40044
rect 19984 39992 20036 40044
rect 20812 39992 20864 40044
rect 21272 39992 21324 40044
rect 18052 39924 18104 39976
rect 22376 40035 22428 40044
rect 22376 40001 22385 40035
rect 22385 40001 22419 40035
rect 22419 40001 22428 40035
rect 22376 39992 22428 40001
rect 23296 40035 23348 40044
rect 23296 40001 23305 40035
rect 23305 40001 23339 40035
rect 23339 40001 23348 40035
rect 23296 39992 23348 40001
rect 22836 39967 22888 39976
rect 22836 39933 22845 39967
rect 22845 39933 22879 39967
rect 22879 39933 22888 39967
rect 22836 39924 22888 39933
rect 23940 40035 23992 40044
rect 23940 40001 23949 40035
rect 23949 40001 23983 40035
rect 23983 40001 23992 40035
rect 24216 40035 24268 40044
rect 23940 39992 23992 40001
rect 24216 40001 24225 40035
rect 24225 40001 24259 40035
rect 24259 40001 24268 40035
rect 24216 39992 24268 40001
rect 24584 39992 24636 40044
rect 25780 40128 25832 40180
rect 27068 40128 27120 40180
rect 28080 40171 28132 40180
rect 28080 40137 28089 40171
rect 28089 40137 28123 40171
rect 28123 40137 28132 40171
rect 28080 40128 28132 40137
rect 31208 40128 31260 40180
rect 32220 40171 32272 40180
rect 32220 40137 32229 40171
rect 32229 40137 32263 40171
rect 32263 40137 32272 40171
rect 32220 40128 32272 40137
rect 33508 40128 33560 40180
rect 39396 40171 39448 40180
rect 26608 40060 26660 40112
rect 27160 40060 27212 40112
rect 27528 40060 27580 40112
rect 26332 39992 26384 40044
rect 27344 40035 27396 40044
rect 27344 40001 27353 40035
rect 27353 40001 27387 40035
rect 27387 40001 27396 40035
rect 27344 39992 27396 40001
rect 29736 40060 29788 40112
rect 34152 40060 34204 40112
rect 24124 39967 24176 39976
rect 24124 39933 24133 39967
rect 24133 39933 24167 39967
rect 24167 39933 24176 39967
rect 24124 39924 24176 39933
rect 24952 39924 25004 39976
rect 17316 39788 17368 39840
rect 17500 39788 17552 39840
rect 24216 39856 24268 39908
rect 27068 39967 27120 39976
rect 27068 39933 27077 39967
rect 27077 39933 27111 39967
rect 27111 39933 27120 39967
rect 27068 39924 27120 39933
rect 27436 39924 27488 39976
rect 30012 39967 30064 39976
rect 30012 39933 30021 39967
rect 30021 39933 30055 39967
rect 30055 39933 30064 39967
rect 30012 39924 30064 39933
rect 30564 39992 30616 40044
rect 31116 40035 31168 40044
rect 31116 40001 31125 40035
rect 31125 40001 31159 40035
rect 31159 40001 31168 40035
rect 31116 39992 31168 40001
rect 31760 39992 31812 40044
rect 32956 39992 33008 40044
rect 33324 40035 33376 40044
rect 30748 39924 30800 39976
rect 33324 40001 33333 40035
rect 33333 40001 33367 40035
rect 33367 40001 33376 40035
rect 33324 39992 33376 40001
rect 34796 39992 34848 40044
rect 33508 39924 33560 39976
rect 34152 39924 34204 39976
rect 18788 39831 18840 39840
rect 18788 39797 18797 39831
rect 18797 39797 18831 39831
rect 18831 39797 18840 39831
rect 18788 39788 18840 39797
rect 21180 39831 21232 39840
rect 21180 39797 21189 39831
rect 21189 39797 21223 39831
rect 21223 39797 21232 39831
rect 21180 39788 21232 39797
rect 23480 39788 23532 39840
rect 24492 39788 24544 39840
rect 24952 39788 25004 39840
rect 27344 39856 27396 39908
rect 28080 39856 28132 39908
rect 31668 39856 31720 39908
rect 25504 39831 25556 39840
rect 25504 39797 25513 39831
rect 25513 39797 25547 39831
rect 25547 39797 25556 39831
rect 25504 39788 25556 39797
rect 27160 39831 27212 39840
rect 27160 39797 27169 39831
rect 27169 39797 27203 39831
rect 27203 39797 27212 39831
rect 27160 39788 27212 39797
rect 33232 39788 33284 39840
rect 39396 40137 39405 40171
rect 39405 40137 39439 40171
rect 39439 40137 39448 40171
rect 39396 40128 39448 40137
rect 40040 40128 40092 40180
rect 40408 40128 40460 40180
rect 41052 40171 41104 40180
rect 41052 40137 41061 40171
rect 41061 40137 41095 40171
rect 41095 40137 41104 40171
rect 41052 40128 41104 40137
rect 36176 40035 36228 40044
rect 36176 40001 36185 40035
rect 36185 40001 36219 40035
rect 36219 40001 36228 40035
rect 36176 39992 36228 40001
rect 36360 40035 36412 40044
rect 36360 40001 36369 40035
rect 36369 40001 36403 40035
rect 36403 40001 36412 40035
rect 36360 39992 36412 40001
rect 37556 39992 37608 40044
rect 38108 40035 38160 40044
rect 38108 40001 38117 40035
rect 38117 40001 38151 40035
rect 38151 40001 38160 40035
rect 38108 39992 38160 40001
rect 38660 40060 38712 40112
rect 38936 40035 38988 40044
rect 38936 40001 38945 40035
rect 38945 40001 38979 40035
rect 38979 40001 38988 40035
rect 39672 40035 39724 40044
rect 38936 39992 38988 40001
rect 38660 39924 38712 39976
rect 39672 40001 39681 40035
rect 39681 40001 39715 40035
rect 39715 40001 39724 40035
rect 39672 39992 39724 40001
rect 39856 40035 39908 40044
rect 39856 40001 39865 40035
rect 39865 40001 39899 40035
rect 39899 40001 39908 40035
rect 39856 39992 39908 40001
rect 41052 39924 41104 39976
rect 53564 40035 53616 40044
rect 53564 40001 53573 40035
rect 53573 40001 53607 40035
rect 53607 40001 53616 40035
rect 53564 39992 53616 40001
rect 35808 39856 35860 39908
rect 38292 39899 38344 39908
rect 38292 39865 38301 39899
rect 38301 39865 38335 39899
rect 38335 39865 38344 39899
rect 38292 39856 38344 39865
rect 39856 39856 39908 39908
rect 52828 39856 52880 39908
rect 35624 39788 35676 39840
rect 37464 39788 37516 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 21180 39584 21232 39636
rect 22192 39584 22244 39636
rect 22376 39627 22428 39636
rect 22376 39593 22385 39627
rect 22385 39593 22419 39627
rect 22419 39593 22428 39627
rect 22376 39584 22428 39593
rect 22468 39584 22520 39636
rect 23664 39584 23716 39636
rect 26884 39584 26936 39636
rect 31484 39584 31536 39636
rect 32680 39627 32732 39636
rect 32680 39593 32689 39627
rect 32689 39593 32723 39627
rect 32723 39593 32732 39627
rect 32680 39584 32732 39593
rect 33140 39584 33192 39636
rect 33324 39627 33376 39636
rect 33324 39593 33333 39627
rect 33333 39593 33367 39627
rect 33367 39593 33376 39627
rect 33324 39584 33376 39593
rect 33784 39584 33836 39636
rect 34152 39584 34204 39636
rect 35348 39584 35400 39636
rect 38568 39584 38620 39636
rect 41512 39627 41564 39636
rect 41512 39593 41521 39627
rect 41521 39593 41555 39627
rect 41555 39593 41564 39627
rect 41512 39584 41564 39593
rect 15476 39448 15528 39500
rect 18052 39448 18104 39500
rect 18788 39448 18840 39500
rect 16764 39423 16816 39432
rect 16764 39389 16773 39423
rect 16773 39389 16807 39423
rect 16807 39389 16816 39423
rect 16764 39380 16816 39389
rect 16948 39423 17000 39432
rect 16948 39389 16957 39423
rect 16957 39389 16991 39423
rect 16991 39389 17000 39423
rect 16948 39380 17000 39389
rect 17316 39380 17368 39432
rect 17776 39423 17828 39432
rect 17776 39389 17785 39423
rect 17785 39389 17819 39423
rect 17819 39389 17828 39423
rect 17776 39380 17828 39389
rect 19340 39380 19392 39432
rect 20444 39423 20496 39432
rect 20444 39389 20453 39423
rect 20453 39389 20487 39423
rect 20487 39389 20496 39423
rect 20444 39380 20496 39389
rect 16304 39312 16356 39364
rect 17408 39312 17460 39364
rect 20812 39312 20864 39364
rect 25504 39516 25556 39568
rect 23480 39491 23532 39500
rect 23480 39457 23489 39491
rect 23489 39457 23523 39491
rect 23523 39457 23532 39491
rect 23480 39448 23532 39457
rect 22376 39380 22428 39432
rect 23664 39423 23716 39432
rect 22560 39355 22612 39364
rect 22560 39321 22569 39355
rect 22569 39321 22603 39355
rect 22603 39321 22612 39355
rect 22560 39312 22612 39321
rect 22744 39355 22796 39364
rect 22744 39321 22753 39355
rect 22753 39321 22787 39355
rect 22787 39321 22796 39355
rect 22744 39312 22796 39321
rect 23112 39312 23164 39364
rect 23664 39389 23673 39423
rect 23673 39389 23707 39423
rect 23707 39389 23716 39423
rect 23664 39380 23716 39389
rect 23756 39380 23808 39432
rect 24492 39380 24544 39432
rect 15476 39287 15528 39296
rect 15476 39253 15485 39287
rect 15485 39253 15519 39287
rect 15519 39253 15528 39287
rect 15476 39244 15528 39253
rect 15936 39244 15988 39296
rect 17500 39287 17552 39296
rect 17500 39253 17509 39287
rect 17509 39253 17543 39287
rect 17543 39253 17552 39287
rect 17500 39244 17552 39253
rect 19432 39244 19484 39296
rect 20720 39244 20772 39296
rect 22468 39244 22520 39296
rect 23296 39244 23348 39296
rect 24308 39244 24360 39296
rect 24860 39380 24912 39432
rect 24952 39423 25004 39432
rect 24952 39389 24961 39423
rect 24961 39389 24995 39423
rect 24995 39389 25004 39423
rect 24952 39380 25004 39389
rect 30840 39516 30892 39568
rect 26976 39491 27028 39500
rect 26976 39457 26985 39491
rect 26985 39457 27019 39491
rect 27019 39457 27028 39491
rect 26976 39448 27028 39457
rect 31116 39448 31168 39500
rect 34428 39516 34480 39568
rect 30748 39423 30800 39432
rect 30748 39389 30757 39423
rect 30757 39389 30791 39423
rect 30791 39389 30800 39423
rect 30748 39380 30800 39389
rect 26424 39312 26476 39364
rect 26516 39355 26568 39364
rect 26516 39321 26525 39355
rect 26525 39321 26559 39355
rect 26559 39321 26568 39355
rect 26516 39312 26568 39321
rect 29920 39312 29972 39364
rect 25136 39287 25188 39296
rect 25136 39253 25145 39287
rect 25145 39253 25179 39287
rect 25179 39253 25188 39287
rect 25136 39244 25188 39253
rect 26332 39287 26384 39296
rect 26332 39253 26341 39287
rect 26341 39253 26375 39287
rect 26375 39253 26384 39287
rect 26332 39244 26384 39253
rect 27252 39244 27304 39296
rect 30656 39355 30708 39364
rect 30656 39321 30665 39355
rect 30665 39321 30699 39355
rect 30699 39321 30708 39355
rect 32588 39448 32640 39500
rect 33324 39448 33376 39500
rect 33416 39380 33468 39432
rect 35348 39448 35400 39500
rect 36176 39448 36228 39500
rect 40040 39516 40092 39568
rect 38292 39448 38344 39500
rect 34796 39380 34848 39432
rect 35256 39380 35308 39432
rect 35624 39423 35676 39432
rect 35624 39389 35633 39423
rect 35633 39389 35667 39423
rect 35667 39389 35676 39423
rect 35624 39380 35676 39389
rect 36360 39423 36412 39432
rect 36360 39389 36369 39423
rect 36369 39389 36403 39423
rect 36403 39389 36412 39423
rect 36360 39380 36412 39389
rect 37372 39380 37424 39432
rect 37556 39380 37608 39432
rect 38476 39423 38528 39432
rect 38476 39389 38485 39423
rect 38485 39389 38519 39423
rect 38519 39389 38528 39423
rect 38476 39380 38528 39389
rect 30656 39312 30708 39321
rect 32956 39312 33008 39364
rect 33508 39355 33560 39364
rect 33508 39321 33517 39355
rect 33517 39321 33551 39355
rect 33551 39321 33560 39355
rect 33508 39312 33560 39321
rect 34980 39355 35032 39364
rect 34980 39321 34989 39355
rect 34989 39321 35023 39355
rect 35023 39321 35032 39355
rect 34980 39312 35032 39321
rect 38200 39312 38252 39364
rect 39856 39312 39908 39364
rect 30840 39244 30892 39296
rect 31024 39244 31076 39296
rect 31392 39287 31444 39296
rect 31392 39253 31401 39287
rect 31401 39253 31435 39287
rect 31435 39253 31444 39287
rect 31392 39244 31444 39253
rect 33048 39244 33100 39296
rect 33784 39244 33836 39296
rect 34704 39244 34756 39296
rect 35808 39244 35860 39296
rect 37280 39287 37332 39296
rect 37280 39253 37289 39287
rect 37289 39253 37323 39287
rect 37323 39253 37332 39287
rect 37280 39244 37332 39253
rect 39028 39244 39080 39296
rect 40408 39287 40460 39296
rect 40408 39253 40417 39287
rect 40417 39253 40451 39287
rect 40451 39253 40460 39287
rect 40408 39244 40460 39253
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 15936 39040 15988 39092
rect 17776 39040 17828 39092
rect 19340 39040 19392 39092
rect 20168 39083 20220 39092
rect 16764 38972 16816 39024
rect 18696 39015 18748 39024
rect 1584 38904 1636 38956
rect 15936 38947 15988 38956
rect 15936 38913 15945 38947
rect 15945 38913 15979 38947
rect 15979 38913 15988 38947
rect 15936 38904 15988 38913
rect 16672 38904 16724 38956
rect 17408 38904 17460 38956
rect 18328 38904 18380 38956
rect 18696 38981 18705 39015
rect 18705 38981 18739 39015
rect 18739 38981 18748 39015
rect 18696 38972 18748 38981
rect 20168 39049 20177 39083
rect 20177 39049 20211 39083
rect 20211 39049 20220 39083
rect 20168 39040 20220 39049
rect 20444 39040 20496 39092
rect 20628 39083 20680 39092
rect 20628 39049 20637 39083
rect 20637 39049 20671 39083
rect 20671 39049 20680 39083
rect 20628 39040 20680 39049
rect 22376 39083 22428 39092
rect 22376 39049 22385 39083
rect 22385 39049 22419 39083
rect 22419 39049 22428 39083
rect 22376 39040 22428 39049
rect 22836 39040 22888 39092
rect 20720 38972 20772 39024
rect 23756 39040 23808 39092
rect 24952 38972 25004 39024
rect 26240 39040 26292 39092
rect 26332 39040 26384 39092
rect 29552 39083 29604 39092
rect 29552 39049 29561 39083
rect 29561 39049 29595 39083
rect 29595 39049 29604 39083
rect 29552 39040 29604 39049
rect 29920 39083 29972 39092
rect 29920 39049 29929 39083
rect 29929 39049 29963 39083
rect 29963 39049 29972 39083
rect 29920 39040 29972 39049
rect 26516 38972 26568 39024
rect 20812 38904 20864 38956
rect 21088 38947 21140 38956
rect 21088 38913 21097 38947
rect 21097 38913 21131 38947
rect 21131 38913 21140 38947
rect 21088 38904 21140 38913
rect 21824 38904 21876 38956
rect 22008 38947 22060 38956
rect 22008 38913 22017 38947
rect 22017 38913 22051 38947
rect 22051 38913 22060 38947
rect 22008 38904 22060 38913
rect 22560 38904 22612 38956
rect 23296 38947 23348 38956
rect 23296 38913 23305 38947
rect 23305 38913 23339 38947
rect 23339 38913 23348 38947
rect 23296 38904 23348 38913
rect 23940 38904 23992 38956
rect 24860 38904 24912 38956
rect 25228 38904 25280 38956
rect 27160 38947 27212 38956
rect 27160 38913 27169 38947
rect 27169 38913 27203 38947
rect 27203 38913 27212 38947
rect 27160 38904 27212 38913
rect 27252 38904 27304 38956
rect 27436 38947 27488 38956
rect 27436 38913 27445 38947
rect 27445 38913 27479 38947
rect 27479 38913 27488 38947
rect 27436 38904 27488 38913
rect 19524 38836 19576 38888
rect 20996 38879 21048 38888
rect 19432 38768 19484 38820
rect 20996 38845 21005 38879
rect 21005 38845 21039 38879
rect 21039 38845 21048 38879
rect 20996 38836 21048 38845
rect 21272 38879 21324 38888
rect 21272 38845 21281 38879
rect 21281 38845 21315 38879
rect 21315 38845 21324 38879
rect 21272 38836 21324 38845
rect 22192 38836 22244 38888
rect 30564 38904 30616 38956
rect 31392 38972 31444 39024
rect 31576 39015 31628 39024
rect 31576 38981 31585 39015
rect 31585 38981 31619 39015
rect 31619 38981 31628 39015
rect 31576 38972 31628 38981
rect 30932 38947 30984 38956
rect 15384 38700 15436 38752
rect 17500 38700 17552 38752
rect 25228 38768 25280 38820
rect 27252 38768 27304 38820
rect 20996 38700 21048 38752
rect 21456 38700 21508 38752
rect 22192 38700 22244 38752
rect 24400 38700 24452 38752
rect 24676 38700 24728 38752
rect 26332 38743 26384 38752
rect 26332 38709 26341 38743
rect 26341 38709 26375 38743
rect 26375 38709 26384 38743
rect 26332 38700 26384 38709
rect 30472 38836 30524 38888
rect 30932 38913 30941 38947
rect 30941 38913 30975 38947
rect 30975 38913 30984 38947
rect 30932 38904 30984 38913
rect 31024 38947 31076 38956
rect 31024 38913 31033 38947
rect 31033 38913 31067 38947
rect 31067 38913 31076 38947
rect 31024 38904 31076 38913
rect 32956 38904 33008 38956
rect 31208 38836 31260 38888
rect 30288 38768 30340 38820
rect 36360 39040 36412 39092
rect 37280 39040 37332 39092
rect 38384 39040 38436 39092
rect 38568 39040 38620 39092
rect 40040 39083 40092 39092
rect 40040 39049 40049 39083
rect 40049 39049 40083 39083
rect 40083 39049 40092 39083
rect 40040 39040 40092 39049
rect 34980 38972 35032 39024
rect 35532 38972 35584 39024
rect 34152 38904 34204 38956
rect 34428 38947 34480 38956
rect 34428 38913 34437 38947
rect 34437 38913 34471 38947
rect 34471 38913 34480 38947
rect 34428 38904 34480 38913
rect 35256 38947 35308 38956
rect 35256 38913 35265 38947
rect 35265 38913 35299 38947
rect 35299 38913 35308 38947
rect 35256 38904 35308 38913
rect 35624 38904 35676 38956
rect 33416 38836 33468 38888
rect 37280 38904 37332 38956
rect 38384 38904 38436 38956
rect 38660 38904 38712 38956
rect 37464 38836 37516 38888
rect 38936 38879 38988 38888
rect 38936 38845 38945 38879
rect 38945 38845 38979 38879
rect 38979 38845 38988 38879
rect 38936 38836 38988 38845
rect 38844 38768 38896 38820
rect 31208 38700 31260 38752
rect 32496 38700 32548 38752
rect 33416 38700 33468 38752
rect 33784 38700 33836 38752
rect 34060 38743 34112 38752
rect 34060 38709 34069 38743
rect 34069 38709 34103 38743
rect 34103 38709 34112 38743
rect 34060 38700 34112 38709
rect 34796 38700 34848 38752
rect 35992 38743 36044 38752
rect 35992 38709 36001 38743
rect 36001 38709 36035 38743
rect 36035 38709 36044 38743
rect 35992 38700 36044 38709
rect 36452 38743 36504 38752
rect 36452 38709 36461 38743
rect 36461 38709 36495 38743
rect 36495 38709 36504 38743
rect 36452 38700 36504 38709
rect 37280 38743 37332 38752
rect 37280 38709 37289 38743
rect 37289 38709 37323 38743
rect 37323 38709 37332 38743
rect 37280 38700 37332 38709
rect 37464 38743 37516 38752
rect 37464 38709 37473 38743
rect 37473 38709 37507 38743
rect 37507 38709 37516 38743
rect 37464 38700 37516 38709
rect 40040 38700 40092 38752
rect 40408 38700 40460 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 1584 38539 1636 38548
rect 1584 38505 1593 38539
rect 1593 38505 1627 38539
rect 1627 38505 1636 38539
rect 1584 38496 1636 38505
rect 16672 38539 16724 38548
rect 16672 38505 16681 38539
rect 16681 38505 16715 38539
rect 16715 38505 16724 38539
rect 16672 38496 16724 38505
rect 26516 38496 26568 38548
rect 27712 38496 27764 38548
rect 30012 38496 30064 38548
rect 30932 38496 30984 38548
rect 32956 38539 33008 38548
rect 32956 38505 32965 38539
rect 32965 38505 32999 38539
rect 32999 38505 33008 38539
rect 32956 38496 33008 38505
rect 34796 38539 34848 38548
rect 34796 38505 34805 38539
rect 34805 38505 34839 38539
rect 34839 38505 34848 38539
rect 34796 38496 34848 38505
rect 35348 38496 35400 38548
rect 36452 38496 36504 38548
rect 25320 38428 25372 38480
rect 15476 38292 15528 38344
rect 16304 38267 16356 38276
rect 16304 38233 16313 38267
rect 16313 38233 16347 38267
rect 16347 38233 16356 38267
rect 16304 38224 16356 38233
rect 16488 38267 16540 38276
rect 16488 38233 16497 38267
rect 16497 38233 16531 38267
rect 16531 38233 16540 38267
rect 16488 38224 16540 38233
rect 16396 38156 16448 38208
rect 17224 38335 17276 38344
rect 17224 38301 17233 38335
rect 17233 38301 17267 38335
rect 17267 38301 17276 38335
rect 17224 38292 17276 38301
rect 17500 38335 17552 38344
rect 17500 38301 17509 38335
rect 17509 38301 17543 38335
rect 17543 38301 17552 38335
rect 17500 38292 17552 38301
rect 18144 38335 18196 38344
rect 18144 38301 18153 38335
rect 18153 38301 18187 38335
rect 18187 38301 18196 38335
rect 18144 38292 18196 38301
rect 18328 38335 18380 38344
rect 18328 38301 18337 38335
rect 18337 38301 18371 38335
rect 18371 38301 18380 38335
rect 18328 38292 18380 38301
rect 19248 38335 19300 38344
rect 19248 38301 19257 38335
rect 19257 38301 19291 38335
rect 19291 38301 19300 38335
rect 19248 38292 19300 38301
rect 19524 38292 19576 38344
rect 20168 38335 20220 38344
rect 20168 38301 20177 38335
rect 20177 38301 20211 38335
rect 20211 38301 20220 38335
rect 20168 38292 20220 38301
rect 21272 38360 21324 38412
rect 22008 38360 22060 38412
rect 20904 38335 20956 38344
rect 16948 38224 17000 38276
rect 20904 38301 20913 38335
rect 20913 38301 20947 38335
rect 20947 38301 20956 38335
rect 20904 38292 20956 38301
rect 21180 38335 21232 38344
rect 21180 38301 21189 38335
rect 21189 38301 21223 38335
rect 21223 38301 21232 38335
rect 21180 38292 21232 38301
rect 21640 38292 21692 38344
rect 22192 38335 22244 38344
rect 22192 38301 22201 38335
rect 22201 38301 22235 38335
rect 22235 38301 22244 38335
rect 22192 38292 22244 38301
rect 22836 38335 22888 38344
rect 22836 38301 22845 38335
rect 22845 38301 22879 38335
rect 22879 38301 22888 38335
rect 22836 38292 22888 38301
rect 24400 38335 24452 38344
rect 24400 38301 24409 38335
rect 24409 38301 24443 38335
rect 24443 38301 24452 38335
rect 24400 38292 24452 38301
rect 21088 38224 21140 38276
rect 24032 38224 24084 38276
rect 26056 38335 26108 38344
rect 26056 38301 26065 38335
rect 26065 38301 26099 38335
rect 26099 38301 26108 38335
rect 26056 38292 26108 38301
rect 26700 38471 26752 38480
rect 26700 38437 26709 38471
rect 26709 38437 26743 38471
rect 26743 38437 26752 38471
rect 26700 38428 26752 38437
rect 27344 38428 27396 38480
rect 29920 38403 29972 38412
rect 24676 38224 24728 38276
rect 26608 38224 26660 38276
rect 26884 38292 26936 38344
rect 27436 38292 27488 38344
rect 29920 38369 29929 38403
rect 29929 38369 29963 38403
rect 29963 38369 29972 38403
rect 29920 38360 29972 38369
rect 30840 38428 30892 38480
rect 35808 38428 35860 38480
rect 17684 38199 17736 38208
rect 17684 38165 17693 38199
rect 17693 38165 17727 38199
rect 17727 38165 17736 38199
rect 17684 38156 17736 38165
rect 17776 38156 17828 38208
rect 20720 38156 20772 38208
rect 20996 38199 21048 38208
rect 20996 38165 21005 38199
rect 21005 38165 21039 38199
rect 21039 38165 21048 38199
rect 20996 38156 21048 38165
rect 21364 38199 21416 38208
rect 21364 38165 21373 38199
rect 21373 38165 21407 38199
rect 21407 38165 21416 38199
rect 21364 38156 21416 38165
rect 21824 38156 21876 38208
rect 22100 38199 22152 38208
rect 22100 38165 22109 38199
rect 22109 38165 22143 38199
rect 22143 38165 22152 38199
rect 24768 38199 24820 38208
rect 22100 38156 22152 38165
rect 24768 38165 24777 38199
rect 24777 38165 24811 38199
rect 24811 38165 24820 38199
rect 24768 38156 24820 38165
rect 25228 38199 25280 38208
rect 25228 38165 25237 38199
rect 25237 38165 25271 38199
rect 25271 38165 25280 38199
rect 25228 38156 25280 38165
rect 27068 38224 27120 38276
rect 27160 38156 27212 38208
rect 30104 38156 30156 38208
rect 30564 38156 30616 38208
rect 30932 38199 30984 38208
rect 30932 38165 30941 38199
rect 30941 38165 30975 38199
rect 30975 38165 30984 38199
rect 30932 38156 30984 38165
rect 31944 38335 31996 38344
rect 31944 38301 31953 38335
rect 31953 38301 31987 38335
rect 31987 38301 31996 38335
rect 31944 38292 31996 38301
rect 32036 38335 32088 38344
rect 32036 38301 32045 38335
rect 32045 38301 32079 38335
rect 32079 38301 32088 38335
rect 32036 38292 32088 38301
rect 33416 38292 33468 38344
rect 33600 38335 33652 38344
rect 33600 38301 33609 38335
rect 33609 38301 33643 38335
rect 33643 38301 33652 38335
rect 33600 38292 33652 38301
rect 33692 38335 33744 38344
rect 33692 38301 33701 38335
rect 33701 38301 33735 38335
rect 33735 38301 33744 38335
rect 33692 38292 33744 38301
rect 32588 38224 32640 38276
rect 34060 38224 34112 38276
rect 34704 38224 34756 38276
rect 35164 38267 35216 38276
rect 35164 38233 35173 38267
rect 35173 38233 35207 38267
rect 35207 38233 35216 38267
rect 35164 38224 35216 38233
rect 35348 38292 35400 38344
rect 37188 38292 37240 38344
rect 37280 38335 37332 38344
rect 37280 38301 37289 38335
rect 37289 38301 37323 38335
rect 37323 38301 37332 38335
rect 37280 38292 37332 38301
rect 38476 38335 38528 38344
rect 38476 38301 38485 38335
rect 38485 38301 38519 38335
rect 38519 38301 38528 38335
rect 38476 38292 38528 38301
rect 35900 38224 35952 38276
rect 38384 38224 38436 38276
rect 40040 38224 40092 38276
rect 33416 38199 33468 38208
rect 33416 38165 33425 38199
rect 33425 38165 33459 38199
rect 33459 38165 33468 38199
rect 33416 38156 33468 38165
rect 35532 38156 35584 38208
rect 36636 38156 36688 38208
rect 37188 38199 37240 38208
rect 37188 38165 37197 38199
rect 37197 38165 37231 38199
rect 37231 38165 37240 38199
rect 37188 38156 37240 38165
rect 38660 38156 38712 38208
rect 39856 38199 39908 38208
rect 39856 38165 39865 38199
rect 39865 38165 39899 38199
rect 39899 38165 39908 38199
rect 39856 38156 39908 38165
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 16304 37952 16356 38004
rect 17684 37952 17736 38004
rect 19432 37952 19484 38004
rect 21180 37952 21232 38004
rect 25228 37995 25280 38004
rect 25228 37961 25237 37995
rect 25237 37961 25271 37995
rect 25271 37961 25280 37995
rect 25228 37952 25280 37961
rect 26056 37952 26108 38004
rect 17408 37859 17460 37868
rect 17408 37825 17417 37859
rect 17417 37825 17451 37859
rect 17451 37825 17460 37859
rect 17408 37816 17460 37825
rect 17776 37816 17828 37868
rect 18512 37884 18564 37936
rect 20904 37884 20956 37936
rect 16028 37655 16080 37664
rect 16028 37621 16037 37655
rect 16037 37621 16071 37655
rect 16071 37621 16080 37655
rect 18696 37748 18748 37800
rect 20076 37816 20128 37868
rect 20168 37859 20220 37868
rect 20168 37825 20177 37859
rect 20177 37825 20211 37859
rect 20211 37825 20220 37859
rect 21088 37859 21140 37868
rect 20168 37816 20220 37825
rect 21088 37825 21097 37859
rect 21097 37825 21131 37859
rect 21131 37825 21140 37859
rect 21088 37816 21140 37825
rect 21364 37884 21416 37936
rect 20720 37748 20772 37800
rect 21272 37748 21324 37800
rect 21824 37791 21876 37800
rect 21824 37757 21833 37791
rect 21833 37757 21867 37791
rect 21867 37757 21876 37791
rect 21824 37748 21876 37757
rect 21088 37680 21140 37732
rect 22836 37816 22888 37868
rect 23388 37859 23440 37868
rect 23388 37825 23397 37859
rect 23397 37825 23431 37859
rect 23431 37825 23440 37859
rect 23388 37816 23440 37825
rect 22468 37748 22520 37800
rect 24308 37816 24360 37868
rect 24768 37816 24820 37868
rect 25412 37816 25464 37868
rect 26424 37859 26476 37868
rect 24676 37748 24728 37800
rect 25320 37791 25372 37800
rect 25320 37757 25329 37791
rect 25329 37757 25363 37791
rect 25363 37757 25372 37791
rect 25320 37748 25372 37757
rect 26424 37825 26433 37859
rect 26433 37825 26467 37859
rect 26467 37825 26476 37859
rect 26424 37816 26476 37825
rect 30288 37952 30340 38004
rect 30840 37952 30892 38004
rect 33416 37952 33468 38004
rect 33600 37952 33652 38004
rect 35164 37952 35216 38004
rect 35532 37952 35584 38004
rect 27068 37816 27120 37868
rect 26700 37748 26752 37800
rect 28356 37748 28408 37800
rect 30472 37748 30524 37800
rect 31024 37816 31076 37868
rect 31576 37816 31628 37868
rect 32036 37816 32088 37868
rect 32588 37859 32640 37868
rect 32588 37825 32597 37859
rect 32597 37825 32631 37859
rect 32631 37825 32640 37859
rect 32588 37816 32640 37825
rect 33048 37859 33100 37868
rect 33048 37825 33057 37859
rect 33057 37825 33091 37859
rect 33091 37825 33100 37859
rect 33048 37816 33100 37825
rect 33232 37816 33284 37868
rect 33968 37859 34020 37868
rect 33968 37825 33977 37859
rect 33977 37825 34011 37859
rect 34011 37825 34020 37859
rect 33968 37816 34020 37825
rect 34612 37816 34664 37868
rect 35808 37816 35860 37868
rect 37280 37884 37332 37936
rect 36452 37816 36504 37868
rect 37740 37859 37792 37868
rect 37740 37825 37779 37859
rect 37779 37825 37792 37859
rect 37740 37816 37792 37825
rect 38752 37816 38804 37868
rect 31944 37748 31996 37800
rect 16028 37612 16080 37621
rect 18512 37612 18564 37664
rect 19708 37655 19760 37664
rect 19708 37621 19717 37655
rect 19717 37621 19751 37655
rect 19751 37621 19760 37655
rect 19708 37612 19760 37621
rect 21456 37612 21508 37664
rect 23848 37612 23900 37664
rect 24032 37655 24084 37664
rect 24032 37621 24041 37655
rect 24041 37621 24075 37655
rect 24075 37621 24084 37655
rect 24032 37612 24084 37621
rect 26608 37680 26660 37732
rect 24676 37612 24728 37664
rect 26700 37612 26752 37664
rect 31668 37680 31720 37732
rect 33140 37680 33192 37732
rect 37556 37723 37608 37732
rect 37556 37689 37565 37723
rect 37565 37689 37599 37723
rect 37599 37689 37608 37723
rect 37556 37680 37608 37689
rect 32128 37655 32180 37664
rect 32128 37621 32137 37655
rect 32137 37621 32171 37655
rect 32171 37621 32180 37655
rect 32128 37612 32180 37621
rect 32496 37655 32548 37664
rect 32496 37621 32505 37655
rect 32505 37621 32539 37655
rect 32539 37621 32548 37655
rect 32496 37612 32548 37621
rect 33600 37612 33652 37664
rect 34152 37612 34204 37664
rect 38384 37655 38436 37664
rect 38384 37621 38393 37655
rect 38393 37621 38427 37655
rect 38427 37621 38436 37655
rect 38384 37612 38436 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 16396 37408 16448 37460
rect 17500 37451 17552 37460
rect 17500 37417 17509 37451
rect 17509 37417 17543 37451
rect 17543 37417 17552 37451
rect 17500 37408 17552 37417
rect 18236 37408 18288 37460
rect 19708 37408 19760 37460
rect 20812 37408 20864 37460
rect 17316 37340 17368 37392
rect 17776 37340 17828 37392
rect 18328 37340 18380 37392
rect 16028 37315 16080 37324
rect 16028 37281 16037 37315
rect 16037 37281 16071 37315
rect 16071 37281 16080 37315
rect 16028 37272 16080 37281
rect 17868 37315 17920 37324
rect 17868 37281 17877 37315
rect 17877 37281 17911 37315
rect 17911 37281 17920 37315
rect 17868 37272 17920 37281
rect 19432 37272 19484 37324
rect 17224 37204 17276 37256
rect 18420 37247 18472 37256
rect 18420 37213 18429 37247
rect 18429 37213 18463 37247
rect 18463 37213 18472 37247
rect 18420 37204 18472 37213
rect 18696 37247 18748 37256
rect 18696 37213 18705 37247
rect 18705 37213 18739 37247
rect 18739 37213 18748 37247
rect 18696 37204 18748 37213
rect 19248 37136 19300 37188
rect 20076 37247 20128 37256
rect 20076 37213 20085 37247
rect 20085 37213 20119 37247
rect 20119 37213 20128 37247
rect 20076 37204 20128 37213
rect 23940 37408 23992 37460
rect 26608 37408 26660 37460
rect 29920 37408 29972 37460
rect 33508 37451 33560 37460
rect 33508 37417 33517 37451
rect 33517 37417 33551 37451
rect 33551 37417 33560 37451
rect 33508 37408 33560 37417
rect 34704 37408 34756 37460
rect 35992 37408 36044 37460
rect 36360 37451 36412 37460
rect 36360 37417 36369 37451
rect 36369 37417 36403 37451
rect 36403 37417 36412 37451
rect 36360 37408 36412 37417
rect 36636 37408 36688 37460
rect 38200 37451 38252 37460
rect 22376 37383 22428 37392
rect 22376 37349 22385 37383
rect 22385 37349 22419 37383
rect 22419 37349 22428 37383
rect 22376 37340 22428 37349
rect 23664 37340 23716 37392
rect 24308 37340 24360 37392
rect 20904 37204 20956 37256
rect 22192 37272 22244 37324
rect 22284 37272 22336 37324
rect 23388 37272 23440 37324
rect 24032 37272 24084 37324
rect 24492 37204 24544 37256
rect 24676 37247 24728 37256
rect 24676 37213 24685 37247
rect 24685 37213 24719 37247
rect 24719 37213 24728 37247
rect 24676 37204 24728 37213
rect 19984 37136 20036 37188
rect 22468 37136 22520 37188
rect 24308 37136 24360 37188
rect 24860 37247 24912 37256
rect 24860 37213 24869 37247
rect 24869 37213 24903 37247
rect 24903 37213 24912 37247
rect 26700 37340 26752 37392
rect 27068 37383 27120 37392
rect 27068 37349 27077 37383
rect 27077 37349 27111 37383
rect 27111 37349 27120 37383
rect 27068 37340 27120 37349
rect 29828 37383 29880 37392
rect 29828 37349 29837 37383
rect 29837 37349 29871 37383
rect 29871 37349 29880 37383
rect 29828 37340 29880 37349
rect 24860 37204 24912 37213
rect 25412 37204 25464 37256
rect 25136 37136 25188 37188
rect 25228 37136 25280 37188
rect 26424 37272 26476 37324
rect 32404 37340 32456 37392
rect 34612 37340 34664 37392
rect 34888 37340 34940 37392
rect 37188 37340 37240 37392
rect 30932 37272 30984 37324
rect 27160 37204 27212 37256
rect 27528 37204 27580 37256
rect 27712 37204 27764 37256
rect 28356 37247 28408 37256
rect 28356 37213 28365 37247
rect 28365 37213 28399 37247
rect 28399 37213 28408 37247
rect 28356 37204 28408 37213
rect 28540 37247 28592 37256
rect 28540 37213 28549 37247
rect 28549 37213 28583 37247
rect 28583 37213 28592 37247
rect 28540 37204 28592 37213
rect 29736 37247 29788 37256
rect 29736 37213 29745 37247
rect 29745 37213 29779 37247
rect 29779 37213 29788 37247
rect 29736 37204 29788 37213
rect 29920 37247 29972 37256
rect 29920 37213 29929 37247
rect 29929 37213 29963 37247
rect 29963 37213 29972 37247
rect 29920 37204 29972 37213
rect 26884 37179 26936 37188
rect 26884 37145 26909 37179
rect 26909 37145 26936 37179
rect 26884 37136 26936 37145
rect 28908 37136 28960 37188
rect 29644 37136 29696 37188
rect 30104 37204 30156 37256
rect 30656 37204 30708 37256
rect 32588 37272 32640 37324
rect 16948 37068 17000 37120
rect 18512 37111 18564 37120
rect 18512 37077 18521 37111
rect 18521 37077 18555 37111
rect 18555 37077 18564 37111
rect 18512 37068 18564 37077
rect 20996 37111 21048 37120
rect 20996 37077 21005 37111
rect 21005 37077 21039 37111
rect 21039 37077 21048 37111
rect 20996 37068 21048 37077
rect 24216 37068 24268 37120
rect 24400 37111 24452 37120
rect 24400 37077 24409 37111
rect 24409 37077 24443 37111
rect 24443 37077 24452 37111
rect 24400 37068 24452 37077
rect 24584 37068 24636 37120
rect 27988 37068 28040 37120
rect 28724 37068 28776 37120
rect 30748 37068 30800 37120
rect 31484 37204 31536 37256
rect 31760 37247 31812 37256
rect 31760 37213 31769 37247
rect 31769 37213 31803 37247
rect 31803 37213 31812 37247
rect 31760 37204 31812 37213
rect 32220 37204 32272 37256
rect 32128 37136 32180 37188
rect 32956 37136 33008 37188
rect 33416 37136 33468 37188
rect 34244 37204 34296 37256
rect 34704 37247 34756 37256
rect 34704 37213 34713 37247
rect 34713 37213 34747 37247
rect 34747 37213 34756 37247
rect 34704 37204 34756 37213
rect 35072 37204 35124 37256
rect 35348 37136 35400 37188
rect 32404 37111 32456 37120
rect 32404 37077 32413 37111
rect 32413 37077 32447 37111
rect 32447 37077 32456 37111
rect 32404 37068 32456 37077
rect 33876 37068 33928 37120
rect 34796 37111 34848 37120
rect 34796 37077 34805 37111
rect 34805 37077 34839 37111
rect 34839 37077 34848 37111
rect 34796 37068 34848 37077
rect 37280 37204 37332 37256
rect 37556 37340 37608 37392
rect 38200 37417 38209 37451
rect 38209 37417 38243 37451
rect 38243 37417 38252 37451
rect 38200 37408 38252 37417
rect 38660 37408 38712 37460
rect 52828 37451 52880 37460
rect 52828 37417 52837 37451
rect 52837 37417 52871 37451
rect 52871 37417 52880 37451
rect 52828 37408 52880 37417
rect 37648 37247 37700 37256
rect 37372 37136 37424 37188
rect 37648 37213 37657 37247
rect 37657 37213 37691 37247
rect 37691 37213 37700 37247
rect 37648 37204 37700 37213
rect 52828 37204 52880 37256
rect 38016 37136 38068 37188
rect 38384 37136 38436 37188
rect 38292 37068 38344 37120
rect 53564 37111 53616 37120
rect 53564 37077 53573 37111
rect 53573 37077 53607 37111
rect 53607 37077 53616 37111
rect 53564 37068 53616 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 17684 36864 17736 36916
rect 18144 36864 18196 36916
rect 19984 36864 20036 36916
rect 21640 36864 21692 36916
rect 21824 36864 21876 36916
rect 22560 36864 22612 36916
rect 17316 36728 17368 36780
rect 17592 36728 17644 36780
rect 18512 36796 18564 36848
rect 18328 36728 18380 36780
rect 19064 36728 19116 36780
rect 22376 36796 22428 36848
rect 21364 36728 21416 36780
rect 23020 36771 23072 36780
rect 23020 36737 23029 36771
rect 23029 36737 23063 36771
rect 23063 36737 23072 36771
rect 23020 36728 23072 36737
rect 24860 36864 24912 36916
rect 26148 36864 26200 36916
rect 29920 36864 29972 36916
rect 33968 36864 34020 36916
rect 20168 36660 20220 36712
rect 23664 36771 23716 36780
rect 23664 36737 23673 36771
rect 23673 36737 23707 36771
rect 23707 36737 23716 36771
rect 23664 36728 23716 36737
rect 23848 36771 23900 36780
rect 23848 36737 23857 36771
rect 23857 36737 23891 36771
rect 23891 36737 23900 36771
rect 23848 36728 23900 36737
rect 24308 36728 24360 36780
rect 24768 36728 24820 36780
rect 29552 36796 29604 36848
rect 30380 36839 30432 36848
rect 30380 36805 30389 36839
rect 30389 36805 30423 36839
rect 30423 36805 30432 36839
rect 30380 36796 30432 36805
rect 31116 36796 31168 36848
rect 33784 36796 33836 36848
rect 35072 36864 35124 36916
rect 37280 36864 37332 36916
rect 38200 36864 38252 36916
rect 23756 36660 23808 36712
rect 24032 36660 24084 36712
rect 18420 36592 18472 36644
rect 21088 36592 21140 36644
rect 21732 36592 21784 36644
rect 23940 36592 23992 36644
rect 25228 36660 25280 36712
rect 25412 36703 25464 36712
rect 25412 36669 25421 36703
rect 25421 36669 25455 36703
rect 25455 36669 25464 36703
rect 25412 36660 25464 36669
rect 26884 36728 26936 36780
rect 27068 36771 27120 36780
rect 27068 36737 27077 36771
rect 27077 36737 27111 36771
rect 27111 36737 27120 36771
rect 27068 36728 27120 36737
rect 27436 36728 27488 36780
rect 30840 36771 30892 36780
rect 30840 36737 30849 36771
rect 30849 36737 30883 36771
rect 30883 36737 30892 36771
rect 30840 36728 30892 36737
rect 31024 36771 31076 36780
rect 31024 36737 31033 36771
rect 31033 36737 31067 36771
rect 31067 36737 31076 36771
rect 31024 36728 31076 36737
rect 33416 36771 33468 36780
rect 33416 36737 33425 36771
rect 33425 36737 33459 36771
rect 33459 36737 33468 36771
rect 33416 36728 33468 36737
rect 34244 36728 34296 36780
rect 34796 36796 34848 36848
rect 35164 36771 35216 36780
rect 35164 36737 35173 36771
rect 35173 36737 35207 36771
rect 35207 36737 35216 36771
rect 35164 36728 35216 36737
rect 35532 36728 35584 36780
rect 37832 36728 37884 36780
rect 26516 36660 26568 36712
rect 27344 36660 27396 36712
rect 29184 36660 29236 36712
rect 31116 36660 31168 36712
rect 33692 36660 33744 36712
rect 33968 36660 34020 36712
rect 34704 36660 34756 36712
rect 36636 36703 36688 36712
rect 36636 36669 36645 36703
rect 36645 36669 36679 36703
rect 36679 36669 36688 36703
rect 36636 36660 36688 36669
rect 38016 36660 38068 36712
rect 38752 36728 38804 36780
rect 26240 36592 26292 36644
rect 26976 36592 27028 36644
rect 18604 36567 18656 36576
rect 18604 36533 18613 36567
rect 18613 36533 18647 36567
rect 18647 36533 18656 36567
rect 18604 36524 18656 36533
rect 19248 36524 19300 36576
rect 22284 36524 22336 36576
rect 24768 36524 24820 36576
rect 25872 36567 25924 36576
rect 25872 36533 25881 36567
rect 25881 36533 25915 36567
rect 25915 36533 25924 36567
rect 25872 36524 25924 36533
rect 26332 36567 26384 36576
rect 26332 36533 26341 36567
rect 26341 36533 26375 36567
rect 26375 36533 26384 36567
rect 26332 36524 26384 36533
rect 27160 36567 27212 36576
rect 27160 36533 27169 36567
rect 27169 36533 27203 36567
rect 27203 36533 27212 36567
rect 27160 36524 27212 36533
rect 30656 36524 30708 36576
rect 31760 36524 31812 36576
rect 32036 36524 32088 36576
rect 33140 36592 33192 36644
rect 33508 36592 33560 36644
rect 33784 36592 33836 36644
rect 39028 36660 39080 36712
rect 33324 36524 33376 36576
rect 33968 36524 34020 36576
rect 34152 36524 34204 36576
rect 35164 36524 35216 36576
rect 35348 36567 35400 36576
rect 35348 36533 35357 36567
rect 35357 36533 35391 36567
rect 35391 36533 35400 36567
rect 35348 36524 35400 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 21088 36320 21140 36372
rect 23020 36320 23072 36372
rect 25412 36320 25464 36372
rect 28540 36320 28592 36372
rect 17592 36252 17644 36304
rect 17960 36295 18012 36304
rect 17960 36261 17969 36295
rect 17969 36261 18003 36295
rect 18003 36261 18012 36295
rect 17960 36252 18012 36261
rect 18236 36252 18288 36304
rect 18144 36184 18196 36236
rect 17316 36116 17368 36168
rect 18052 36159 18104 36168
rect 18052 36125 18061 36159
rect 18061 36125 18095 36159
rect 18095 36125 18104 36159
rect 18236 36159 18288 36168
rect 18052 36116 18104 36125
rect 18236 36125 18245 36159
rect 18245 36125 18279 36159
rect 18279 36125 18288 36159
rect 18236 36116 18288 36125
rect 18512 36116 18564 36168
rect 20168 36184 20220 36236
rect 21916 36252 21968 36304
rect 29644 36295 29696 36304
rect 21640 36227 21692 36236
rect 21640 36193 21649 36227
rect 21649 36193 21683 36227
rect 21683 36193 21692 36227
rect 21640 36184 21692 36193
rect 21456 36159 21508 36168
rect 1860 36091 1912 36100
rect 1860 36057 1869 36091
rect 1869 36057 1903 36091
rect 1903 36057 1912 36091
rect 1860 36048 1912 36057
rect 16396 36048 16448 36100
rect 18696 36048 18748 36100
rect 21456 36125 21465 36159
rect 21465 36125 21499 36159
rect 21499 36125 21508 36159
rect 21456 36116 21508 36125
rect 21732 36116 21784 36168
rect 29644 36261 29653 36295
rect 29653 36261 29687 36295
rect 29687 36261 29696 36295
rect 29644 36252 29696 36261
rect 30104 36252 30156 36304
rect 33692 36320 33744 36372
rect 25872 36184 25924 36236
rect 26976 36184 27028 36236
rect 28724 36227 28776 36236
rect 28724 36193 28733 36227
rect 28733 36193 28767 36227
rect 28767 36193 28776 36227
rect 28724 36184 28776 36193
rect 33048 36252 33100 36304
rect 33784 36252 33836 36304
rect 34612 36320 34664 36372
rect 38752 36363 38804 36372
rect 38752 36329 38761 36363
rect 38761 36329 38795 36363
rect 38795 36329 38804 36363
rect 38752 36320 38804 36329
rect 34888 36252 34940 36304
rect 24584 36159 24636 36168
rect 24584 36125 24593 36159
rect 24593 36125 24627 36159
rect 24627 36125 24636 36159
rect 24584 36116 24636 36125
rect 24768 36159 24820 36168
rect 24768 36125 24777 36159
rect 24777 36125 24811 36159
rect 24811 36125 24820 36159
rect 24768 36116 24820 36125
rect 15476 35980 15528 36032
rect 16948 35980 17000 36032
rect 17592 36023 17644 36032
rect 17592 35989 17601 36023
rect 17601 35989 17635 36023
rect 17635 35989 17644 36023
rect 17592 35980 17644 35989
rect 17960 35980 18012 36032
rect 21364 36048 21416 36100
rect 23664 36091 23716 36100
rect 23664 36057 23673 36091
rect 23673 36057 23707 36091
rect 23707 36057 23716 36091
rect 23664 36048 23716 36057
rect 23848 36091 23900 36100
rect 23848 36057 23857 36091
rect 23857 36057 23891 36091
rect 23891 36057 23900 36091
rect 26332 36116 26384 36168
rect 27712 36116 27764 36168
rect 29000 36159 29052 36168
rect 29000 36125 29009 36159
rect 29009 36125 29043 36159
rect 29043 36125 29052 36159
rect 29000 36116 29052 36125
rect 29552 36116 29604 36168
rect 30472 36116 30524 36168
rect 23848 36048 23900 36057
rect 26884 36048 26936 36100
rect 30196 36048 30248 36100
rect 30748 36159 30800 36168
rect 30748 36125 30757 36159
rect 30757 36125 30791 36159
rect 30791 36125 30800 36159
rect 30748 36116 30800 36125
rect 31116 36159 31168 36168
rect 30656 36048 30708 36100
rect 31116 36125 31125 36159
rect 31125 36125 31159 36159
rect 31159 36125 31168 36159
rect 31116 36116 31168 36125
rect 32864 36116 32916 36168
rect 33508 36116 33560 36168
rect 31944 36048 31996 36100
rect 33876 36227 33928 36236
rect 33876 36193 33885 36227
rect 33885 36193 33919 36227
rect 33919 36193 33928 36227
rect 33876 36184 33928 36193
rect 35164 36184 35216 36236
rect 34336 36116 34388 36168
rect 35532 36116 35584 36168
rect 35808 36184 35860 36236
rect 39028 36252 39080 36304
rect 38292 36227 38344 36236
rect 38292 36193 38301 36227
rect 38301 36193 38335 36227
rect 38335 36193 38344 36227
rect 38292 36184 38344 36193
rect 36176 36116 36228 36168
rect 37372 36116 37424 36168
rect 38752 36159 38804 36168
rect 19984 35980 20036 36032
rect 20904 35980 20956 36032
rect 21272 36023 21324 36032
rect 21272 35989 21281 36023
rect 21281 35989 21315 36023
rect 21315 35989 21324 36023
rect 21272 35980 21324 35989
rect 24032 35980 24084 36032
rect 29184 35980 29236 36032
rect 31576 36023 31628 36032
rect 31576 35989 31585 36023
rect 31585 35989 31619 36023
rect 31619 35989 31628 36023
rect 31576 35980 31628 35989
rect 31852 35980 31904 36032
rect 34888 36048 34940 36100
rect 34428 35980 34480 36032
rect 35992 36048 36044 36100
rect 37648 36048 37700 36100
rect 37832 36048 37884 36100
rect 38752 36125 38761 36159
rect 38761 36125 38795 36159
rect 38795 36125 38804 36159
rect 38752 36116 38804 36125
rect 39764 36048 39816 36100
rect 52368 35980 52420 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 1860 35776 1912 35828
rect 18052 35819 18104 35828
rect 18052 35785 18061 35819
rect 18061 35785 18095 35819
rect 18095 35785 18104 35819
rect 18052 35776 18104 35785
rect 18604 35776 18656 35828
rect 19248 35819 19300 35828
rect 19248 35785 19257 35819
rect 19257 35785 19291 35819
rect 19291 35785 19300 35819
rect 19248 35776 19300 35785
rect 19984 35819 20036 35828
rect 17960 35708 18012 35760
rect 18880 35640 18932 35692
rect 19984 35785 20009 35819
rect 20009 35785 20036 35819
rect 20168 35819 20220 35828
rect 19984 35776 20036 35785
rect 20168 35785 20177 35819
rect 20177 35785 20211 35819
rect 20211 35785 20220 35819
rect 20168 35776 20220 35785
rect 20628 35776 20680 35828
rect 18236 35572 18288 35624
rect 18696 35572 18748 35624
rect 19156 35572 19208 35624
rect 20628 35683 20680 35692
rect 20628 35649 20637 35683
rect 20637 35649 20671 35683
rect 20671 35649 20680 35683
rect 20628 35640 20680 35649
rect 20812 35683 20864 35692
rect 20812 35649 20821 35683
rect 20821 35649 20855 35683
rect 20855 35649 20864 35683
rect 20812 35640 20864 35649
rect 20904 35615 20956 35624
rect 20904 35581 20913 35615
rect 20913 35581 20947 35615
rect 20947 35581 20956 35615
rect 20904 35572 20956 35581
rect 25320 35776 25372 35828
rect 26240 35776 26292 35828
rect 31760 35776 31812 35828
rect 34336 35819 34388 35828
rect 21640 35640 21692 35692
rect 22744 35640 22796 35692
rect 27988 35708 28040 35760
rect 30380 35751 30432 35760
rect 30380 35717 30389 35751
rect 30389 35717 30423 35751
rect 30423 35717 30432 35751
rect 30380 35708 30432 35717
rect 30748 35708 30800 35760
rect 24124 35683 24176 35692
rect 24124 35649 24133 35683
rect 24133 35649 24167 35683
rect 24167 35649 24176 35683
rect 24124 35640 24176 35649
rect 24216 35640 24268 35692
rect 24768 35640 24820 35692
rect 27068 35640 27120 35692
rect 27436 35640 27488 35692
rect 32036 35640 32088 35692
rect 34336 35785 34345 35819
rect 34345 35785 34379 35819
rect 34379 35785 34388 35819
rect 34336 35776 34388 35785
rect 34704 35776 34756 35828
rect 36636 35776 36688 35828
rect 21088 35504 21140 35556
rect 21456 35572 21508 35624
rect 15936 35436 15988 35488
rect 16396 35436 16448 35488
rect 16856 35479 16908 35488
rect 16856 35445 16865 35479
rect 16865 35445 16899 35479
rect 16899 35445 16908 35479
rect 16856 35436 16908 35445
rect 18144 35436 18196 35488
rect 19248 35436 19300 35488
rect 20904 35436 20956 35488
rect 21180 35436 21232 35488
rect 21824 35436 21876 35488
rect 23388 35479 23440 35488
rect 23388 35445 23397 35479
rect 23397 35445 23431 35479
rect 23431 35445 23440 35479
rect 23388 35436 23440 35445
rect 23572 35436 23624 35488
rect 25044 35504 25096 35556
rect 26884 35572 26936 35624
rect 29552 35572 29604 35624
rect 33968 35640 34020 35692
rect 34152 35683 34204 35692
rect 34152 35649 34161 35683
rect 34161 35649 34195 35683
rect 34195 35649 34204 35683
rect 34152 35640 34204 35649
rect 35348 35708 35400 35760
rect 37740 35776 37792 35828
rect 39672 35776 39724 35828
rect 37464 35751 37516 35760
rect 37464 35717 37491 35751
rect 37491 35717 37516 35751
rect 37464 35708 37516 35717
rect 37648 35751 37700 35760
rect 37648 35717 37657 35751
rect 37657 35717 37691 35751
rect 37691 35717 37700 35751
rect 37648 35708 37700 35717
rect 38568 35708 38620 35760
rect 35072 35683 35124 35692
rect 35072 35649 35081 35683
rect 35081 35649 35115 35683
rect 35115 35649 35124 35683
rect 35072 35640 35124 35649
rect 36452 35683 36504 35692
rect 34612 35572 34664 35624
rect 35164 35615 35216 35624
rect 35164 35581 35173 35615
rect 35173 35581 35207 35615
rect 35207 35581 35216 35615
rect 35164 35572 35216 35581
rect 36452 35649 36461 35683
rect 36461 35649 36495 35683
rect 36495 35649 36504 35683
rect 36452 35640 36504 35649
rect 38292 35683 38344 35692
rect 38292 35649 38301 35683
rect 38301 35649 38335 35683
rect 38335 35649 38344 35683
rect 38292 35640 38344 35649
rect 38752 35683 38804 35692
rect 38752 35649 38761 35683
rect 38761 35649 38795 35683
rect 38795 35649 38804 35683
rect 38752 35640 38804 35649
rect 39764 35640 39816 35692
rect 27068 35504 27120 35556
rect 29000 35504 29052 35556
rect 30288 35504 30340 35556
rect 32128 35504 32180 35556
rect 32404 35504 32456 35556
rect 24584 35436 24636 35488
rect 29552 35436 29604 35488
rect 30932 35479 30984 35488
rect 30932 35445 30941 35479
rect 30941 35445 30975 35479
rect 30975 35445 30984 35479
rect 30932 35436 30984 35445
rect 32680 35436 32732 35488
rect 33232 35479 33284 35488
rect 33232 35445 33241 35479
rect 33241 35445 33275 35479
rect 33275 35445 33284 35479
rect 33232 35436 33284 35445
rect 34060 35436 34112 35488
rect 36176 35572 36228 35624
rect 37740 35436 37792 35488
rect 38384 35436 38436 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 18236 35232 18288 35284
rect 20628 35232 20680 35284
rect 20904 35232 20956 35284
rect 21088 35232 21140 35284
rect 21272 35232 21324 35284
rect 23388 35232 23440 35284
rect 23848 35232 23900 35284
rect 24400 35232 24452 35284
rect 24768 35275 24820 35284
rect 24768 35241 24777 35275
rect 24777 35241 24811 35275
rect 24811 35241 24820 35275
rect 24768 35232 24820 35241
rect 28356 35232 28408 35284
rect 16948 35096 17000 35148
rect 19064 35164 19116 35216
rect 16764 35028 16816 35080
rect 17408 35096 17460 35148
rect 17868 35096 17920 35148
rect 17960 35139 18012 35148
rect 17960 35105 17969 35139
rect 17969 35105 18003 35139
rect 18003 35105 18012 35139
rect 17960 35096 18012 35105
rect 17592 35028 17644 35080
rect 18052 35071 18104 35080
rect 18052 35037 18061 35071
rect 18061 35037 18095 35071
rect 18095 35037 18104 35071
rect 18052 35028 18104 35037
rect 18512 35071 18564 35080
rect 18512 35037 18521 35071
rect 18521 35037 18555 35071
rect 18555 35037 18564 35071
rect 18512 35028 18564 35037
rect 19248 35096 19300 35148
rect 19432 35071 19484 35080
rect 19432 35037 19441 35071
rect 19441 35037 19475 35071
rect 19475 35037 19484 35071
rect 19432 35028 19484 35037
rect 20720 35096 20772 35148
rect 19984 35028 20036 35080
rect 20628 35028 20680 35080
rect 21916 35096 21968 35148
rect 22744 35139 22796 35148
rect 22744 35105 22753 35139
rect 22753 35105 22787 35139
rect 22787 35105 22796 35139
rect 22744 35096 22796 35105
rect 24124 35164 24176 35216
rect 25872 35164 25924 35216
rect 22560 35071 22612 35080
rect 19340 34960 19392 35012
rect 21272 35003 21324 35012
rect 15936 34892 15988 34944
rect 19156 34892 19208 34944
rect 21272 34969 21281 35003
rect 21281 34969 21315 35003
rect 21315 34969 21324 35003
rect 22560 35037 22569 35071
rect 22569 35037 22603 35071
rect 22603 35037 22612 35071
rect 22560 35028 22612 35037
rect 22928 35071 22980 35080
rect 22928 35037 22937 35071
rect 22937 35037 22971 35071
rect 22971 35037 22980 35071
rect 22928 35028 22980 35037
rect 23848 35028 23900 35080
rect 26976 35096 27028 35148
rect 31300 35232 31352 35284
rect 35808 35232 35860 35284
rect 37464 35275 37516 35284
rect 37464 35241 37473 35275
rect 37473 35241 37507 35275
rect 37507 35241 37516 35275
rect 37464 35232 37516 35241
rect 29092 35164 29144 35216
rect 33416 35164 33468 35216
rect 29184 35096 29236 35148
rect 27160 35028 27212 35080
rect 21272 34960 21324 34969
rect 25044 34960 25096 35012
rect 29644 35003 29696 35012
rect 29644 34969 29653 35003
rect 29653 34969 29687 35003
rect 29687 34969 29696 35003
rect 29644 34960 29696 34969
rect 31852 35028 31904 35080
rect 32128 35028 32180 35080
rect 32680 35071 32732 35080
rect 32680 35037 32714 35071
rect 32714 35037 32732 35071
rect 32680 35028 32732 35037
rect 36084 35096 36136 35148
rect 34612 35028 34664 35080
rect 34796 35028 34848 35080
rect 35348 35028 35400 35080
rect 35532 35028 35584 35080
rect 36544 35164 36596 35216
rect 39764 35232 39816 35284
rect 37832 35071 37884 35080
rect 37832 35037 37841 35071
rect 37841 35037 37875 35071
rect 37875 35037 37884 35071
rect 37832 35028 37884 35037
rect 20076 34935 20128 34944
rect 20076 34901 20085 34935
rect 20085 34901 20119 34935
rect 20119 34901 20128 34935
rect 20076 34892 20128 34901
rect 25780 34892 25832 34944
rect 27712 34892 27764 34944
rect 29552 34892 29604 34944
rect 30564 34935 30616 34944
rect 30564 34901 30573 34935
rect 30573 34901 30607 34935
rect 30607 34901 30616 34935
rect 30564 34892 30616 34901
rect 31392 34892 31444 34944
rect 31668 34892 31720 34944
rect 33232 34892 33284 34944
rect 34336 34892 34388 34944
rect 36452 34960 36504 35012
rect 37648 35003 37700 35012
rect 37648 34969 37657 35003
rect 37657 34969 37691 35003
rect 37691 34969 37700 35003
rect 37648 34960 37700 34969
rect 53564 35003 53616 35012
rect 53564 34969 53573 35003
rect 53573 34969 53607 35003
rect 53607 34969 53616 35003
rect 53564 34960 53616 34969
rect 35348 34892 35400 34944
rect 36636 34892 36688 34944
rect 38844 34935 38896 34944
rect 38844 34901 38853 34935
rect 38853 34901 38887 34935
rect 38887 34901 38896 34935
rect 38844 34892 38896 34901
rect 52460 34892 52512 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 15476 34731 15528 34740
rect 15476 34697 15485 34731
rect 15485 34697 15519 34731
rect 15519 34697 15528 34731
rect 15476 34688 15528 34697
rect 16948 34688 17000 34740
rect 18512 34688 18564 34740
rect 18880 34731 18932 34740
rect 18880 34697 18889 34731
rect 18889 34697 18923 34731
rect 18923 34697 18932 34731
rect 18880 34688 18932 34697
rect 22560 34688 22612 34740
rect 22928 34688 22980 34740
rect 25320 34688 25372 34740
rect 26424 34731 26476 34740
rect 26424 34697 26433 34731
rect 26433 34697 26467 34731
rect 26467 34697 26476 34731
rect 26424 34688 26476 34697
rect 27160 34688 27212 34740
rect 30748 34731 30800 34740
rect 30748 34697 30757 34731
rect 30757 34697 30791 34731
rect 30791 34697 30800 34731
rect 30748 34688 30800 34697
rect 32404 34688 32456 34740
rect 16856 34620 16908 34672
rect 1584 34552 1636 34604
rect 18052 34620 18104 34672
rect 19064 34663 19116 34672
rect 19064 34629 19073 34663
rect 19073 34629 19107 34663
rect 19107 34629 19116 34663
rect 19064 34620 19116 34629
rect 22284 34620 22336 34672
rect 23664 34620 23716 34672
rect 25044 34620 25096 34672
rect 25872 34620 25924 34672
rect 30472 34620 30524 34672
rect 31392 34663 31444 34672
rect 31392 34629 31401 34663
rect 31401 34629 31435 34663
rect 31435 34629 31444 34663
rect 31392 34620 31444 34629
rect 17592 34552 17644 34604
rect 18236 34595 18288 34604
rect 18236 34561 18245 34595
rect 18245 34561 18279 34595
rect 18279 34561 18288 34595
rect 18236 34552 18288 34561
rect 2044 34527 2096 34536
rect 2044 34493 2053 34527
rect 2053 34493 2087 34527
rect 2087 34493 2096 34527
rect 2044 34484 2096 34493
rect 16764 34484 16816 34536
rect 19432 34552 19484 34604
rect 20628 34552 20680 34604
rect 21088 34595 21140 34604
rect 21088 34561 21097 34595
rect 21097 34561 21131 34595
rect 21131 34561 21140 34595
rect 21088 34552 21140 34561
rect 18420 34527 18472 34536
rect 18420 34493 18429 34527
rect 18429 34493 18463 34527
rect 18463 34493 18472 34527
rect 18420 34484 18472 34493
rect 19340 34484 19392 34536
rect 19800 34527 19852 34536
rect 19800 34493 19809 34527
rect 19809 34493 19843 34527
rect 19843 34493 19852 34527
rect 19800 34484 19852 34493
rect 21272 34527 21324 34536
rect 21272 34493 21281 34527
rect 21281 34493 21315 34527
rect 21315 34493 21324 34527
rect 21272 34484 21324 34493
rect 15476 34416 15528 34468
rect 16396 34416 16448 34468
rect 24676 34552 24728 34604
rect 24860 34552 24912 34604
rect 25504 34595 25556 34604
rect 25504 34561 25513 34595
rect 25513 34561 25547 34595
rect 25547 34561 25556 34595
rect 25504 34552 25556 34561
rect 25780 34595 25832 34604
rect 22008 34416 22060 34468
rect 25780 34561 25789 34595
rect 25789 34561 25823 34595
rect 25823 34561 25832 34595
rect 25780 34552 25832 34561
rect 26884 34552 26936 34604
rect 28816 34595 28868 34604
rect 26056 34484 26108 34536
rect 28816 34561 28825 34595
rect 28825 34561 28859 34595
rect 28859 34561 28868 34595
rect 28816 34552 28868 34561
rect 29092 34595 29144 34604
rect 29092 34561 29101 34595
rect 29101 34561 29135 34595
rect 29135 34561 29144 34595
rect 29092 34552 29144 34561
rect 29000 34527 29052 34536
rect 29000 34493 29009 34527
rect 29009 34493 29043 34527
rect 29043 34493 29052 34527
rect 30288 34552 30340 34604
rect 30656 34595 30708 34604
rect 30656 34561 30665 34595
rect 30665 34561 30699 34595
rect 30699 34561 30708 34595
rect 30656 34552 30708 34561
rect 31300 34595 31352 34604
rect 29000 34484 29052 34493
rect 29920 34527 29972 34536
rect 29920 34493 29929 34527
rect 29929 34493 29963 34527
rect 29963 34493 29972 34527
rect 30196 34527 30248 34536
rect 29920 34484 29972 34493
rect 30196 34493 30205 34527
rect 30205 34493 30239 34527
rect 30239 34493 30248 34527
rect 30196 34484 30248 34493
rect 31300 34561 31309 34595
rect 31309 34561 31343 34595
rect 31343 34561 31352 34595
rect 31300 34552 31352 34561
rect 32404 34595 32456 34604
rect 32404 34561 32413 34595
rect 32413 34561 32447 34595
rect 32447 34561 32456 34595
rect 32404 34552 32456 34561
rect 36544 34731 36596 34740
rect 36544 34697 36553 34731
rect 36553 34697 36587 34731
rect 36587 34697 36596 34731
rect 36544 34688 36596 34697
rect 38292 34688 38344 34740
rect 33048 34620 33100 34672
rect 32588 34595 32640 34604
rect 32588 34561 32597 34595
rect 32597 34561 32631 34595
rect 32631 34561 32640 34595
rect 32588 34552 32640 34561
rect 17408 34391 17460 34400
rect 17408 34357 17417 34391
rect 17417 34357 17451 34391
rect 17451 34357 17460 34391
rect 17408 34348 17460 34357
rect 18144 34348 18196 34400
rect 22652 34348 22704 34400
rect 24676 34391 24728 34400
rect 24676 34357 24685 34391
rect 24685 34357 24719 34391
rect 24719 34357 24728 34391
rect 24676 34348 24728 34357
rect 27344 34416 27396 34468
rect 29828 34416 29880 34468
rect 30104 34416 30156 34468
rect 32864 34552 32916 34604
rect 34336 34620 34388 34672
rect 34612 34620 34664 34672
rect 34796 34552 34848 34604
rect 35348 34595 35400 34604
rect 35348 34561 35357 34595
rect 35357 34561 35391 34595
rect 35391 34561 35400 34595
rect 35348 34552 35400 34561
rect 35808 34595 35860 34604
rect 35808 34561 35817 34595
rect 35817 34561 35851 34595
rect 35851 34561 35860 34595
rect 35808 34552 35860 34561
rect 35992 34595 36044 34604
rect 35992 34561 36001 34595
rect 36001 34561 36035 34595
rect 36035 34561 36044 34595
rect 35992 34552 36044 34561
rect 36452 34552 36504 34604
rect 37648 34552 37700 34604
rect 39672 34688 39724 34740
rect 34704 34484 34756 34536
rect 27436 34348 27488 34400
rect 28172 34391 28224 34400
rect 28172 34357 28181 34391
rect 28181 34357 28215 34391
rect 28215 34357 28224 34391
rect 28172 34348 28224 34357
rect 31300 34348 31352 34400
rect 32404 34348 32456 34400
rect 33232 34391 33284 34400
rect 33232 34357 33241 34391
rect 33241 34357 33275 34391
rect 33275 34357 33284 34391
rect 33232 34348 33284 34357
rect 33416 34391 33468 34400
rect 33416 34357 33425 34391
rect 33425 34357 33459 34391
rect 33459 34357 33468 34391
rect 33416 34348 33468 34357
rect 35900 34391 35952 34400
rect 35900 34357 35909 34391
rect 35909 34357 35943 34391
rect 35943 34357 35952 34391
rect 35900 34348 35952 34357
rect 38016 34391 38068 34400
rect 38016 34357 38025 34391
rect 38025 34357 38059 34391
rect 38059 34357 38068 34391
rect 38844 34484 38896 34536
rect 39672 34484 39724 34536
rect 50712 34484 50764 34536
rect 38016 34348 38068 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 16856 34144 16908 34196
rect 1584 34119 1636 34128
rect 1584 34085 1593 34119
rect 1593 34085 1627 34119
rect 1627 34085 1636 34119
rect 1584 34076 1636 34085
rect 18052 34144 18104 34196
rect 19432 34144 19484 34196
rect 19800 34144 19852 34196
rect 20812 34144 20864 34196
rect 25504 34187 25556 34196
rect 25504 34153 25513 34187
rect 25513 34153 25547 34187
rect 25547 34153 25556 34187
rect 25504 34144 25556 34153
rect 26056 34187 26108 34196
rect 26056 34153 26065 34187
rect 26065 34153 26099 34187
rect 26099 34153 26108 34187
rect 26056 34144 26108 34153
rect 26240 34187 26292 34196
rect 26240 34153 26249 34187
rect 26249 34153 26283 34187
rect 26283 34153 26292 34187
rect 26240 34144 26292 34153
rect 26884 34187 26936 34196
rect 26884 34153 26893 34187
rect 26893 34153 26927 34187
rect 26927 34153 26936 34187
rect 26884 34144 26936 34153
rect 29920 34144 29972 34196
rect 32588 34144 32640 34196
rect 32680 34187 32732 34196
rect 32680 34153 32689 34187
rect 32689 34153 32723 34187
rect 32723 34153 32732 34187
rect 32680 34144 32732 34153
rect 18420 34076 18472 34128
rect 22192 34076 22244 34128
rect 24860 34076 24912 34128
rect 18236 34008 18288 34060
rect 20076 34051 20128 34060
rect 20076 34017 20085 34051
rect 20085 34017 20119 34051
rect 20119 34017 20128 34051
rect 20076 34008 20128 34017
rect 23572 34051 23624 34060
rect 18144 33983 18196 33992
rect 18144 33949 18153 33983
rect 18153 33949 18187 33983
rect 18187 33949 18196 33983
rect 18144 33940 18196 33949
rect 19432 33940 19484 33992
rect 22008 33983 22060 33992
rect 22008 33949 22017 33983
rect 22017 33949 22051 33983
rect 22051 33949 22060 33983
rect 22008 33940 22060 33949
rect 22192 33983 22244 33992
rect 22192 33949 22201 33983
rect 22201 33949 22235 33983
rect 22235 33949 22244 33983
rect 22192 33940 22244 33949
rect 22652 33983 22704 33992
rect 22652 33949 22661 33983
rect 22661 33949 22695 33983
rect 22695 33949 22704 33983
rect 22652 33940 22704 33949
rect 23572 34017 23581 34051
rect 23581 34017 23615 34051
rect 23615 34017 23624 34051
rect 23572 34008 23624 34017
rect 24676 34008 24728 34060
rect 26424 34076 26476 34128
rect 23296 33940 23348 33992
rect 18328 33915 18380 33924
rect 18328 33881 18337 33915
rect 18337 33881 18371 33915
rect 18371 33881 18380 33915
rect 18328 33872 18380 33881
rect 23756 33940 23808 33992
rect 16764 33804 16816 33856
rect 21456 33847 21508 33856
rect 21456 33813 21465 33847
rect 21465 33813 21499 33847
rect 21499 33813 21508 33847
rect 21456 33804 21508 33813
rect 24492 33847 24544 33856
rect 24492 33813 24501 33847
rect 24501 33813 24535 33847
rect 24535 33813 24544 33847
rect 24492 33804 24544 33813
rect 26240 33940 26292 33992
rect 27068 33940 27120 33992
rect 28816 34076 28868 34128
rect 29000 34076 29052 34128
rect 29276 34076 29328 34128
rect 29736 34076 29788 34128
rect 28264 34008 28316 34060
rect 28356 34008 28408 34060
rect 26424 33915 26476 33924
rect 26424 33881 26433 33915
rect 26433 33881 26467 33915
rect 26467 33881 26476 33915
rect 26424 33872 26476 33881
rect 28172 33940 28224 33992
rect 29092 34008 29144 34060
rect 29552 34008 29604 34060
rect 29828 34051 29880 34060
rect 29828 34017 29837 34051
rect 29837 34017 29871 34051
rect 29871 34017 29880 34051
rect 29828 34008 29880 34017
rect 28816 33940 28868 33992
rect 29736 33983 29788 33992
rect 29736 33949 29745 33983
rect 29745 33949 29779 33983
rect 29779 33949 29788 33983
rect 29736 33940 29788 33949
rect 30104 33940 30156 33992
rect 31392 34008 31444 34060
rect 31300 33983 31352 33992
rect 31300 33949 31309 33983
rect 31309 33949 31343 33983
rect 31343 33949 31352 33983
rect 32772 33983 32824 33992
rect 31300 33940 31352 33949
rect 32772 33949 32781 33983
rect 32781 33949 32815 33983
rect 32815 33949 32824 33983
rect 32772 33940 32824 33949
rect 33232 33940 33284 33992
rect 35348 34144 35400 34196
rect 36544 34187 36596 34196
rect 36544 34153 36553 34187
rect 36553 34153 36587 34187
rect 36587 34153 36596 34187
rect 36544 34144 36596 34153
rect 34704 34076 34756 34128
rect 35900 34008 35952 34060
rect 34612 33940 34664 33992
rect 35348 33940 35400 33992
rect 35532 33940 35584 33992
rect 27160 33804 27212 33856
rect 27252 33804 27304 33856
rect 35992 33872 36044 33924
rect 38936 33940 38988 33992
rect 53656 33940 53708 33992
rect 38016 33872 38068 33924
rect 30380 33804 30432 33856
rect 30472 33804 30524 33856
rect 31576 33804 31628 33856
rect 32588 33804 32640 33856
rect 32864 33804 32916 33856
rect 34336 33804 34388 33856
rect 35716 33847 35768 33856
rect 35716 33813 35725 33847
rect 35725 33813 35759 33847
rect 35759 33813 35768 33847
rect 35716 33804 35768 33813
rect 37648 33847 37700 33856
rect 37648 33813 37657 33847
rect 37657 33813 37691 33847
rect 37691 33813 37700 33847
rect 37648 33804 37700 33813
rect 38200 33847 38252 33856
rect 38200 33813 38209 33847
rect 38209 33813 38243 33847
rect 38243 33813 38252 33847
rect 38200 33804 38252 33813
rect 40408 33804 40460 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 18328 33600 18380 33652
rect 18972 33643 19024 33652
rect 18972 33609 18981 33643
rect 18981 33609 19015 33643
rect 19015 33609 19024 33643
rect 18972 33600 19024 33609
rect 24676 33643 24728 33652
rect 24676 33609 24685 33643
rect 24685 33609 24719 33643
rect 24719 33609 24728 33643
rect 24676 33600 24728 33609
rect 26516 33600 26568 33652
rect 16396 33464 16448 33516
rect 21916 33532 21968 33584
rect 24492 33532 24544 33584
rect 26240 33532 26292 33584
rect 18236 33464 18288 33516
rect 22560 33464 22612 33516
rect 22652 33507 22704 33516
rect 22652 33473 22661 33507
rect 22661 33473 22695 33507
rect 22695 33473 22704 33507
rect 23296 33507 23348 33516
rect 22652 33464 22704 33473
rect 23296 33473 23305 33507
rect 23305 33473 23339 33507
rect 23339 33473 23348 33507
rect 23296 33464 23348 33473
rect 23388 33464 23440 33516
rect 27252 33507 27304 33516
rect 27252 33473 27261 33507
rect 27261 33473 27295 33507
rect 27295 33473 27304 33507
rect 29276 33600 29328 33652
rect 29644 33600 29696 33652
rect 29736 33600 29788 33652
rect 32680 33600 32732 33652
rect 33324 33600 33376 33652
rect 34704 33600 34756 33652
rect 34796 33600 34848 33652
rect 35256 33600 35308 33652
rect 35532 33600 35584 33652
rect 35992 33600 36044 33652
rect 28264 33532 28316 33584
rect 30472 33575 30524 33584
rect 27252 33464 27304 33473
rect 21272 33396 21324 33448
rect 23756 33396 23808 33448
rect 27436 33439 27488 33448
rect 27436 33405 27445 33439
rect 27445 33405 27479 33439
rect 27479 33405 27488 33439
rect 27436 33396 27488 33405
rect 21364 33328 21416 33380
rect 24492 33328 24544 33380
rect 19340 33260 19392 33312
rect 20812 33260 20864 33312
rect 21456 33260 21508 33312
rect 23112 33303 23164 33312
rect 23112 33269 23121 33303
rect 23121 33269 23155 33303
rect 23155 33269 23164 33303
rect 23112 33260 23164 33269
rect 23572 33260 23624 33312
rect 23848 33260 23900 33312
rect 25780 33303 25832 33312
rect 25780 33269 25789 33303
rect 25789 33269 25823 33303
rect 25823 33269 25832 33303
rect 25780 33260 25832 33269
rect 26424 33260 26476 33312
rect 28724 33507 28776 33516
rect 28724 33473 28733 33507
rect 28733 33473 28767 33507
rect 28767 33473 28776 33507
rect 28724 33464 28776 33473
rect 29092 33464 29144 33516
rect 29368 33396 29420 33448
rect 29000 33328 29052 33380
rect 29184 33328 29236 33380
rect 29920 33464 29972 33516
rect 30472 33541 30481 33575
rect 30481 33541 30515 33575
rect 30515 33541 30524 33575
rect 30472 33532 30524 33541
rect 31392 33532 31444 33584
rect 33048 33532 33100 33584
rect 34520 33532 34572 33584
rect 35624 33532 35676 33584
rect 30104 33396 30156 33448
rect 32496 33396 32548 33448
rect 32588 33396 32640 33448
rect 33416 33464 33468 33516
rect 35256 33507 35308 33516
rect 32864 33396 32916 33448
rect 34336 33439 34388 33448
rect 29920 33328 29972 33380
rect 33324 33328 33376 33380
rect 34060 33371 34112 33380
rect 34060 33337 34069 33371
rect 34069 33337 34103 33371
rect 34103 33337 34112 33371
rect 34060 33328 34112 33337
rect 34336 33405 34345 33439
rect 34345 33405 34379 33439
rect 34379 33405 34388 33439
rect 34336 33396 34388 33405
rect 35256 33473 35265 33507
rect 35265 33473 35299 33507
rect 35299 33473 35308 33507
rect 35256 33464 35308 33473
rect 36544 33532 36596 33584
rect 36084 33507 36136 33516
rect 36084 33473 36093 33507
rect 36093 33473 36127 33507
rect 36127 33473 36136 33507
rect 36084 33464 36136 33473
rect 36176 33464 36228 33516
rect 38200 33532 38252 33584
rect 37464 33507 37516 33516
rect 37464 33473 37473 33507
rect 37473 33473 37507 33507
rect 37507 33473 37516 33507
rect 37464 33464 37516 33473
rect 35900 33396 35952 33448
rect 37372 33439 37424 33448
rect 37372 33405 37381 33439
rect 37381 33405 37415 33439
rect 37415 33405 37424 33439
rect 37372 33396 37424 33405
rect 38752 33396 38804 33448
rect 40408 33328 40460 33380
rect 30840 33303 30892 33312
rect 30840 33269 30849 33303
rect 30849 33269 30883 33303
rect 30883 33269 30892 33303
rect 30840 33260 30892 33269
rect 32404 33260 32456 33312
rect 53104 33260 53156 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 2044 33056 2096 33108
rect 17960 33056 18012 33108
rect 26240 32988 26292 33040
rect 28264 32988 28316 33040
rect 29092 32988 29144 33040
rect 30748 32988 30800 33040
rect 33692 33056 33744 33108
rect 35348 33099 35400 33108
rect 35348 33065 35357 33099
rect 35357 33065 35391 33099
rect 35391 33065 35400 33099
rect 35348 33056 35400 33065
rect 36084 33056 36136 33108
rect 38292 33056 38344 33108
rect 38936 33099 38988 33108
rect 38936 33065 38945 33099
rect 38945 33065 38979 33099
rect 38979 33065 38988 33099
rect 38936 33056 38988 33065
rect 18420 32920 18472 32972
rect 18972 32920 19024 32972
rect 17960 32852 18012 32904
rect 18512 32852 18564 32904
rect 18604 32852 18656 32904
rect 20076 32895 20128 32904
rect 20076 32861 20085 32895
rect 20085 32861 20119 32895
rect 20119 32861 20128 32895
rect 20076 32852 20128 32861
rect 20260 32895 20312 32904
rect 20260 32861 20269 32895
rect 20269 32861 20303 32895
rect 20303 32861 20312 32895
rect 20260 32852 20312 32861
rect 23296 32920 23348 32972
rect 24492 32963 24544 32972
rect 24492 32929 24501 32963
rect 24501 32929 24535 32963
rect 24535 32929 24544 32963
rect 24492 32920 24544 32929
rect 21456 32852 21508 32904
rect 22008 32852 22060 32904
rect 22560 32852 22612 32904
rect 23204 32852 23256 32904
rect 25596 32895 25648 32904
rect 21916 32827 21968 32836
rect 21916 32793 21925 32827
rect 21925 32793 21959 32827
rect 21959 32793 21968 32827
rect 21916 32784 21968 32793
rect 25596 32861 25605 32895
rect 25605 32861 25639 32895
rect 25639 32861 25648 32895
rect 25596 32852 25648 32861
rect 26424 32920 26476 32972
rect 25780 32895 25832 32904
rect 25780 32861 25789 32895
rect 25789 32861 25823 32895
rect 25823 32861 25832 32895
rect 25780 32852 25832 32861
rect 26516 32852 26568 32904
rect 26976 32852 27028 32904
rect 28724 32852 28776 32904
rect 29552 32920 29604 32972
rect 29920 32920 29972 32972
rect 30840 32852 30892 32904
rect 31392 32920 31444 32972
rect 31668 32920 31720 32972
rect 31208 32852 31260 32904
rect 31576 32852 31628 32904
rect 32496 32920 32548 32972
rect 34244 32920 34296 32972
rect 38016 32988 38068 33040
rect 29644 32784 29696 32836
rect 16856 32759 16908 32768
rect 16856 32725 16865 32759
rect 16865 32725 16899 32759
rect 16899 32725 16908 32759
rect 16856 32716 16908 32725
rect 18144 32716 18196 32768
rect 18328 32759 18380 32768
rect 18328 32725 18337 32759
rect 18337 32725 18371 32759
rect 18371 32725 18380 32759
rect 18328 32716 18380 32725
rect 19248 32716 19300 32768
rect 19432 32716 19484 32768
rect 20720 32716 20772 32768
rect 21364 32759 21416 32768
rect 21364 32725 21373 32759
rect 21373 32725 21407 32759
rect 21407 32725 21416 32759
rect 21364 32716 21416 32725
rect 22652 32716 22704 32768
rect 23020 32716 23072 32768
rect 23296 32759 23348 32768
rect 23296 32725 23305 32759
rect 23305 32725 23339 32759
rect 23339 32725 23348 32759
rect 23296 32716 23348 32725
rect 23940 32716 23992 32768
rect 25504 32716 25556 32768
rect 25780 32716 25832 32768
rect 30288 32716 30340 32768
rect 30380 32716 30432 32768
rect 30932 32759 30984 32768
rect 30932 32725 30941 32759
rect 30941 32725 30975 32759
rect 30975 32725 30984 32759
rect 30932 32716 30984 32725
rect 31944 32784 31996 32836
rect 32864 32784 32916 32836
rect 33508 32852 33560 32904
rect 35072 32895 35124 32904
rect 35072 32861 35081 32895
rect 35081 32861 35115 32895
rect 35115 32861 35124 32895
rect 35072 32852 35124 32861
rect 35716 32852 35768 32904
rect 37648 32920 37700 32972
rect 35532 32784 35584 32836
rect 38016 32784 38068 32836
rect 38660 32784 38712 32836
rect 35716 32716 35768 32768
rect 36636 32716 36688 32768
rect 36728 32759 36780 32768
rect 36728 32725 36737 32759
rect 36737 32725 36771 32759
rect 36771 32725 36780 32759
rect 36728 32716 36780 32725
rect 38200 32716 38252 32768
rect 40408 32759 40460 32768
rect 40408 32725 40417 32759
rect 40417 32725 40451 32759
rect 40451 32725 40460 32759
rect 40408 32716 40460 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 16028 32376 16080 32428
rect 18052 32512 18104 32564
rect 17684 32444 17736 32496
rect 18604 32512 18656 32564
rect 20260 32512 20312 32564
rect 25596 32555 25648 32564
rect 25596 32521 25605 32555
rect 25605 32521 25639 32555
rect 25639 32521 25648 32555
rect 25596 32512 25648 32521
rect 27344 32512 27396 32564
rect 28448 32555 28500 32564
rect 28448 32521 28457 32555
rect 28457 32521 28491 32555
rect 28491 32521 28500 32555
rect 28448 32512 28500 32521
rect 28724 32512 28776 32564
rect 29644 32555 29696 32564
rect 29644 32521 29653 32555
rect 29653 32521 29687 32555
rect 29687 32521 29696 32555
rect 29644 32512 29696 32521
rect 31484 32512 31536 32564
rect 33140 32512 33192 32564
rect 33324 32512 33376 32564
rect 18972 32487 19024 32496
rect 18972 32453 18981 32487
rect 18981 32453 19015 32487
rect 19015 32453 19024 32487
rect 18972 32444 19024 32453
rect 19248 32444 19300 32496
rect 17684 32351 17736 32360
rect 17684 32317 17693 32351
rect 17693 32317 17727 32351
rect 17727 32317 17736 32351
rect 18052 32376 18104 32428
rect 18420 32419 18472 32428
rect 18420 32385 18429 32419
rect 18429 32385 18463 32419
rect 18463 32385 18472 32419
rect 22008 32444 22060 32496
rect 18420 32376 18472 32385
rect 19524 32376 19576 32428
rect 20812 32419 20864 32428
rect 20812 32385 20821 32419
rect 20821 32385 20855 32419
rect 20855 32385 20864 32419
rect 20812 32376 20864 32385
rect 21916 32419 21968 32428
rect 21916 32385 21925 32419
rect 21925 32385 21959 32419
rect 21959 32385 21968 32419
rect 21916 32376 21968 32385
rect 23756 32444 23808 32496
rect 22560 32419 22612 32428
rect 22560 32385 22569 32419
rect 22569 32385 22603 32419
rect 22603 32385 22612 32419
rect 22560 32376 22612 32385
rect 23112 32376 23164 32428
rect 23204 32419 23256 32428
rect 23204 32385 23213 32419
rect 23213 32385 23247 32419
rect 23247 32385 23256 32419
rect 23204 32376 23256 32385
rect 23664 32376 23716 32428
rect 24400 32419 24452 32428
rect 24400 32385 24409 32419
rect 24409 32385 24443 32419
rect 24443 32385 24452 32419
rect 24400 32376 24452 32385
rect 25320 32444 25372 32496
rect 25504 32419 25556 32428
rect 25504 32385 25513 32419
rect 25513 32385 25547 32419
rect 25547 32385 25556 32419
rect 25504 32376 25556 32385
rect 30104 32444 30156 32496
rect 30840 32444 30892 32496
rect 33600 32444 33652 32496
rect 34152 32512 34204 32564
rect 35808 32555 35860 32564
rect 35808 32521 35817 32555
rect 35817 32521 35851 32555
rect 35851 32521 35860 32555
rect 35808 32512 35860 32521
rect 37464 32512 37516 32564
rect 38200 32555 38252 32564
rect 38200 32521 38209 32555
rect 38209 32521 38243 32555
rect 38243 32521 38252 32555
rect 38200 32512 38252 32521
rect 38660 32555 38712 32564
rect 38660 32521 38669 32555
rect 38669 32521 38703 32555
rect 38703 32521 38712 32555
rect 38660 32512 38712 32521
rect 35072 32444 35124 32496
rect 29552 32419 29604 32428
rect 29552 32385 29561 32419
rect 29561 32385 29595 32419
rect 29595 32385 29604 32419
rect 29552 32376 29604 32385
rect 29736 32419 29788 32428
rect 29736 32385 29745 32419
rect 29745 32385 29779 32419
rect 29779 32385 29788 32419
rect 29736 32376 29788 32385
rect 20720 32351 20772 32360
rect 17684 32308 17736 32317
rect 20720 32317 20729 32351
rect 20729 32317 20763 32351
rect 20763 32317 20772 32351
rect 20720 32308 20772 32317
rect 28908 32308 28960 32360
rect 20076 32283 20128 32292
rect 1492 32215 1544 32224
rect 1492 32181 1501 32215
rect 1501 32181 1535 32215
rect 1535 32181 1544 32215
rect 1492 32172 1544 32181
rect 17960 32172 18012 32224
rect 18696 32172 18748 32224
rect 20076 32249 20085 32283
rect 20085 32249 20119 32283
rect 20119 32249 20128 32283
rect 20076 32240 20128 32249
rect 23388 32240 23440 32292
rect 28448 32240 28500 32292
rect 30380 32308 30432 32360
rect 30472 32240 30524 32292
rect 31208 32376 31260 32428
rect 31668 32376 31720 32428
rect 31944 32308 31996 32360
rect 32220 32376 32272 32428
rect 32680 32376 32732 32428
rect 32864 32419 32916 32428
rect 32864 32385 32873 32419
rect 32873 32385 32907 32419
rect 32907 32385 32916 32419
rect 32864 32376 32916 32385
rect 32956 32376 33008 32428
rect 36176 32444 36228 32496
rect 35716 32376 35768 32428
rect 36084 32376 36136 32428
rect 36268 32419 36320 32428
rect 36268 32385 36277 32419
rect 36277 32385 36311 32419
rect 36311 32385 36320 32419
rect 36268 32376 36320 32385
rect 36636 32376 36688 32428
rect 53564 32419 53616 32428
rect 53564 32385 53573 32419
rect 53573 32385 53607 32419
rect 53607 32385 53616 32419
rect 53564 32376 53616 32385
rect 32496 32240 32548 32292
rect 33048 32240 33100 32292
rect 22652 32215 22704 32224
rect 22652 32181 22661 32215
rect 22661 32181 22695 32215
rect 22695 32181 22704 32215
rect 22652 32172 22704 32181
rect 23296 32215 23348 32224
rect 23296 32181 23305 32215
rect 23305 32181 23339 32215
rect 23339 32181 23348 32215
rect 23296 32172 23348 32181
rect 23756 32215 23808 32224
rect 23756 32181 23765 32215
rect 23765 32181 23799 32215
rect 23799 32181 23808 32215
rect 23756 32172 23808 32181
rect 23848 32172 23900 32224
rect 24676 32215 24728 32224
rect 24676 32181 24685 32215
rect 24685 32181 24719 32215
rect 24719 32181 24728 32215
rect 24676 32172 24728 32181
rect 25596 32172 25648 32224
rect 27712 32172 27764 32224
rect 29736 32172 29788 32224
rect 30932 32172 30984 32224
rect 31392 32215 31444 32224
rect 31392 32181 31401 32215
rect 31401 32181 31435 32215
rect 31435 32181 31444 32215
rect 31392 32172 31444 32181
rect 31484 32215 31536 32224
rect 31484 32181 31493 32215
rect 31493 32181 31527 32215
rect 31527 32181 31536 32215
rect 31484 32172 31536 32181
rect 31668 32172 31720 32224
rect 36728 32308 36780 32360
rect 37648 32351 37700 32360
rect 37648 32317 37657 32351
rect 37657 32317 37691 32351
rect 37691 32317 37700 32351
rect 37648 32308 37700 32317
rect 53380 32283 53432 32292
rect 53380 32249 53389 32283
rect 53389 32249 53423 32283
rect 53423 32249 53432 32283
rect 53380 32240 53432 32249
rect 34336 32172 34388 32224
rect 34704 32215 34756 32224
rect 34704 32181 34713 32215
rect 34713 32181 34747 32215
rect 34747 32181 34756 32215
rect 34704 32172 34756 32181
rect 36360 32215 36412 32224
rect 36360 32181 36369 32215
rect 36369 32181 36403 32215
rect 36403 32181 36412 32215
rect 36360 32172 36412 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 15384 31968 15436 32020
rect 18144 32011 18196 32020
rect 18144 31977 18153 32011
rect 18153 31977 18187 32011
rect 18187 31977 18196 32011
rect 18144 31968 18196 31977
rect 18512 32011 18564 32020
rect 18512 31977 18521 32011
rect 18521 31977 18555 32011
rect 18555 31977 18564 32011
rect 18512 31968 18564 31977
rect 26148 31968 26200 32020
rect 31392 31968 31444 32020
rect 31668 32011 31720 32020
rect 31668 31977 31677 32011
rect 31677 31977 31711 32011
rect 31711 31977 31720 32011
rect 31668 31968 31720 31977
rect 16396 31900 16448 31952
rect 2228 31832 2280 31884
rect 16028 31832 16080 31884
rect 18420 31900 18472 31952
rect 27252 31900 27304 31952
rect 29000 31943 29052 31952
rect 29000 31909 29009 31943
rect 29009 31909 29043 31943
rect 29043 31909 29052 31943
rect 29000 31900 29052 31909
rect 29920 31900 29972 31952
rect 34060 31968 34112 32020
rect 16396 31764 16448 31816
rect 21364 31832 21416 31884
rect 16856 31764 16908 31816
rect 18052 31807 18104 31816
rect 18052 31773 18061 31807
rect 18061 31773 18095 31807
rect 18095 31773 18104 31807
rect 18052 31764 18104 31773
rect 19340 31764 19392 31816
rect 20260 31764 20312 31816
rect 20720 31807 20772 31816
rect 20720 31773 20729 31807
rect 20729 31773 20763 31807
rect 20763 31773 20772 31807
rect 20720 31764 20772 31773
rect 20996 31764 21048 31816
rect 22192 31807 22244 31816
rect 22192 31773 22201 31807
rect 22201 31773 22235 31807
rect 22235 31773 22244 31807
rect 22192 31764 22244 31773
rect 24032 31832 24084 31884
rect 22652 31764 22704 31816
rect 17960 31696 18012 31748
rect 16948 31628 17000 31680
rect 17224 31671 17276 31680
rect 17224 31637 17233 31671
rect 17233 31637 17267 31671
rect 17267 31637 17276 31671
rect 17224 31628 17276 31637
rect 17592 31628 17644 31680
rect 20536 31696 20588 31748
rect 20812 31696 20864 31748
rect 21272 31739 21324 31748
rect 21272 31705 21281 31739
rect 21281 31705 21315 31739
rect 21315 31705 21324 31739
rect 21272 31696 21324 31705
rect 23112 31696 23164 31748
rect 23572 31764 23624 31816
rect 20444 31628 20496 31680
rect 22560 31628 22612 31680
rect 23204 31628 23256 31680
rect 25872 31807 25924 31816
rect 25872 31773 25881 31807
rect 25881 31773 25915 31807
rect 25915 31773 25924 31807
rect 25872 31764 25924 31773
rect 26148 31764 26200 31816
rect 32680 31832 32732 31884
rect 33140 31900 33192 31952
rect 34336 31900 34388 31952
rect 36268 31900 36320 31952
rect 37096 31900 37148 31952
rect 37464 31900 37516 31952
rect 33784 31832 33836 31884
rect 36636 31875 36688 31884
rect 25596 31739 25648 31748
rect 25596 31705 25605 31739
rect 25605 31705 25639 31739
rect 25639 31705 25648 31739
rect 25596 31696 25648 31705
rect 25504 31628 25556 31680
rect 27712 31696 27764 31748
rect 28908 31696 28960 31748
rect 29552 31628 29604 31680
rect 30840 31764 30892 31816
rect 30932 31764 30984 31816
rect 31484 31807 31536 31816
rect 31484 31773 31493 31807
rect 31493 31773 31527 31807
rect 31527 31773 31536 31807
rect 31484 31764 31536 31773
rect 31760 31807 31812 31816
rect 31760 31773 31769 31807
rect 31769 31773 31803 31807
rect 31803 31773 31812 31807
rect 31760 31764 31812 31773
rect 32312 31764 32364 31816
rect 33048 31807 33100 31816
rect 33048 31773 33057 31807
rect 33057 31773 33091 31807
rect 33091 31773 33100 31807
rect 33048 31764 33100 31773
rect 32956 31696 33008 31748
rect 33876 31807 33928 31816
rect 33876 31773 33885 31807
rect 33885 31773 33919 31807
rect 33919 31773 33928 31807
rect 33876 31764 33928 31773
rect 36636 31841 36645 31875
rect 36645 31841 36679 31875
rect 36679 31841 36688 31875
rect 36636 31832 36688 31841
rect 37648 31832 37700 31884
rect 34704 31764 34756 31816
rect 34060 31739 34112 31748
rect 34060 31705 34069 31739
rect 34069 31705 34103 31739
rect 34103 31705 34112 31739
rect 34060 31696 34112 31705
rect 35992 31696 36044 31748
rect 36728 31764 36780 31816
rect 37372 31764 37424 31816
rect 51724 31764 51776 31816
rect 31024 31628 31076 31680
rect 31392 31628 31444 31680
rect 32680 31628 32732 31680
rect 33416 31628 33468 31680
rect 37280 31671 37332 31680
rect 37280 31637 37289 31671
rect 37289 31637 37323 31671
rect 37323 31637 37332 31671
rect 37280 31628 37332 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 16028 31467 16080 31476
rect 16028 31433 16037 31467
rect 16037 31433 16071 31467
rect 16071 31433 16080 31467
rect 16028 31424 16080 31433
rect 18052 31424 18104 31476
rect 18420 31424 18472 31476
rect 16948 31331 17000 31340
rect 16948 31297 16957 31331
rect 16957 31297 16991 31331
rect 16991 31297 17000 31331
rect 16948 31288 17000 31297
rect 17224 31288 17276 31340
rect 17592 31331 17644 31340
rect 17592 31297 17601 31331
rect 17601 31297 17635 31331
rect 17635 31297 17644 31331
rect 17592 31288 17644 31297
rect 17960 31288 18012 31340
rect 18512 31331 18564 31340
rect 18512 31297 18521 31331
rect 18521 31297 18555 31331
rect 18555 31297 18564 31331
rect 18512 31288 18564 31297
rect 18696 31288 18748 31340
rect 19524 31331 19576 31340
rect 19524 31297 19533 31331
rect 19533 31297 19567 31331
rect 19567 31297 19576 31331
rect 19524 31288 19576 31297
rect 19616 31263 19668 31272
rect 19616 31229 19625 31263
rect 19625 31229 19659 31263
rect 19659 31229 19668 31263
rect 19616 31220 19668 31229
rect 20720 31288 20772 31340
rect 23480 31424 23532 31476
rect 23756 31424 23808 31476
rect 25872 31424 25924 31476
rect 22652 31399 22704 31408
rect 22652 31365 22661 31399
rect 22661 31365 22695 31399
rect 22695 31365 22704 31399
rect 22652 31356 22704 31365
rect 24676 31356 24728 31408
rect 22560 31331 22612 31340
rect 20444 31263 20496 31272
rect 20444 31229 20453 31263
rect 20453 31229 20487 31263
rect 20487 31229 20496 31263
rect 20444 31220 20496 31229
rect 22560 31297 22569 31331
rect 22569 31297 22603 31331
rect 22603 31297 22612 31331
rect 22560 31288 22612 31297
rect 23204 31288 23256 31340
rect 23756 31331 23808 31340
rect 23756 31297 23765 31331
rect 23765 31297 23799 31331
rect 23799 31297 23808 31331
rect 23756 31288 23808 31297
rect 22192 31220 22244 31272
rect 23388 31263 23440 31272
rect 23388 31229 23397 31263
rect 23397 31229 23431 31263
rect 23431 31229 23440 31263
rect 25504 31288 25556 31340
rect 25688 31331 25740 31340
rect 25688 31297 25697 31331
rect 25697 31297 25731 31331
rect 25731 31297 25740 31331
rect 25688 31288 25740 31297
rect 25780 31331 25832 31340
rect 25780 31297 25789 31331
rect 25789 31297 25823 31331
rect 25823 31297 25832 31331
rect 26976 31331 27028 31340
rect 25780 31288 25832 31297
rect 26976 31297 26985 31331
rect 26985 31297 27019 31331
rect 27019 31297 27028 31331
rect 26976 31288 27028 31297
rect 27252 31331 27304 31340
rect 27252 31297 27261 31331
rect 27261 31297 27295 31331
rect 27295 31297 27304 31331
rect 27252 31288 27304 31297
rect 28908 31288 28960 31340
rect 29552 31331 29604 31340
rect 29552 31297 29561 31331
rect 29561 31297 29595 31331
rect 29595 31297 29604 31331
rect 29552 31288 29604 31297
rect 32956 31424 33008 31476
rect 33876 31424 33928 31476
rect 37648 31467 37700 31476
rect 37648 31433 37657 31467
rect 37657 31433 37691 31467
rect 37691 31433 37700 31467
rect 37648 31424 37700 31433
rect 32220 31331 32272 31340
rect 32220 31297 32229 31331
rect 32229 31297 32263 31331
rect 32263 31297 32272 31331
rect 32496 31331 32548 31340
rect 32220 31288 32272 31297
rect 32496 31297 32505 31331
rect 32505 31297 32539 31331
rect 32539 31297 32548 31331
rect 32496 31288 32548 31297
rect 33140 31331 33192 31340
rect 33140 31297 33149 31331
rect 33149 31297 33183 31331
rect 33183 31297 33192 31331
rect 33140 31288 33192 31297
rect 34060 31331 34112 31340
rect 34060 31297 34069 31331
rect 34069 31297 34103 31331
rect 34103 31297 34112 31331
rect 34060 31288 34112 31297
rect 35716 31356 35768 31408
rect 23388 31220 23440 31229
rect 31852 31220 31904 31272
rect 27988 31152 28040 31204
rect 16948 31127 17000 31136
rect 16948 31093 16957 31127
rect 16957 31093 16991 31127
rect 16991 31093 17000 31127
rect 16948 31084 17000 31093
rect 18880 31127 18932 31136
rect 18880 31093 18889 31127
rect 18889 31093 18923 31127
rect 18923 31093 18932 31127
rect 18880 31084 18932 31093
rect 22008 31127 22060 31136
rect 22008 31093 22017 31127
rect 22017 31093 22051 31127
rect 22051 31093 22060 31127
rect 22008 31084 22060 31093
rect 24216 31084 24268 31136
rect 24584 31127 24636 31136
rect 24584 31093 24593 31127
rect 24593 31093 24627 31127
rect 24627 31093 24636 31127
rect 24584 31084 24636 31093
rect 28356 31127 28408 31136
rect 28356 31093 28365 31127
rect 28365 31093 28399 31127
rect 28399 31093 28408 31127
rect 28356 31084 28408 31093
rect 29828 31084 29880 31136
rect 30380 31152 30432 31204
rect 30840 31152 30892 31204
rect 31760 31152 31812 31204
rect 31944 31152 31996 31204
rect 32772 31220 32824 31272
rect 33416 31220 33468 31272
rect 33784 31220 33836 31272
rect 35440 31288 35492 31340
rect 36268 31331 36320 31340
rect 36268 31297 36277 31331
rect 36277 31297 36311 31331
rect 36311 31297 36320 31331
rect 36268 31288 36320 31297
rect 34704 31220 34756 31272
rect 37280 31356 37332 31408
rect 36544 31288 36596 31340
rect 36452 31152 36504 31204
rect 32496 31127 32548 31136
rect 32496 31093 32505 31127
rect 32505 31093 32539 31127
rect 32539 31093 32548 31127
rect 32496 31084 32548 31093
rect 32956 31127 33008 31136
rect 32956 31093 32965 31127
rect 32965 31093 32999 31127
rect 32999 31093 33008 31127
rect 32956 31084 33008 31093
rect 36636 31084 36688 31136
rect 38200 31127 38252 31136
rect 38200 31093 38209 31127
rect 38209 31093 38243 31127
rect 38243 31093 38252 31127
rect 38200 31084 38252 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 22192 30880 22244 30932
rect 23664 30880 23716 30932
rect 25688 30880 25740 30932
rect 26056 30923 26108 30932
rect 26056 30889 26065 30923
rect 26065 30889 26099 30923
rect 26099 30889 26108 30923
rect 26056 30880 26108 30889
rect 19616 30812 19668 30864
rect 18328 30787 18380 30796
rect 18328 30753 18337 30787
rect 18337 30753 18371 30787
rect 18371 30753 18380 30787
rect 18328 30744 18380 30753
rect 16948 30676 17000 30728
rect 25320 30812 25372 30864
rect 22008 30744 22060 30796
rect 24952 30744 25004 30796
rect 27344 30880 27396 30932
rect 31208 30880 31260 30932
rect 31944 30923 31996 30932
rect 31944 30889 31953 30923
rect 31953 30889 31987 30923
rect 31987 30889 31996 30923
rect 31944 30880 31996 30889
rect 32220 30880 32272 30932
rect 32772 30923 32824 30932
rect 32772 30889 32781 30923
rect 32781 30889 32815 30923
rect 32815 30889 32824 30923
rect 32772 30880 32824 30889
rect 34704 30923 34756 30932
rect 34704 30889 34713 30923
rect 34713 30889 34747 30923
rect 34747 30889 34756 30923
rect 34704 30880 34756 30889
rect 36084 30880 36136 30932
rect 36544 30880 36596 30932
rect 32128 30744 32180 30796
rect 33784 30787 33836 30796
rect 33784 30753 33793 30787
rect 33793 30753 33827 30787
rect 33827 30753 33836 30787
rect 33784 30744 33836 30753
rect 36360 30787 36412 30796
rect 36360 30753 36369 30787
rect 36369 30753 36403 30787
rect 36403 30753 36412 30787
rect 36360 30744 36412 30753
rect 37372 30812 37424 30864
rect 36636 30787 36688 30796
rect 36636 30753 36645 30787
rect 36645 30753 36679 30787
rect 36679 30753 36688 30787
rect 36636 30744 36688 30753
rect 20260 30676 20312 30728
rect 19524 30608 19576 30660
rect 21364 30676 21416 30728
rect 23204 30719 23256 30728
rect 21272 30608 21324 30660
rect 23204 30685 23213 30719
rect 23213 30685 23247 30719
rect 23247 30685 23256 30719
rect 23204 30676 23256 30685
rect 23572 30676 23624 30728
rect 24584 30676 24636 30728
rect 24768 30719 24820 30728
rect 24768 30685 24777 30719
rect 24777 30685 24811 30719
rect 24811 30685 24820 30719
rect 24768 30676 24820 30685
rect 26148 30719 26200 30728
rect 26148 30685 26157 30719
rect 26157 30685 26191 30719
rect 26191 30685 26200 30719
rect 26148 30676 26200 30685
rect 28356 30676 28408 30728
rect 29828 30719 29880 30728
rect 29828 30685 29837 30719
rect 29837 30685 29871 30719
rect 29871 30685 29880 30719
rect 29828 30676 29880 30685
rect 31852 30676 31904 30728
rect 2136 30540 2188 30592
rect 17592 30540 17644 30592
rect 20812 30583 20864 30592
rect 20812 30549 20821 30583
rect 20821 30549 20855 30583
rect 20855 30549 20864 30583
rect 20812 30540 20864 30549
rect 23756 30608 23808 30660
rect 32956 30676 33008 30728
rect 34060 30676 34112 30728
rect 35440 30676 35492 30728
rect 35716 30719 35768 30728
rect 32864 30608 32916 30660
rect 35716 30685 35725 30719
rect 35725 30685 35759 30719
rect 35759 30685 35768 30719
rect 35716 30676 35768 30685
rect 37464 30676 37516 30728
rect 24400 30583 24452 30592
rect 24400 30549 24409 30583
rect 24409 30549 24443 30583
rect 24443 30549 24452 30583
rect 24400 30540 24452 30549
rect 27712 30583 27764 30592
rect 27712 30549 27721 30583
rect 27721 30549 27755 30583
rect 27755 30549 27764 30583
rect 27712 30540 27764 30549
rect 36176 30583 36228 30592
rect 36176 30549 36185 30583
rect 36185 30549 36219 30583
rect 36219 30549 36228 30583
rect 36176 30540 36228 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 23388 30336 23440 30388
rect 24768 30336 24820 30388
rect 25780 30336 25832 30388
rect 30656 30336 30708 30388
rect 31024 30379 31076 30388
rect 31024 30345 31033 30379
rect 31033 30345 31067 30379
rect 31067 30345 31076 30379
rect 31024 30336 31076 30345
rect 34060 30379 34112 30388
rect 34060 30345 34069 30379
rect 34069 30345 34103 30379
rect 34103 30345 34112 30379
rect 34060 30336 34112 30345
rect 36268 30379 36320 30388
rect 36268 30345 36277 30379
rect 36277 30345 36311 30379
rect 36311 30345 36320 30379
rect 36268 30336 36320 30345
rect 38200 30336 38252 30388
rect 19432 30268 19484 30320
rect 20904 30268 20956 30320
rect 21456 30268 21508 30320
rect 23480 30268 23532 30320
rect 26056 30268 26108 30320
rect 32496 30268 32548 30320
rect 20720 30200 20772 30252
rect 20996 30243 21048 30252
rect 20996 30209 21005 30243
rect 21005 30209 21039 30243
rect 21039 30209 21048 30243
rect 20996 30200 21048 30209
rect 21824 30243 21876 30252
rect 21824 30209 21833 30243
rect 21833 30209 21867 30243
rect 21867 30209 21876 30243
rect 21824 30200 21876 30209
rect 22100 30200 22152 30252
rect 20260 30132 20312 30184
rect 23388 30200 23440 30252
rect 23572 30243 23624 30252
rect 23572 30209 23581 30243
rect 23581 30209 23615 30243
rect 23615 30209 23624 30243
rect 23572 30200 23624 30209
rect 23756 30243 23808 30252
rect 23756 30209 23765 30243
rect 23765 30209 23799 30243
rect 23799 30209 23808 30243
rect 23756 30200 23808 30209
rect 24400 30243 24452 30252
rect 23664 30132 23716 30184
rect 23940 30132 23992 30184
rect 24400 30209 24409 30243
rect 24409 30209 24443 30243
rect 24443 30209 24452 30243
rect 24400 30200 24452 30209
rect 24860 30243 24912 30252
rect 24860 30209 24869 30243
rect 24869 30209 24903 30243
rect 24903 30209 24912 30243
rect 24860 30200 24912 30209
rect 25596 30200 25648 30252
rect 26240 30200 26292 30252
rect 26976 30243 27028 30252
rect 26976 30209 26985 30243
rect 26985 30209 27019 30243
rect 27019 30209 27028 30243
rect 26976 30200 27028 30209
rect 47584 30268 47636 30320
rect 35164 30243 35216 30252
rect 25320 30132 25372 30184
rect 26148 30132 26200 30184
rect 17960 30039 18012 30048
rect 17960 30005 17969 30039
rect 17969 30005 18003 30039
rect 18003 30005 18012 30039
rect 17960 29996 18012 30005
rect 20352 30039 20404 30048
rect 20352 30005 20361 30039
rect 20361 30005 20395 30039
rect 20395 30005 20404 30039
rect 20352 29996 20404 30005
rect 22008 29996 22060 30048
rect 26056 29996 26108 30048
rect 32128 30175 32180 30184
rect 32128 30141 32137 30175
rect 32137 30141 32171 30175
rect 32171 30141 32180 30175
rect 32128 30132 32180 30141
rect 35164 30209 35173 30243
rect 35173 30209 35207 30243
rect 35207 30209 35216 30243
rect 35164 30200 35216 30209
rect 35716 30200 35768 30252
rect 36084 30200 36136 30252
rect 36452 30200 36504 30252
rect 53564 30243 53616 30252
rect 53564 30209 53573 30243
rect 53573 30209 53607 30243
rect 53607 30209 53616 30243
rect 53564 30200 53616 30209
rect 35808 30132 35860 30184
rect 32496 29996 32548 30048
rect 35992 29996 36044 30048
rect 36452 29996 36504 30048
rect 53472 30039 53524 30048
rect 53472 30005 53481 30039
rect 53481 30005 53515 30039
rect 53515 30005 53524 30039
rect 53472 29996 53524 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 22928 29792 22980 29844
rect 23204 29792 23256 29844
rect 23756 29792 23808 29844
rect 24860 29792 24912 29844
rect 26148 29835 26200 29844
rect 26148 29801 26157 29835
rect 26157 29801 26191 29835
rect 26191 29801 26200 29835
rect 26148 29792 26200 29801
rect 31208 29792 31260 29844
rect 33048 29835 33100 29844
rect 33048 29801 33057 29835
rect 33057 29801 33091 29835
rect 33091 29801 33100 29835
rect 33048 29792 33100 29801
rect 33324 29792 33376 29844
rect 34152 29792 34204 29844
rect 36452 29835 36504 29844
rect 36452 29801 36461 29835
rect 36461 29801 36495 29835
rect 36495 29801 36504 29835
rect 36452 29792 36504 29801
rect 20352 29724 20404 29776
rect 20904 29724 20956 29776
rect 20812 29656 20864 29708
rect 21272 29656 21324 29708
rect 1400 29631 1452 29640
rect 1400 29597 1409 29631
rect 1409 29597 1443 29631
rect 1443 29597 1452 29631
rect 1400 29588 1452 29597
rect 19248 29588 19300 29640
rect 19984 29588 20036 29640
rect 21456 29588 21508 29640
rect 23296 29724 23348 29776
rect 23388 29656 23440 29708
rect 22008 29588 22060 29640
rect 20168 29520 20220 29572
rect 18144 29495 18196 29504
rect 18144 29461 18153 29495
rect 18153 29461 18187 29495
rect 18187 29461 18196 29495
rect 18144 29452 18196 29461
rect 19340 29452 19392 29504
rect 22284 29520 22336 29572
rect 23112 29588 23164 29640
rect 24952 29656 25004 29708
rect 25504 29656 25556 29708
rect 23204 29520 23256 29572
rect 23848 29588 23900 29640
rect 31668 29724 31720 29776
rect 26976 29656 27028 29708
rect 27804 29656 27856 29708
rect 31484 29656 31536 29708
rect 32772 29724 32824 29776
rect 53472 29724 53524 29776
rect 33324 29656 33376 29708
rect 33784 29656 33836 29708
rect 23756 29520 23808 29572
rect 22836 29495 22888 29504
rect 22836 29461 22845 29495
rect 22845 29461 22879 29495
rect 22879 29461 22888 29495
rect 22836 29452 22888 29461
rect 25780 29588 25832 29640
rect 27252 29588 27304 29640
rect 28816 29631 28868 29640
rect 28816 29597 28825 29631
rect 28825 29597 28859 29631
rect 28859 29597 28868 29631
rect 28816 29588 28868 29597
rect 29828 29588 29880 29640
rect 31668 29633 31720 29640
rect 31668 29599 31677 29633
rect 31677 29599 31711 29633
rect 31711 29599 31720 29633
rect 31852 29631 31904 29640
rect 31668 29588 31720 29599
rect 31852 29597 31861 29631
rect 31861 29597 31895 29631
rect 31895 29597 31904 29631
rect 31852 29588 31904 29597
rect 25412 29452 25464 29504
rect 26056 29452 26108 29504
rect 27620 29452 27672 29504
rect 29092 29452 29144 29504
rect 30380 29452 30432 29504
rect 31392 29452 31444 29504
rect 32588 29588 32640 29640
rect 33140 29588 33192 29640
rect 36176 29656 36228 29708
rect 35716 29631 35768 29640
rect 35716 29597 35725 29631
rect 35725 29597 35759 29631
rect 35759 29597 35768 29631
rect 35716 29588 35768 29597
rect 36636 29588 36688 29640
rect 33416 29520 33468 29572
rect 32404 29495 32456 29504
rect 32404 29461 32413 29495
rect 32413 29461 32447 29495
rect 32447 29461 32456 29495
rect 32404 29452 32456 29461
rect 33324 29452 33376 29504
rect 36268 29495 36320 29504
rect 36268 29461 36277 29495
rect 36277 29461 36311 29495
rect 36311 29461 36320 29495
rect 36268 29452 36320 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 1400 29291 1452 29300
rect 1400 29257 1409 29291
rect 1409 29257 1443 29291
rect 1443 29257 1452 29291
rect 1400 29248 1452 29257
rect 19248 29291 19300 29300
rect 19248 29257 19257 29291
rect 19257 29257 19291 29291
rect 19291 29257 19300 29291
rect 19248 29248 19300 29257
rect 20812 29248 20864 29300
rect 22100 29248 22152 29300
rect 23480 29248 23532 29300
rect 23848 29291 23900 29300
rect 23848 29257 23857 29291
rect 23857 29257 23891 29291
rect 23891 29257 23900 29291
rect 23848 29248 23900 29257
rect 18144 29223 18196 29232
rect 18144 29189 18153 29223
rect 18153 29189 18187 29223
rect 18187 29189 18196 29223
rect 20168 29223 20220 29232
rect 18144 29180 18196 29189
rect 20168 29189 20177 29223
rect 20177 29189 20211 29223
rect 20211 29189 20220 29223
rect 33600 29248 33652 29300
rect 20168 29180 20220 29189
rect 20260 29112 20312 29164
rect 20904 29155 20956 29164
rect 20904 29121 20913 29155
rect 20913 29121 20947 29155
rect 20947 29121 20956 29155
rect 20904 29112 20956 29121
rect 21732 29112 21784 29164
rect 22100 29155 22152 29164
rect 22100 29121 22109 29155
rect 22109 29121 22143 29155
rect 22143 29121 22152 29155
rect 22100 29112 22152 29121
rect 22836 29112 22888 29164
rect 23112 29155 23164 29164
rect 23112 29121 23121 29155
rect 23121 29121 23155 29155
rect 23155 29121 23164 29155
rect 25412 29180 25464 29232
rect 23112 29112 23164 29121
rect 25780 29112 25832 29164
rect 26240 29180 26292 29232
rect 26056 29155 26108 29164
rect 26056 29121 26065 29155
rect 26065 29121 26099 29155
rect 26099 29121 26108 29155
rect 26056 29112 26108 29121
rect 23296 29087 23348 29096
rect 23296 29053 23305 29087
rect 23305 29053 23339 29087
rect 23339 29053 23348 29087
rect 23296 29044 23348 29053
rect 26148 29087 26200 29096
rect 26148 29053 26157 29087
rect 26157 29053 26191 29087
rect 26191 29053 26200 29087
rect 26148 29044 26200 29053
rect 26332 29044 26384 29096
rect 20352 28976 20404 29028
rect 20720 28976 20772 29028
rect 22008 28976 22060 29028
rect 24860 28976 24912 29028
rect 27804 29112 27856 29164
rect 28540 29112 28592 29164
rect 31576 29180 31628 29232
rect 33876 29248 33928 29300
rect 53380 29248 53432 29300
rect 31300 29112 31352 29164
rect 32036 29112 32088 29164
rect 32588 29112 32640 29164
rect 19800 28951 19852 28960
rect 19800 28917 19809 28951
rect 19809 28917 19843 28951
rect 19843 28917 19852 28951
rect 19800 28908 19852 28917
rect 20904 28951 20956 28960
rect 20904 28917 20913 28951
rect 20913 28917 20947 28951
rect 20947 28917 20956 28951
rect 20904 28908 20956 28917
rect 22376 28908 22428 28960
rect 22560 28951 22612 28960
rect 22560 28917 22569 28951
rect 22569 28917 22603 28951
rect 22603 28917 22612 28951
rect 22560 28908 22612 28917
rect 24952 28951 25004 28960
rect 24952 28917 24961 28951
rect 24961 28917 24995 28951
rect 24995 28917 25004 28951
rect 24952 28908 25004 28917
rect 25136 28951 25188 28960
rect 25136 28917 25145 28951
rect 25145 28917 25179 28951
rect 25179 28917 25188 28951
rect 25136 28908 25188 28917
rect 25504 28908 25556 28960
rect 27436 28976 27488 29028
rect 27712 28976 27764 29028
rect 26976 28951 27028 28960
rect 26976 28917 26985 28951
rect 26985 28917 27019 28951
rect 27019 28917 27028 28951
rect 26976 28908 27028 28917
rect 28724 28908 28776 28960
rect 29644 28976 29696 29028
rect 29828 29019 29880 29028
rect 29828 28985 29837 29019
rect 29837 28985 29871 29019
rect 29871 28985 29880 29019
rect 29828 28976 29880 28985
rect 31300 28976 31352 29028
rect 34428 29044 34480 29096
rect 36176 29112 36228 29164
rect 35348 29044 35400 29096
rect 35624 29044 35676 29096
rect 36452 29087 36504 29096
rect 36452 29053 36461 29087
rect 36461 29053 36495 29087
rect 36495 29053 36504 29087
rect 36452 29044 36504 29053
rect 35808 28976 35860 29028
rect 30656 28908 30708 28960
rect 31944 28908 31996 28960
rect 33968 28908 34020 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 18880 28704 18932 28756
rect 19432 28704 19484 28756
rect 21272 28747 21324 28756
rect 18788 28636 18840 28688
rect 19984 28636 20036 28688
rect 21272 28713 21281 28747
rect 21281 28713 21315 28747
rect 21315 28713 21324 28747
rect 21272 28704 21324 28713
rect 23664 28636 23716 28688
rect 19340 28568 19392 28620
rect 17224 28500 17276 28552
rect 20076 28568 20128 28620
rect 19616 28543 19668 28552
rect 19616 28509 19625 28543
rect 19625 28509 19659 28543
rect 19659 28509 19668 28543
rect 19616 28500 19668 28509
rect 19800 28543 19852 28552
rect 19800 28509 19809 28543
rect 19809 28509 19843 28543
rect 19843 28509 19852 28543
rect 19800 28500 19852 28509
rect 20904 28500 20956 28552
rect 21272 28543 21324 28552
rect 21272 28509 21281 28543
rect 21281 28509 21315 28543
rect 21315 28509 21324 28543
rect 21272 28500 21324 28509
rect 22100 28543 22152 28552
rect 22100 28509 22109 28543
rect 22109 28509 22143 28543
rect 22143 28509 22152 28543
rect 22100 28500 22152 28509
rect 22284 28543 22336 28552
rect 22284 28509 22293 28543
rect 22293 28509 22327 28543
rect 22327 28509 22336 28543
rect 22284 28500 22336 28509
rect 19340 28407 19392 28416
rect 19340 28373 19349 28407
rect 19349 28373 19383 28407
rect 19383 28373 19392 28407
rect 19340 28364 19392 28373
rect 22008 28432 22060 28484
rect 23112 28432 23164 28484
rect 23388 28475 23440 28484
rect 23388 28441 23397 28475
rect 23397 28441 23431 28475
rect 23431 28441 23440 28475
rect 23388 28432 23440 28441
rect 20812 28364 20864 28416
rect 22652 28364 22704 28416
rect 23940 28364 23992 28416
rect 24124 28364 24176 28416
rect 25136 28636 25188 28688
rect 25320 28636 25372 28688
rect 28540 28704 28592 28756
rect 27804 28611 27856 28620
rect 27804 28577 27813 28611
rect 27813 28577 27847 28611
rect 27847 28577 27856 28611
rect 27804 28568 27856 28577
rect 25136 28543 25188 28552
rect 25136 28509 25145 28543
rect 25145 28509 25179 28543
rect 25179 28509 25188 28543
rect 25136 28500 25188 28509
rect 25320 28543 25372 28552
rect 25320 28509 25329 28543
rect 25329 28509 25363 28543
rect 25363 28509 25372 28543
rect 25320 28500 25372 28509
rect 26976 28500 27028 28552
rect 28448 28543 28500 28552
rect 28448 28509 28457 28543
rect 28457 28509 28491 28543
rect 28491 28509 28500 28543
rect 28448 28500 28500 28509
rect 29000 28500 29052 28552
rect 29828 28543 29880 28552
rect 29828 28509 29837 28543
rect 29837 28509 29871 28543
rect 29871 28509 29880 28543
rect 29828 28500 29880 28509
rect 32312 28704 32364 28756
rect 32588 28704 32640 28756
rect 35808 28747 35860 28756
rect 35808 28713 35817 28747
rect 35817 28713 35851 28747
rect 35851 28713 35860 28747
rect 35808 28704 35860 28713
rect 35532 28636 35584 28688
rect 37832 28636 37884 28688
rect 32496 28611 32548 28620
rect 32496 28577 32505 28611
rect 32505 28577 32539 28611
rect 32539 28577 32548 28611
rect 32496 28568 32548 28577
rect 33416 28568 33468 28620
rect 25412 28432 25464 28484
rect 27804 28432 27856 28484
rect 30380 28432 30432 28484
rect 32404 28500 32456 28552
rect 32956 28543 33008 28552
rect 32956 28509 32965 28543
rect 32965 28509 32999 28543
rect 32999 28509 33008 28543
rect 32956 28500 33008 28509
rect 33968 28543 34020 28552
rect 33968 28509 33977 28543
rect 33977 28509 34011 28543
rect 34011 28509 34020 28543
rect 33968 28500 34020 28509
rect 34980 28543 35032 28552
rect 26332 28364 26384 28416
rect 28080 28364 28132 28416
rect 30840 28364 30892 28416
rect 31392 28364 31444 28416
rect 31576 28364 31628 28416
rect 34980 28509 34988 28543
rect 34988 28509 35022 28543
rect 35022 28509 35032 28543
rect 34980 28500 35032 28509
rect 36268 28568 36320 28620
rect 35348 28543 35400 28552
rect 35348 28509 35357 28543
rect 35357 28509 35391 28543
rect 35391 28509 35400 28543
rect 35348 28500 35400 28509
rect 35900 28500 35952 28552
rect 35532 28432 35584 28484
rect 35900 28364 35952 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 19984 28160 20036 28212
rect 22008 28160 22060 28212
rect 22376 28160 22428 28212
rect 23388 28160 23440 28212
rect 23940 28203 23992 28212
rect 23940 28169 23949 28203
rect 23949 28169 23983 28203
rect 23983 28169 23992 28203
rect 23940 28160 23992 28169
rect 25320 28203 25372 28212
rect 25320 28169 25329 28203
rect 25329 28169 25363 28203
rect 25363 28169 25372 28203
rect 25320 28160 25372 28169
rect 26332 28203 26384 28212
rect 26332 28169 26341 28203
rect 26341 28169 26375 28203
rect 26375 28169 26384 28203
rect 26332 28160 26384 28169
rect 27804 28203 27856 28212
rect 27804 28169 27813 28203
rect 27813 28169 27847 28203
rect 27847 28169 27856 28203
rect 27804 28160 27856 28169
rect 20352 28092 20404 28144
rect 20720 28135 20772 28144
rect 20720 28101 20745 28135
rect 20745 28101 20772 28135
rect 20720 28092 20772 28101
rect 21916 28092 21968 28144
rect 23664 28092 23716 28144
rect 24124 28135 24176 28144
rect 24124 28101 24133 28135
rect 24133 28101 24167 28135
rect 24167 28101 24176 28135
rect 24124 28092 24176 28101
rect 20168 28024 20220 28076
rect 22008 28067 22060 28076
rect 22008 28033 22017 28067
rect 22017 28033 22051 28067
rect 22051 28033 22060 28067
rect 22008 28024 22060 28033
rect 23112 28067 23164 28076
rect 20260 27956 20312 28008
rect 21456 27956 21508 28008
rect 23112 28033 23121 28067
rect 23121 28033 23155 28067
rect 23155 28033 23164 28067
rect 23112 28024 23164 28033
rect 23388 28067 23440 28076
rect 23388 28033 23397 28067
rect 23397 28033 23431 28067
rect 23431 28033 23440 28067
rect 23388 28024 23440 28033
rect 24584 28067 24636 28076
rect 24584 28033 24593 28067
rect 24593 28033 24627 28067
rect 24627 28033 24636 28067
rect 24584 28024 24636 28033
rect 24952 28024 25004 28076
rect 25596 28092 25648 28144
rect 26148 28092 26200 28144
rect 28724 28135 28776 28144
rect 28724 28101 28733 28135
rect 28733 28101 28767 28135
rect 28767 28101 28776 28135
rect 28724 28092 28776 28101
rect 28816 28092 28868 28144
rect 31852 28160 31904 28212
rect 35348 28160 35400 28212
rect 36452 28160 36504 28212
rect 37832 28203 37884 28212
rect 37832 28169 37841 28203
rect 37841 28169 37875 28203
rect 37875 28169 37884 28203
rect 37832 28160 37884 28169
rect 31300 28135 31352 28144
rect 31300 28101 31309 28135
rect 31309 28101 31343 28135
rect 31343 28101 31352 28135
rect 31300 28092 31352 28101
rect 32128 28092 32180 28144
rect 33968 28092 34020 28144
rect 24768 27956 24820 28008
rect 25872 28024 25924 28076
rect 27436 28024 27488 28076
rect 28080 28067 28132 28076
rect 28080 28033 28089 28067
rect 28089 28033 28123 28067
rect 28123 28033 28132 28067
rect 28080 28024 28132 28033
rect 27896 27956 27948 28008
rect 29828 28024 29880 28076
rect 30840 28024 30892 28076
rect 30932 28067 30984 28076
rect 30932 28033 30941 28067
rect 30941 28033 30975 28067
rect 30975 28033 30984 28067
rect 30932 28024 30984 28033
rect 29092 27956 29144 28008
rect 31576 28024 31628 28076
rect 32312 28067 32364 28076
rect 32312 28033 32321 28067
rect 32321 28033 32355 28067
rect 32355 28033 32364 28067
rect 32312 28024 32364 28033
rect 32680 28024 32732 28076
rect 32036 27956 32088 28008
rect 20812 27820 20864 27872
rect 21272 27820 21324 27872
rect 23204 27820 23256 27872
rect 24952 27888 25004 27940
rect 26056 27888 26108 27940
rect 27252 27931 27304 27940
rect 27252 27897 27261 27931
rect 27261 27897 27295 27931
rect 27295 27897 27304 27931
rect 27252 27888 27304 27897
rect 28448 27888 28500 27940
rect 25320 27820 25372 27872
rect 25504 27863 25556 27872
rect 25504 27829 25513 27863
rect 25513 27829 25547 27863
rect 25547 27829 25556 27863
rect 25504 27820 25556 27829
rect 28724 27820 28776 27872
rect 30380 27888 30432 27940
rect 30932 27888 30984 27940
rect 31024 27888 31076 27940
rect 31668 27888 31720 27940
rect 34428 28024 34480 28076
rect 35624 28092 35676 28144
rect 35532 28067 35584 28076
rect 35532 28033 35541 28067
rect 35541 28033 35575 28067
rect 35575 28033 35584 28067
rect 35532 28024 35584 28033
rect 35900 28024 35952 28076
rect 34244 27999 34296 28008
rect 34244 27965 34253 27999
rect 34253 27965 34287 27999
rect 34287 27965 34296 27999
rect 34244 27956 34296 27965
rect 34060 27888 34112 27940
rect 36452 28024 36504 28076
rect 53380 27999 53432 28008
rect 53380 27965 53389 27999
rect 53389 27965 53423 27999
rect 53423 27965 53432 27999
rect 53380 27956 53432 27965
rect 53656 27999 53708 28008
rect 53656 27965 53665 27999
rect 53665 27965 53699 27999
rect 53699 27965 53708 27999
rect 53656 27956 53708 27965
rect 37556 27888 37608 27940
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 18880 27616 18932 27668
rect 21364 27616 21416 27668
rect 22376 27616 22428 27668
rect 23388 27616 23440 27668
rect 25688 27616 25740 27668
rect 27896 27659 27948 27668
rect 27896 27625 27905 27659
rect 27905 27625 27939 27659
rect 27939 27625 27948 27659
rect 27896 27616 27948 27625
rect 31300 27659 31352 27668
rect 31300 27625 31309 27659
rect 31309 27625 31343 27659
rect 31343 27625 31352 27659
rect 31300 27616 31352 27625
rect 36452 27659 36504 27668
rect 20720 27548 20772 27600
rect 25872 27591 25924 27600
rect 25872 27557 25881 27591
rect 25881 27557 25915 27591
rect 25915 27557 25924 27591
rect 25872 27548 25924 27557
rect 21456 27523 21508 27532
rect 21456 27489 21465 27523
rect 21465 27489 21499 27523
rect 21499 27489 21508 27523
rect 21456 27480 21508 27489
rect 23664 27480 23716 27532
rect 28816 27548 28868 27600
rect 29000 27591 29052 27600
rect 29000 27557 29009 27591
rect 29009 27557 29043 27591
rect 29043 27557 29052 27591
rect 29000 27548 29052 27557
rect 29644 27591 29696 27600
rect 29644 27557 29653 27591
rect 29653 27557 29687 27591
rect 29687 27557 29696 27591
rect 29644 27548 29696 27557
rect 30932 27548 30984 27600
rect 31484 27591 31536 27600
rect 31484 27557 31493 27591
rect 31493 27557 31527 27591
rect 31527 27557 31536 27591
rect 31484 27548 31536 27557
rect 19432 27412 19484 27464
rect 20076 27412 20128 27464
rect 21088 27412 21140 27464
rect 21916 27412 21968 27464
rect 22560 27412 22612 27464
rect 24124 27412 24176 27464
rect 16580 27344 16632 27396
rect 22192 27344 22244 27396
rect 22652 27387 22704 27396
rect 22652 27353 22661 27387
rect 22661 27353 22695 27387
rect 22695 27353 22704 27387
rect 22652 27344 22704 27353
rect 1492 27319 1544 27328
rect 1492 27285 1501 27319
rect 1501 27285 1535 27319
rect 1535 27285 1544 27319
rect 1492 27276 1544 27285
rect 22284 27276 22336 27328
rect 25320 27412 25372 27464
rect 27620 27480 27672 27532
rect 29552 27480 29604 27532
rect 31576 27480 31628 27532
rect 31944 27523 31996 27532
rect 31944 27489 31953 27523
rect 31953 27489 31987 27523
rect 31987 27489 31996 27523
rect 31944 27480 31996 27489
rect 25688 27455 25740 27464
rect 25688 27421 25697 27455
rect 25697 27421 25731 27455
rect 25731 27421 25740 27455
rect 25688 27412 25740 27421
rect 26056 27412 26108 27464
rect 26608 27455 26660 27464
rect 26608 27421 26617 27455
rect 26617 27421 26651 27455
rect 26651 27421 26660 27455
rect 26608 27412 26660 27421
rect 28172 27412 28224 27464
rect 28724 27455 28776 27464
rect 28724 27421 28733 27455
rect 28733 27421 28767 27455
rect 28767 27421 28776 27455
rect 28724 27412 28776 27421
rect 29092 27412 29144 27464
rect 30012 27412 30064 27464
rect 32128 27455 32180 27464
rect 25964 27276 26016 27328
rect 27620 27344 27672 27396
rect 28632 27387 28684 27396
rect 28632 27353 28641 27387
rect 28641 27353 28675 27387
rect 28675 27353 28684 27387
rect 28632 27344 28684 27353
rect 31024 27344 31076 27396
rect 32128 27421 32137 27455
rect 32137 27421 32171 27455
rect 32171 27421 32180 27455
rect 32128 27412 32180 27421
rect 32404 27412 32456 27464
rect 36452 27625 36461 27659
rect 36461 27625 36495 27659
rect 36495 27625 36504 27659
rect 36452 27616 36504 27625
rect 37556 27659 37608 27668
rect 37556 27625 37565 27659
rect 37565 27625 37599 27659
rect 37599 27625 37608 27659
rect 37556 27616 37608 27625
rect 53656 27659 53708 27668
rect 53656 27625 53665 27659
rect 53665 27625 53699 27659
rect 53699 27625 53708 27659
rect 53656 27616 53708 27625
rect 34152 27480 34204 27532
rect 33784 27455 33836 27464
rect 33784 27421 33793 27455
rect 33793 27421 33827 27455
rect 33827 27421 33836 27455
rect 33784 27412 33836 27421
rect 35348 27455 35400 27464
rect 35348 27421 35357 27455
rect 35357 27421 35391 27455
rect 35391 27421 35400 27455
rect 35348 27412 35400 27421
rect 31484 27344 31536 27396
rect 27804 27276 27856 27328
rect 30380 27276 30432 27328
rect 35900 27319 35952 27328
rect 35900 27285 35909 27319
rect 35909 27285 35943 27319
rect 35943 27285 35952 27319
rect 35900 27276 35952 27285
rect 37556 27276 37608 27328
rect 41512 27276 41564 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 20168 27072 20220 27124
rect 24124 27072 24176 27124
rect 25136 27072 25188 27124
rect 25412 27072 25464 27124
rect 26148 27115 26200 27124
rect 26148 27081 26157 27115
rect 26157 27081 26191 27115
rect 26191 27081 26200 27115
rect 26148 27072 26200 27081
rect 28632 27115 28684 27124
rect 20260 27004 20312 27056
rect 23204 27047 23256 27056
rect 23204 27013 23213 27047
rect 23213 27013 23247 27047
rect 23247 27013 23256 27047
rect 23204 27004 23256 27013
rect 25596 27004 25648 27056
rect 28632 27081 28641 27115
rect 28641 27081 28675 27115
rect 28675 27081 28684 27115
rect 28632 27072 28684 27081
rect 29552 27115 29604 27124
rect 29552 27081 29561 27115
rect 29561 27081 29595 27115
rect 29595 27081 29604 27115
rect 29552 27072 29604 27081
rect 30380 27115 30432 27124
rect 30380 27081 30389 27115
rect 30389 27081 30423 27115
rect 30423 27081 30432 27115
rect 30380 27072 30432 27081
rect 30840 27072 30892 27124
rect 27620 27004 27672 27056
rect 20996 26979 21048 26988
rect 20996 26945 21005 26979
rect 21005 26945 21039 26979
rect 21039 26945 21048 26979
rect 20996 26936 21048 26945
rect 21456 26936 21508 26988
rect 22192 26979 22244 26988
rect 22192 26945 22201 26979
rect 22201 26945 22235 26979
rect 22235 26945 22244 26979
rect 22192 26936 22244 26945
rect 22284 26979 22336 26988
rect 22284 26945 22293 26979
rect 22293 26945 22327 26979
rect 22327 26945 22336 26979
rect 22284 26936 22336 26945
rect 22560 26936 22612 26988
rect 24216 26979 24268 26988
rect 24216 26945 24225 26979
rect 24225 26945 24259 26979
rect 24259 26945 24268 26979
rect 24216 26936 24268 26945
rect 24492 26936 24544 26988
rect 26240 26979 26292 26988
rect 26240 26945 26249 26979
rect 26249 26945 26283 26979
rect 26283 26945 26292 26979
rect 26240 26936 26292 26945
rect 21272 26911 21324 26920
rect 21272 26877 21281 26911
rect 21281 26877 21315 26911
rect 21315 26877 21324 26911
rect 21272 26868 21324 26877
rect 22652 26868 22704 26920
rect 25228 26868 25280 26920
rect 26148 26868 26200 26920
rect 27344 26936 27396 26988
rect 27896 26979 27948 26988
rect 27896 26945 27905 26979
rect 27905 26945 27939 26979
rect 27939 26945 27948 26979
rect 27896 26936 27948 26945
rect 27988 26979 28040 26988
rect 27988 26945 27997 26979
rect 27997 26945 28031 26979
rect 28031 26945 28040 26979
rect 27988 26936 28040 26945
rect 28264 26936 28316 26988
rect 30104 26979 30156 26988
rect 30104 26945 30113 26979
rect 30113 26945 30147 26979
rect 30147 26945 30156 26979
rect 30104 26936 30156 26945
rect 29184 26911 29236 26920
rect 26424 26800 26476 26852
rect 29184 26877 29193 26911
rect 29193 26877 29227 26911
rect 29227 26877 29236 26911
rect 29184 26868 29236 26877
rect 29276 26868 29328 26920
rect 30380 26911 30432 26920
rect 30380 26877 30389 26911
rect 30389 26877 30423 26911
rect 30423 26877 30432 26911
rect 30380 26868 30432 26877
rect 32956 27072 33008 27124
rect 32128 27004 32180 27056
rect 32404 27047 32456 27056
rect 32404 27013 32413 27047
rect 32413 27013 32447 27047
rect 32447 27013 32456 27047
rect 32404 27004 32456 27013
rect 33784 27004 33836 27056
rect 31484 26936 31536 26988
rect 34336 26936 34388 26988
rect 34612 26936 34664 26988
rect 36084 26936 36136 26988
rect 34060 26911 34112 26920
rect 34060 26877 34069 26911
rect 34069 26877 34103 26911
rect 34103 26877 34112 26911
rect 34060 26868 34112 26877
rect 28172 26843 28224 26852
rect 28172 26809 28181 26843
rect 28181 26809 28215 26843
rect 28215 26809 28224 26843
rect 28172 26800 28224 26809
rect 29828 26800 29880 26852
rect 25964 26775 26016 26784
rect 25964 26741 25973 26775
rect 25973 26741 26007 26775
rect 26007 26741 26016 26775
rect 25964 26732 26016 26741
rect 27160 26775 27212 26784
rect 27160 26741 27169 26775
rect 27169 26741 27203 26775
rect 27203 26741 27212 26775
rect 27160 26732 27212 26741
rect 30196 26775 30248 26784
rect 30196 26741 30205 26775
rect 30205 26741 30239 26775
rect 30239 26741 30248 26775
rect 30196 26732 30248 26741
rect 35900 26732 35952 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 22192 26528 22244 26580
rect 24492 26571 24544 26580
rect 24492 26537 24501 26571
rect 24501 26537 24535 26571
rect 24535 26537 24544 26571
rect 24492 26528 24544 26537
rect 25964 26571 26016 26580
rect 25964 26537 25973 26571
rect 25973 26537 26007 26571
rect 26007 26537 26016 26571
rect 25964 26528 26016 26537
rect 27620 26571 27672 26580
rect 27620 26537 27629 26571
rect 27629 26537 27663 26571
rect 27663 26537 27672 26571
rect 27620 26528 27672 26537
rect 28080 26528 28132 26580
rect 30196 26528 30248 26580
rect 31300 26528 31352 26580
rect 31668 26528 31720 26580
rect 21456 26460 21508 26512
rect 19340 26392 19392 26444
rect 20168 26392 20220 26444
rect 21732 26392 21784 26444
rect 20076 26367 20128 26376
rect 20076 26333 20085 26367
rect 20085 26333 20119 26367
rect 20119 26333 20128 26367
rect 20076 26324 20128 26333
rect 25872 26392 25924 26444
rect 26148 26435 26200 26444
rect 26148 26401 26157 26435
rect 26157 26401 26191 26435
rect 26191 26401 26200 26435
rect 26148 26392 26200 26401
rect 26424 26435 26476 26444
rect 26424 26401 26433 26435
rect 26433 26401 26467 26435
rect 26467 26401 26476 26435
rect 26424 26392 26476 26401
rect 24400 26367 24452 26376
rect 22468 26256 22520 26308
rect 24400 26333 24409 26367
rect 24409 26333 24443 26367
rect 24443 26333 24452 26367
rect 24400 26324 24452 26333
rect 24860 26324 24912 26376
rect 25412 26324 25464 26376
rect 26056 26324 26108 26376
rect 23756 26299 23808 26308
rect 23756 26265 23765 26299
rect 23765 26265 23799 26299
rect 23799 26265 23808 26299
rect 23756 26256 23808 26265
rect 21088 26231 21140 26240
rect 21088 26197 21097 26231
rect 21097 26197 21131 26231
rect 21131 26197 21140 26231
rect 21088 26188 21140 26197
rect 26332 26367 26384 26376
rect 26332 26333 26341 26367
rect 26341 26333 26375 26367
rect 26375 26333 26384 26367
rect 27160 26392 27212 26444
rect 26332 26324 26384 26333
rect 27068 26367 27120 26376
rect 27068 26333 27077 26367
rect 27077 26333 27111 26367
rect 27111 26333 27120 26367
rect 27068 26324 27120 26333
rect 28264 26460 28316 26512
rect 30656 26460 30708 26512
rect 27804 26392 27856 26444
rect 30196 26392 30248 26444
rect 27620 26256 27672 26308
rect 29276 26324 29328 26376
rect 29644 26324 29696 26376
rect 30380 26367 30432 26376
rect 30380 26333 30389 26367
rect 30389 26333 30423 26367
rect 30423 26333 30432 26367
rect 30380 26324 30432 26333
rect 29736 26299 29788 26308
rect 29736 26265 29745 26299
rect 29745 26265 29779 26299
rect 29779 26265 29788 26299
rect 29736 26256 29788 26265
rect 29552 26231 29604 26240
rect 29552 26197 29561 26231
rect 29561 26197 29595 26231
rect 29595 26197 29604 26231
rect 29552 26188 29604 26197
rect 31392 26367 31444 26376
rect 31392 26333 31401 26367
rect 31401 26333 31435 26367
rect 31435 26333 31444 26367
rect 32772 26528 32824 26580
rect 33784 26528 33836 26580
rect 34060 26392 34112 26444
rect 52828 26392 52880 26444
rect 31392 26324 31444 26333
rect 31760 26256 31812 26308
rect 35348 26324 35400 26376
rect 53380 26324 53432 26376
rect 33324 26256 33376 26308
rect 36084 26299 36136 26308
rect 31300 26231 31352 26240
rect 31300 26197 31309 26231
rect 31309 26197 31343 26231
rect 31343 26197 31352 26231
rect 31300 26188 31352 26197
rect 36084 26265 36093 26299
rect 36093 26265 36127 26299
rect 36127 26265 36136 26299
rect 36084 26256 36136 26265
rect 52460 26256 52512 26308
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 20076 26027 20128 26036
rect 20076 25993 20085 26027
rect 20085 25993 20119 26027
rect 20119 25993 20128 26027
rect 20076 25984 20128 25993
rect 24400 26027 24452 26036
rect 24400 25993 24409 26027
rect 24409 25993 24443 26027
rect 24443 25993 24452 26027
rect 24400 25984 24452 25993
rect 24860 26027 24912 26036
rect 24860 25993 24869 26027
rect 24869 25993 24903 26027
rect 24903 25993 24912 26027
rect 24860 25984 24912 25993
rect 26240 25984 26292 26036
rect 27068 25984 27120 26036
rect 19340 25916 19392 25968
rect 19984 25891 20036 25900
rect 19984 25857 19993 25891
rect 19993 25857 20027 25891
rect 20027 25857 20036 25891
rect 19984 25848 20036 25857
rect 19340 25644 19392 25696
rect 20168 25644 20220 25696
rect 22192 25848 22244 25900
rect 23664 25848 23716 25900
rect 24676 25848 24728 25900
rect 24584 25780 24636 25832
rect 26056 25848 26108 25900
rect 25688 25712 25740 25764
rect 26332 25848 26384 25900
rect 27160 25916 27212 25968
rect 27896 25984 27948 26036
rect 27988 25984 28040 26036
rect 30196 26027 30248 26036
rect 30196 25993 30205 26027
rect 30205 25993 30239 26027
rect 30239 25993 30248 26027
rect 30196 25984 30248 25993
rect 32772 26027 32824 26036
rect 32772 25993 32781 26027
rect 32781 25993 32815 26027
rect 32815 25993 32824 26027
rect 32772 25984 32824 25993
rect 33324 26027 33376 26036
rect 33324 25993 33333 26027
rect 33333 25993 33367 26027
rect 33367 25993 33376 26027
rect 33324 25984 33376 25993
rect 33784 26027 33836 26036
rect 33784 25993 33793 26027
rect 33793 25993 33827 26027
rect 33827 25993 33836 26027
rect 33784 25984 33836 25993
rect 34336 26027 34388 26036
rect 34336 25993 34345 26027
rect 34345 25993 34379 26027
rect 34379 25993 34388 26027
rect 34336 25984 34388 25993
rect 29368 25916 29420 25968
rect 29644 25916 29696 25968
rect 27436 25848 27488 25900
rect 27344 25823 27396 25832
rect 27344 25789 27353 25823
rect 27353 25789 27387 25823
rect 27387 25789 27396 25823
rect 27344 25780 27396 25789
rect 27620 25780 27672 25832
rect 29552 25848 29604 25900
rect 30012 25891 30064 25900
rect 29184 25780 29236 25832
rect 29644 25780 29696 25832
rect 30012 25857 30021 25891
rect 30021 25857 30055 25891
rect 30055 25857 30064 25891
rect 30012 25848 30064 25857
rect 31392 25848 31444 25900
rect 31760 25848 31812 25900
rect 32772 25848 32824 25900
rect 21088 25644 21140 25696
rect 22468 25687 22520 25696
rect 22468 25653 22477 25687
rect 22477 25653 22511 25687
rect 22511 25653 22520 25687
rect 22468 25644 22520 25653
rect 30472 25644 30524 25696
rect 32220 25687 32272 25696
rect 32220 25653 32229 25687
rect 32229 25653 32263 25687
rect 32263 25653 32272 25687
rect 32220 25644 32272 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 20076 25372 20128 25424
rect 20168 25347 20220 25356
rect 20168 25313 20177 25347
rect 20177 25313 20211 25347
rect 20211 25313 20220 25347
rect 20168 25304 20220 25313
rect 21732 25440 21784 25492
rect 24676 25483 24728 25492
rect 24676 25449 24685 25483
rect 24685 25449 24719 25483
rect 24719 25449 24728 25483
rect 24676 25440 24728 25449
rect 25596 25440 25648 25492
rect 27160 25483 27212 25492
rect 27160 25449 27169 25483
rect 27169 25449 27203 25483
rect 27203 25449 27212 25483
rect 27160 25440 27212 25449
rect 29276 25440 29328 25492
rect 29644 25483 29696 25492
rect 29644 25449 29653 25483
rect 29653 25449 29687 25483
rect 29687 25449 29696 25483
rect 29644 25440 29696 25449
rect 32220 25440 32272 25492
rect 51448 25440 51500 25492
rect 52828 25483 52880 25492
rect 52828 25449 52837 25483
rect 52837 25449 52871 25483
rect 52871 25449 52880 25483
rect 52828 25440 52880 25449
rect 27344 25372 27396 25424
rect 32772 25372 32824 25424
rect 20904 25304 20956 25356
rect 26608 25304 26660 25356
rect 19984 25236 20036 25288
rect 20812 25279 20864 25288
rect 20812 25245 20821 25279
rect 20821 25245 20855 25279
rect 20855 25245 20864 25279
rect 20812 25236 20864 25245
rect 26332 25279 26384 25288
rect 1860 25211 1912 25220
rect 1860 25177 1869 25211
rect 1869 25177 1903 25211
rect 1903 25177 1912 25211
rect 1860 25168 1912 25177
rect 16488 25100 16540 25152
rect 22192 25100 22244 25152
rect 22468 25100 22520 25152
rect 24492 25100 24544 25152
rect 26332 25245 26341 25279
rect 26341 25245 26375 25279
rect 26375 25245 26384 25279
rect 26332 25236 26384 25245
rect 30012 25304 30064 25356
rect 30472 25347 30524 25356
rect 30472 25313 30481 25347
rect 30481 25313 30515 25347
rect 30515 25313 30524 25347
rect 30472 25304 30524 25313
rect 27620 25168 27672 25220
rect 29368 25236 29420 25288
rect 29736 25279 29788 25288
rect 29736 25245 29745 25279
rect 29745 25245 29779 25279
rect 29779 25245 29788 25279
rect 29736 25236 29788 25245
rect 31300 25279 31352 25288
rect 31300 25245 31309 25279
rect 31309 25245 31343 25279
rect 31343 25245 31352 25279
rect 31300 25236 31352 25245
rect 52828 25236 52880 25288
rect 30472 25168 30524 25220
rect 28264 25143 28316 25152
rect 28264 25109 28273 25143
rect 28273 25109 28307 25143
rect 28307 25109 28316 25143
rect 28264 25100 28316 25109
rect 30748 25100 30800 25152
rect 31300 25143 31352 25152
rect 31300 25109 31309 25143
rect 31309 25109 31343 25143
rect 31343 25109 31352 25143
rect 31300 25100 31352 25109
rect 53564 25143 53616 25152
rect 53564 25109 53573 25143
rect 53573 25109 53607 25143
rect 53607 25109 53616 25143
rect 53564 25100 53616 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 1860 24896 1912 24948
rect 19984 24896 20036 24948
rect 20812 24896 20864 24948
rect 24584 24939 24636 24948
rect 24584 24905 24593 24939
rect 24593 24905 24627 24939
rect 24627 24905 24636 24939
rect 24584 24896 24636 24905
rect 25688 24896 25740 24948
rect 29368 24896 29420 24948
rect 30012 24896 30064 24948
rect 32772 24896 32824 24948
rect 20720 24828 20772 24880
rect 22192 24828 22244 24880
rect 20904 24803 20956 24812
rect 20904 24769 20913 24803
rect 20913 24769 20947 24803
rect 20947 24769 20956 24803
rect 20904 24760 20956 24769
rect 21272 24803 21324 24812
rect 21272 24769 21281 24803
rect 21281 24769 21315 24803
rect 21315 24769 21324 24803
rect 21272 24760 21324 24769
rect 22008 24803 22060 24812
rect 22008 24769 22017 24803
rect 22017 24769 22051 24803
rect 22051 24769 22060 24803
rect 22008 24760 22060 24769
rect 28264 24760 28316 24812
rect 21364 24692 21416 24744
rect 30472 24828 30524 24880
rect 31300 24828 31352 24880
rect 30748 24760 30800 24812
rect 30472 24692 30524 24744
rect 30380 24624 30432 24676
rect 19340 24599 19392 24608
rect 19340 24565 19349 24599
rect 19349 24565 19383 24599
rect 19383 24565 19392 24599
rect 19340 24556 19392 24565
rect 27620 24599 27672 24608
rect 27620 24565 27629 24599
rect 27629 24565 27663 24599
rect 27663 24565 27672 24599
rect 28080 24599 28132 24608
rect 27620 24556 27672 24565
rect 28080 24565 28089 24599
rect 28089 24565 28123 24599
rect 28123 24565 28132 24599
rect 28080 24556 28132 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 20720 24352 20772 24404
rect 21364 24395 21416 24404
rect 21364 24361 21373 24395
rect 21373 24361 21407 24395
rect 21407 24361 21416 24395
rect 21364 24352 21416 24361
rect 26332 24352 26384 24404
rect 30472 24395 30524 24404
rect 30472 24361 30481 24395
rect 30481 24361 30515 24395
rect 30515 24361 30524 24395
rect 30472 24352 30524 24361
rect 22008 24284 22060 24336
rect 27620 24216 27672 24268
rect 30104 24259 30156 24268
rect 30104 24225 30113 24259
rect 30113 24225 30147 24259
rect 30147 24225 30156 24259
rect 30104 24216 30156 24225
rect 20536 24123 20588 24132
rect 20536 24089 20545 24123
rect 20545 24089 20579 24123
rect 20579 24089 20588 24123
rect 20536 24080 20588 24089
rect 20812 24080 20864 24132
rect 30656 24012 30708 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 21272 23808 21324 23860
rect 29368 23808 29420 23860
rect 51724 23808 51776 23860
rect 19984 23468 20036 23520
rect 20536 23672 20588 23724
rect 20812 23715 20864 23724
rect 20812 23681 20821 23715
rect 20821 23681 20855 23715
rect 20855 23681 20864 23715
rect 20812 23672 20864 23681
rect 53564 23511 53616 23520
rect 53564 23477 53573 23511
rect 53573 23477 53607 23511
rect 53607 23477 53616 23511
rect 53564 23468 53616 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 20812 23264 20864 23316
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 1400 22627 1452 22636
rect 1400 22593 1409 22627
rect 1409 22593 1443 22627
rect 1443 22593 1452 22627
rect 1400 22584 1452 22593
rect 34796 22516 34848 22568
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 1400 22219 1452 22228
rect 1400 22185 1409 22219
rect 1409 22185 1443 22219
rect 1443 22185 1452 22219
rect 1400 22176 1452 22185
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 39948 21360 40000 21412
rect 53564 21335 53616 21344
rect 53564 21301 53573 21335
rect 53573 21301 53607 21335
rect 53607 21301 53616 21335
rect 53564 21292 53616 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 1400 20927 1452 20936
rect 1400 20893 1409 20927
rect 1409 20893 1443 20927
rect 1443 20893 1452 20927
rect 1400 20884 1452 20893
rect 1584 20791 1636 20800
rect 1584 20757 1593 20791
rect 1593 20757 1627 20791
rect 1627 20757 1636 20791
rect 1584 20748 1636 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 1400 20519 1452 20528
rect 1400 20485 1409 20519
rect 1409 20485 1443 20519
rect 1443 20485 1452 20519
rect 1400 20476 1452 20485
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 36084 18640 36136 18692
rect 53564 18683 53616 18692
rect 53564 18649 53573 18683
rect 53573 18649 53607 18683
rect 53607 18649 53616 18683
rect 53564 18640 53616 18649
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 1584 18232 1636 18284
rect 33140 18028 33192 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 1584 17799 1636 17808
rect 1584 17765 1593 17799
rect 1593 17765 1627 17799
rect 1627 17765 1636 17799
rect 1584 17756 1636 17765
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 30288 16600 30340 16652
rect 53564 16439 53616 16448
rect 53564 16405 53573 16439
rect 53573 16405 53607 16439
rect 53607 16405 53616 16439
rect 53564 16396 53616 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 1400 16099 1452 16108
rect 1400 16065 1409 16099
rect 1409 16065 1443 16099
rect 1443 16065 1452 16099
rect 1400 16056 1452 16065
rect 34520 15852 34572 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 1400 15691 1452 15700
rect 1400 15657 1409 15691
rect 1409 15657 1443 15691
rect 1443 15657 1452 15691
rect 1400 15648 1452 15657
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 21088 13880 21140 13932
rect 53656 13923 53708 13932
rect 53656 13889 53665 13923
rect 53665 13889 53699 13923
rect 53699 13889 53708 13923
rect 53656 13880 53708 13889
rect 42064 13812 42116 13864
rect 1492 13719 1544 13728
rect 1492 13685 1501 13719
rect 1501 13685 1535 13719
rect 1535 13685 1544 13719
rect 1492 13676 1544 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 27436 11568 27488 11620
rect 53564 11611 53616 11620
rect 53564 11577 53573 11611
rect 53573 11577 53607 11611
rect 53607 11577 53616 11611
rect 53564 11568 53616 11577
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 1584 11024 1636 11076
rect 33968 11024 34020 11076
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 1584 10795 1636 10804
rect 1584 10761 1593 10795
rect 1593 10761 1627 10795
rect 1627 10761 1636 10795
rect 1584 10752 1636 10761
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 40408 9868 40460 9920
rect 53564 9979 53616 9988
rect 53564 9945 53573 9979
rect 53573 9945 53607 9979
rect 53607 9945 53616 9979
rect 53564 9936 53616 9945
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 29460 8848 29512 8900
rect 1492 8823 1544 8832
rect 1492 8789 1501 8823
rect 1501 8789 1535 8823
rect 1535 8789 1544 8823
rect 1492 8780 1544 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 1860 7395 1912 7404
rect 1860 7361 1869 7395
rect 1869 7361 1903 7395
rect 1903 7361 1912 7395
rect 1860 7352 1912 7361
rect 53656 7395 53708 7404
rect 53656 7361 53665 7395
rect 53665 7361 53699 7395
rect 53699 7361 53708 7395
rect 53656 7352 53708 7361
rect 13636 7148 13688 7200
rect 17960 7148 18012 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 1584 6944 1636 6996
rect 1860 6944 1912 6996
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 38108 5040 38160 5092
rect 53564 5015 53616 5024
rect 53564 4981 53573 5015
rect 53573 4981 53607 5015
rect 53607 4981 53616 5015
rect 53564 4972 53616 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 15936 4564 15988 4616
rect 1492 4471 1544 4480
rect 1492 4437 1501 4471
rect 1501 4437 1535 4471
rect 1535 4437 1544 4471
rect 1492 4428 1544 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 33508 3408 33560 3460
rect 1308 3340 1360 3392
rect 1860 3340 1912 3392
rect 54116 3340 54168 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 51448 3179 51500 3188
rect 51448 3145 51457 3179
rect 51457 3145 51491 3179
rect 51491 3145 51500 3179
rect 51448 3136 51500 3145
rect 20 3000 72 3052
rect 1308 3000 1360 3052
rect 34428 2932 34480 2984
rect 13268 2864 13320 2916
rect 30564 2864 30616 2916
rect 31116 2864 31168 2916
rect 1952 2796 2004 2848
rect 2780 2839 2832 2848
rect 2780 2805 2789 2839
rect 2789 2805 2823 2839
rect 2823 2805 2832 2839
rect 2780 2796 2832 2805
rect 6460 2839 6512 2848
rect 6460 2805 6469 2839
rect 6469 2805 6503 2839
rect 6503 2805 6512 2839
rect 6460 2796 6512 2805
rect 19340 2839 19392 2848
rect 19340 2805 19349 2839
rect 19349 2805 19383 2839
rect 19383 2805 19392 2839
rect 19340 2796 19392 2805
rect 21272 2796 21324 2848
rect 22284 2796 22336 2848
rect 32220 2839 32272 2848
rect 32220 2805 32229 2839
rect 32229 2805 32263 2839
rect 32263 2805 32272 2839
rect 32220 2796 32272 2805
rect 34520 2796 34572 2848
rect 45100 2839 45152 2848
rect 45100 2805 45109 2839
rect 45109 2805 45143 2839
rect 45143 2805 45152 2839
rect 45100 2796 45152 2805
rect 47676 2796 47728 2848
rect 50344 2839 50396 2848
rect 50344 2805 50353 2839
rect 50353 2805 50387 2839
rect 50387 2805 50396 2839
rect 50344 2796 50396 2805
rect 52460 2796 52512 2848
rect 53564 2839 53616 2848
rect 53564 2805 53573 2839
rect 53573 2805 53607 2839
rect 53607 2805 53616 2839
rect 53564 2796 53616 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 21548 2592 21600 2644
rect 22192 2592 22244 2644
rect 14280 2524 14332 2576
rect 15016 2524 15068 2576
rect 2780 2431 2832 2440
rect 2780 2397 2789 2431
rect 2789 2397 2823 2431
rect 2823 2397 2832 2431
rect 2780 2388 2832 2397
rect 1860 2363 1912 2372
rect 1860 2329 1869 2363
rect 1869 2329 1903 2363
rect 1903 2329 1912 2363
rect 1860 2320 1912 2329
rect 6460 2388 6512 2440
rect 10324 2456 10376 2508
rect 19432 2524 19484 2576
rect 28172 2592 28224 2644
rect 50712 2635 50764 2644
rect 24584 2567 24636 2576
rect 16856 2456 16908 2508
rect 24584 2533 24593 2567
rect 24593 2533 24627 2567
rect 24627 2533 24636 2567
rect 24584 2524 24636 2533
rect 19984 2456 20036 2508
rect 23756 2456 23808 2508
rect 35900 2524 35952 2576
rect 36912 2524 36964 2576
rect 41512 2524 41564 2576
rect 50712 2601 50721 2635
rect 50721 2601 50755 2635
rect 50755 2601 50764 2635
rect 50712 2592 50764 2601
rect 30656 2499 30708 2508
rect 30656 2465 30665 2499
rect 30665 2465 30699 2499
rect 30699 2465 30708 2499
rect 30656 2456 30708 2465
rect 13268 2431 13320 2440
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 13268 2388 13320 2397
rect 14832 2388 14884 2440
rect 16304 2320 16356 2372
rect 19340 2388 19392 2440
rect 22284 2431 22336 2440
rect 22284 2397 22293 2431
rect 22293 2397 22327 2431
rect 22327 2397 22336 2431
rect 22284 2388 22336 2397
rect 30288 2388 30340 2440
rect 32220 2388 32272 2440
rect 25780 2320 25832 2372
rect 27712 2320 27764 2372
rect 35348 2388 35400 2440
rect 37740 2388 37792 2440
rect 38660 2388 38712 2440
rect 34520 2320 34572 2372
rect 41236 2320 41288 2372
rect 45100 2388 45152 2440
rect 49700 2388 49752 2440
rect 50344 2388 50396 2440
rect 51448 2388 51500 2440
rect 47676 2320 47728 2372
rect 52460 2320 52512 2372
rect 53564 2363 53616 2372
rect 53564 2329 53573 2363
rect 53573 2329 53607 2363
rect 53607 2329 53616 2363
rect 53564 2320 53616 2329
rect 3884 2252 3936 2304
rect 4804 2295 4856 2304
rect 4804 2261 4813 2295
rect 4813 2261 4847 2295
rect 4847 2261 4856 2295
rect 4804 2252 4856 2261
rect 8392 2295 8444 2304
rect 8392 2261 8401 2295
rect 8401 2261 8435 2295
rect 8435 2261 8444 2295
rect 8392 2252 8444 2261
rect 9128 2295 9180 2304
rect 9128 2261 9137 2295
rect 9137 2261 9171 2295
rect 9171 2261 9180 2295
rect 9128 2252 9180 2261
rect 12900 2252 12952 2304
rect 16764 2252 16816 2304
rect 17684 2295 17736 2304
rect 17684 2261 17693 2295
rect 17693 2261 17727 2295
rect 17727 2261 17736 2295
rect 17684 2252 17736 2261
rect 23848 2295 23900 2304
rect 23848 2261 23857 2295
rect 23857 2261 23891 2295
rect 23891 2261 23900 2295
rect 23848 2252 23900 2261
rect 36728 2252 36780 2304
rect 42800 2295 42852 2304
rect 42800 2261 42809 2295
rect 42809 2261 42843 2295
rect 42843 2261 42852 2295
rect 42800 2252 42852 2261
rect 43168 2252 43220 2304
rect 45376 2295 45428 2304
rect 45376 2261 45385 2295
rect 45385 2261 45419 2295
rect 45419 2261 45428 2295
rect 45376 2252 45428 2261
rect 48136 2295 48188 2304
rect 48136 2261 48145 2295
rect 48145 2261 48179 2295
rect 48179 2261 48188 2295
rect 48136 2252 48188 2261
rect 51540 2252 51592 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 4804 1980 4856 2032
rect 22468 1980 22520 2032
rect 28356 1980 28408 2032
rect 42800 1980 42852 2032
rect 17684 1912 17736 1964
rect 26792 1912 26844 1964
rect 24952 1844 25004 1896
rect 48136 1844 48188 1896
<< metal2 >>
rect 1306 56841 1362 57641
rect 1582 57216 1638 57225
rect 1582 57151 1638 57160
rect 1320 54262 1348 56841
rect 1596 55214 1624 57151
rect 3882 56841 3938 57641
rect 5814 56841 5870 57641
rect 7746 56841 7802 57641
rect 10322 56841 10378 57641
rect 12254 56841 12310 57641
rect 14186 56841 14242 57641
rect 16762 56841 16818 57641
rect 18694 56841 18750 57641
rect 21270 56841 21326 57641
rect 23202 56841 23258 57641
rect 25134 56841 25190 57641
rect 27710 56841 27766 57641
rect 29642 56841 29698 57641
rect 31574 56841 31630 57641
rect 34150 56841 34206 57641
rect 34256 56902 34468 56930
rect 1412 55186 1624 55214
rect 1412 54670 1440 55186
rect 3896 54738 3924 56841
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 5828 54874 5856 56841
rect 5816 54868 5868 54874
rect 5816 54810 5868 54816
rect 3884 54732 3936 54738
rect 3884 54674 3936 54680
rect 1400 54664 1452 54670
rect 1400 54606 1452 54612
rect 1676 54664 1728 54670
rect 1676 54606 1728 54612
rect 1308 54256 1360 54262
rect 1308 54198 1360 54204
rect 1320 53786 1348 54198
rect 1308 53780 1360 53786
rect 1308 53722 1360 53728
rect 1412 53242 1440 54606
rect 1400 53236 1452 53242
rect 1400 53178 1452 53184
rect 1400 52488 1452 52494
rect 1398 52456 1400 52465
rect 1452 52456 1454 52465
rect 1398 52391 1454 52400
rect 1412 52154 1440 52391
rect 1400 52148 1452 52154
rect 1400 52090 1452 52096
rect 1400 50924 1452 50930
rect 1400 50866 1452 50872
rect 1412 50454 1440 50866
rect 1400 50448 1452 50454
rect 1398 50416 1400 50425
rect 1452 50416 1454 50425
rect 1398 50351 1454 50360
rect 1492 48000 1544 48006
rect 1492 47942 1544 47948
rect 1504 47705 1532 47942
rect 1490 47696 1546 47705
rect 1490 47631 1546 47640
rect 1584 45892 1636 45898
rect 1584 45834 1636 45840
rect 1596 45665 1624 45834
rect 1582 45656 1638 45665
rect 1582 45591 1584 45600
rect 1636 45591 1638 45600
rect 1584 45562 1636 45568
rect 1688 44198 1716 54606
rect 2780 54596 2832 54602
rect 2780 54538 2832 54544
rect 2792 54505 2820 54538
rect 2872 54528 2924 54534
rect 2778 54496 2834 54505
rect 2872 54470 2924 54476
rect 2778 54431 2834 54440
rect 2792 54330 2820 54431
rect 2780 54324 2832 54330
rect 2780 54266 2832 54272
rect 2136 54052 2188 54058
rect 2136 53994 2188 54000
rect 1952 52624 2004 52630
rect 1952 52566 2004 52572
rect 1768 50720 1820 50726
rect 1768 50662 1820 50668
rect 1676 44192 1728 44198
rect 1676 44134 1728 44140
rect 1584 43716 1636 43722
rect 1584 43658 1636 43664
rect 1596 43625 1624 43658
rect 1582 43616 1638 43625
rect 1582 43551 1638 43560
rect 1596 43450 1624 43551
rect 1584 43444 1636 43450
rect 1584 43386 1636 43392
rect 1780 42809 1808 50662
rect 1766 42800 1822 42809
rect 1766 42735 1822 42744
rect 1492 40928 1544 40934
rect 1490 40896 1492 40905
rect 1544 40896 1546 40905
rect 1490 40831 1546 40840
rect 1584 38956 1636 38962
rect 1584 38898 1636 38904
rect 1596 38865 1624 38898
rect 1582 38856 1638 38865
rect 1582 38791 1638 38800
rect 1596 38554 1624 38791
rect 1584 38548 1636 38554
rect 1584 38490 1636 38496
rect 1858 36136 1914 36145
rect 1858 36071 1860 36080
rect 1912 36071 1914 36080
rect 1860 36042 1912 36048
rect 1872 35834 1900 36042
rect 1860 35828 1912 35834
rect 1860 35770 1912 35776
rect 1964 35193 1992 52566
rect 2148 47954 2176 53994
rect 2226 48104 2282 48113
rect 2226 48039 2228 48048
rect 2280 48039 2282 48048
rect 2228 48010 2280 48016
rect 2148 47926 2268 47954
rect 2136 45892 2188 45898
rect 2136 45834 2188 45840
rect 1950 35184 2006 35193
rect 1950 35119 2006 35128
rect 1584 34604 1636 34610
rect 1584 34546 1636 34552
rect 1596 34134 1624 34546
rect 2044 34536 2096 34542
rect 2044 34478 2096 34484
rect 1584 34128 1636 34134
rect 1582 34096 1584 34105
rect 1636 34096 1638 34105
rect 1582 34031 1638 34040
rect 2056 33114 2084 34478
rect 2044 33108 2096 33114
rect 2044 33050 2096 33056
rect 1492 32224 1544 32230
rect 1492 32166 1544 32172
rect 1504 32065 1532 32166
rect 1490 32056 1546 32065
rect 1490 31991 1546 32000
rect 2148 30598 2176 45834
rect 2240 31890 2268 47926
rect 2884 42566 2912 54470
rect 3896 54330 3924 54674
rect 7760 54670 7788 56841
rect 10336 54738 10364 56841
rect 10324 54732 10376 54738
rect 10324 54674 10376 54680
rect 10968 54732 11020 54738
rect 10968 54674 11020 54680
rect 6644 54664 6696 54670
rect 6644 54606 6696 54612
rect 7748 54664 7800 54670
rect 7748 54606 7800 54612
rect 10692 54664 10744 54670
rect 10692 54606 10744 54612
rect 6656 54330 6684 54606
rect 8024 54528 8076 54534
rect 8024 54470 8076 54476
rect 3884 54324 3936 54330
rect 3884 54266 3936 54272
rect 6644 54324 6696 54330
rect 6644 54266 6696 54272
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 2872 42560 2924 42566
rect 2872 42502 2924 42508
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 8036 41177 8064 54470
rect 10704 43994 10732 54606
rect 10980 54330 11008 54674
rect 12268 54670 12296 56841
rect 14200 54874 14228 56841
rect 14188 54868 14240 54874
rect 14188 54810 14240 54816
rect 14648 54800 14700 54806
rect 14648 54742 14700 54748
rect 12256 54664 12308 54670
rect 12256 54606 12308 54612
rect 14660 54602 14688 54742
rect 14648 54596 14700 54602
rect 14648 54538 14700 54544
rect 16776 54534 16804 56841
rect 18708 54670 18736 56841
rect 21284 54670 21312 56841
rect 22192 54800 22244 54806
rect 22192 54742 22244 54748
rect 22376 54800 22428 54806
rect 22376 54742 22428 54748
rect 18696 54664 18748 54670
rect 18696 54606 18748 54612
rect 21272 54664 21324 54670
rect 21272 54606 21324 54612
rect 15108 54528 15160 54534
rect 15108 54470 15160 54476
rect 16764 54528 16816 54534
rect 16764 54470 16816 54476
rect 18880 54528 18932 54534
rect 18880 54470 18932 54476
rect 10968 54324 11020 54330
rect 10968 54266 11020 54272
rect 15120 54126 15148 54470
rect 15108 54120 15160 54126
rect 15108 54062 15160 54068
rect 18892 51074 18920 54470
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 22204 54262 22232 54742
rect 22284 54596 22336 54602
rect 22284 54538 22336 54544
rect 22296 54330 22324 54538
rect 22284 54324 22336 54330
rect 22284 54266 22336 54272
rect 22192 54256 22244 54262
rect 22192 54198 22244 54204
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 22388 51074 22416 54742
rect 23216 54670 23244 56841
rect 25148 54874 25176 56841
rect 24676 54868 24728 54874
rect 24676 54810 24728 54816
rect 25136 54868 25188 54874
rect 25136 54810 25188 54816
rect 23204 54664 23256 54670
rect 23204 54606 23256 54612
rect 23216 54330 23244 54606
rect 24032 54528 24084 54534
rect 24032 54470 24084 54476
rect 23204 54324 23256 54330
rect 23204 54266 23256 54272
rect 24044 53106 24072 54470
rect 24688 54330 24716 54810
rect 25148 54754 25176 54810
rect 25148 54726 25268 54754
rect 27724 54738 27752 56841
rect 29656 54874 29684 56841
rect 29644 54868 29696 54874
rect 29644 54810 29696 54816
rect 25240 54670 25268 54726
rect 27712 54732 27764 54738
rect 27712 54674 27764 54680
rect 25228 54664 25280 54670
rect 25228 54606 25280 54612
rect 27896 54664 27948 54670
rect 27896 54606 27948 54612
rect 28172 54664 28224 54670
rect 28172 54606 28224 54612
rect 30472 54664 30524 54670
rect 30472 54606 30524 54612
rect 24860 54596 24912 54602
rect 24860 54538 24912 54544
rect 24676 54324 24728 54330
rect 24676 54266 24728 54272
rect 24872 53990 24900 54538
rect 24860 53984 24912 53990
rect 24860 53926 24912 53932
rect 25964 53984 26016 53990
rect 25964 53926 26016 53932
rect 26976 53984 27028 53990
rect 26976 53926 27028 53932
rect 24492 53440 24544 53446
rect 24492 53382 24544 53388
rect 24504 53242 24532 53382
rect 24492 53236 24544 53242
rect 24492 53178 24544 53184
rect 24032 53100 24084 53106
rect 24032 53042 24084 53048
rect 23848 52896 23900 52902
rect 23848 52838 23900 52844
rect 23860 52494 23888 52838
rect 24044 52630 24072 53042
rect 24032 52624 24084 52630
rect 24032 52566 24084 52572
rect 23480 52488 23532 52494
rect 23480 52430 23532 52436
rect 23848 52488 23900 52494
rect 23848 52430 23900 52436
rect 23492 52086 23520 52430
rect 23848 52352 23900 52358
rect 23848 52294 23900 52300
rect 23480 52080 23532 52086
rect 23480 52022 23532 52028
rect 23756 52080 23808 52086
rect 23756 52022 23808 52028
rect 23572 52012 23624 52018
rect 23572 51954 23624 51960
rect 23664 52012 23716 52018
rect 23664 51954 23716 51960
rect 23204 51944 23256 51950
rect 23204 51886 23256 51892
rect 22836 51808 22888 51814
rect 22836 51750 22888 51756
rect 22848 51610 22876 51750
rect 23216 51610 23244 51886
rect 22652 51604 22704 51610
rect 22652 51546 22704 51552
rect 22836 51604 22888 51610
rect 22836 51546 22888 51552
rect 23204 51604 23256 51610
rect 23204 51546 23256 51552
rect 22560 51332 22612 51338
rect 22560 51274 22612 51280
rect 18892 51046 19012 51074
rect 18880 46368 18932 46374
rect 18880 46310 18932 46316
rect 18892 46034 18920 46310
rect 18880 46028 18932 46034
rect 18880 45970 18932 45976
rect 17500 45824 17552 45830
rect 17500 45766 17552 45772
rect 16948 45076 17000 45082
rect 16948 45018 17000 45024
rect 17316 45076 17368 45082
rect 17316 45018 17368 45024
rect 16856 44872 16908 44878
rect 16856 44814 16908 44820
rect 16304 44804 16356 44810
rect 16304 44746 16356 44752
rect 15292 44736 15344 44742
rect 15292 44678 15344 44684
rect 15108 44396 15160 44402
rect 15108 44338 15160 44344
rect 14096 44192 14148 44198
rect 14096 44134 14148 44140
rect 14464 44192 14516 44198
rect 14464 44134 14516 44140
rect 15016 44192 15068 44198
rect 15016 44134 15068 44140
rect 10692 43988 10744 43994
rect 10692 43930 10744 43936
rect 14108 43382 14136 44134
rect 14476 43858 14504 44134
rect 14464 43852 14516 43858
rect 14464 43794 14516 43800
rect 14476 43654 14504 43794
rect 14740 43784 14792 43790
rect 14740 43726 14792 43732
rect 14924 43784 14976 43790
rect 14924 43726 14976 43732
rect 14464 43648 14516 43654
rect 14464 43590 14516 43596
rect 14096 43376 14148 43382
rect 14096 43318 14148 43324
rect 14108 42906 14136 43318
rect 14752 43314 14780 43726
rect 14936 43450 14964 43726
rect 14924 43444 14976 43450
rect 14924 43386 14976 43392
rect 14280 43308 14332 43314
rect 14280 43250 14332 43256
rect 14740 43308 14792 43314
rect 14740 43250 14792 43256
rect 14096 42900 14148 42906
rect 14096 42842 14148 42848
rect 14108 42702 14136 42842
rect 14292 42702 14320 43250
rect 14752 42906 14780 43250
rect 14740 42900 14792 42906
rect 14740 42842 14792 42848
rect 14096 42696 14148 42702
rect 14096 42638 14148 42644
rect 14280 42696 14332 42702
rect 14280 42638 14332 42644
rect 13636 42628 13688 42634
rect 13636 42570 13688 42576
rect 13648 42226 13676 42570
rect 13636 42220 13688 42226
rect 13636 42162 13688 42168
rect 13648 42022 13676 42162
rect 14292 42022 14320 42638
rect 14924 42628 14976 42634
rect 14924 42570 14976 42576
rect 14936 42226 14964 42570
rect 14924 42220 14976 42226
rect 14924 42162 14976 42168
rect 13636 42016 13688 42022
rect 13636 41958 13688 41964
rect 14280 42016 14332 42022
rect 14280 41958 14332 41964
rect 13648 41818 13676 41958
rect 13636 41812 13688 41818
rect 13636 41754 13688 41760
rect 8022 41168 8078 41177
rect 8022 41103 8078 41112
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 2228 31884 2280 31890
rect 2228 31826 2280 31832
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 2136 30592 2188 30598
rect 2136 30534 2188 30540
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 1400 29640 1452 29646
rect 1400 29582 1452 29588
rect 1412 29345 1440 29582
rect 1398 29336 1454 29345
rect 1398 29271 1400 29280
rect 1452 29271 1454 29280
rect 1400 29242 1452 29248
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 1492 27328 1544 27334
rect 1490 27296 1492 27305
rect 1544 27296 1546 27305
rect 1490 27231 1546 27240
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 1858 25256 1914 25265
rect 1858 25191 1860 25200
rect 1912 25191 1914 25200
rect 1860 25162 1912 25168
rect 1872 24954 1900 25162
rect 1860 24948 1912 24954
rect 1860 24890 1912 24896
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 1400 22636 1452 22642
rect 1400 22578 1452 22584
rect 1412 22545 1440 22578
rect 1398 22536 1454 22545
rect 1398 22471 1454 22480
rect 1412 22234 1440 22471
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 1400 22228 1452 22234
rect 1400 22170 1452 22176
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 1400 20936 1452 20942
rect 1400 20878 1452 20884
rect 1582 20904 1638 20913
rect 1412 20534 1440 20878
rect 1582 20839 1638 20848
rect 1596 20806 1624 20839
rect 1584 20800 1636 20806
rect 1584 20742 1636 20748
rect 1400 20528 1452 20534
rect 1398 20496 1400 20505
rect 1452 20496 1454 20505
rect 1398 20431 1454 20440
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 1584 18284 1636 18290
rect 1584 18226 1636 18232
rect 1596 17814 1624 18226
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 1584 17808 1636 17814
rect 1582 17776 1584 17785
rect 1636 17776 1638 17785
rect 1582 17711 1638 17720
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1412 15745 1440 16050
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 1398 15736 1454 15745
rect 4214 15739 4522 15748
rect 1398 15671 1400 15680
rect 1452 15671 1454 15680
rect 1400 15642 1452 15648
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 1492 13728 1544 13734
rect 1490 13696 1492 13705
rect 1544 13696 1546 13705
rect 1490 13631 1546 13640
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 1584 11076 1636 11082
rect 1584 11018 1636 11024
rect 1596 10985 1624 11018
rect 1582 10976 1638 10985
rect 1582 10911 1638 10920
rect 1596 10810 1624 10911
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 1490 8936 1546 8945
rect 1490 8871 1546 8880
rect 1504 8838 1532 8871
rect 1492 8832 1544 8838
rect 1492 8774 1544 8780
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 1872 7002 1900 7346
rect 13648 7206 13676 41754
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1860 6996 1912 7002
rect 1860 6938 1912 6944
rect 1596 6905 1624 6938
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 1492 4480 1544 4486
rect 1492 4422 1544 4428
rect 1504 4185 1532 4422
rect 1490 4176 1546 4185
rect 1490 4111 1546 4120
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 1308 3392 1360 3398
rect 1308 3334 1360 3340
rect 1860 3392 1912 3398
rect 1860 3334 1912 3340
rect 1320 3058 1348 3334
rect 20 3052 72 3058
rect 20 2994 72 3000
rect 1308 3052 1360 3058
rect 1308 2994 1360 3000
rect 32 800 60 2994
rect 1872 2378 1900 3334
rect 13268 2916 13320 2922
rect 13268 2858 13320 2864
rect 1952 2848 2004 2854
rect 1952 2790 2004 2796
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 1860 2372 1912 2378
rect 1860 2314 1912 2320
rect 1872 2145 1900 2314
rect 1858 2136 1914 2145
rect 1858 2071 1914 2080
rect 1964 800 1992 2790
rect 2792 2446 2820 2790
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 6472 2446 6500 2790
rect 10324 2508 10376 2514
rect 10324 2450 10376 2456
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 9126 2408 9182 2417
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 4804 2304 4856 2310
rect 4804 2246 4856 2252
rect 3896 800 3924 2246
rect 4816 2038 4844 2246
rect 4804 2032 4856 2038
rect 4804 1974 4856 1980
rect 6472 800 6500 2382
rect 9126 2343 9182 2352
rect 9140 2310 9168 2343
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 8404 800 8432 2246
rect 10336 800 10364 2450
rect 13280 2446 13308 2858
rect 14292 2582 14320 41958
rect 15028 2582 15056 44134
rect 15120 42770 15148 44338
rect 15304 43994 15332 44678
rect 15752 44396 15804 44402
rect 15752 44338 15804 44344
rect 15292 43988 15344 43994
rect 15292 43930 15344 43936
rect 15304 43790 15332 43930
rect 15292 43784 15344 43790
rect 15292 43726 15344 43732
rect 15384 43648 15436 43654
rect 15384 43590 15436 43596
rect 15108 42764 15160 42770
rect 15108 42706 15160 42712
rect 15396 42634 15424 43590
rect 15764 43246 15792 44338
rect 16316 43858 16344 44746
rect 16868 43926 16896 44814
rect 16960 44402 16988 45018
rect 17224 45008 17276 45014
rect 17224 44950 17276 44956
rect 17132 44804 17184 44810
rect 17132 44746 17184 44752
rect 17144 44402 17172 44746
rect 16948 44396 17000 44402
rect 16948 44338 17000 44344
rect 17132 44396 17184 44402
rect 17132 44338 17184 44344
rect 17040 44260 17092 44266
rect 17040 44202 17092 44208
rect 16856 43920 16908 43926
rect 16856 43862 16908 43868
rect 16304 43852 16356 43858
rect 16304 43794 16356 43800
rect 16316 43722 16344 43794
rect 16304 43716 16356 43722
rect 16304 43658 16356 43664
rect 16868 43314 16896 43862
rect 17052 43790 17080 44202
rect 17144 44198 17172 44338
rect 17132 44192 17184 44198
rect 17132 44134 17184 44140
rect 17040 43784 17092 43790
rect 17040 43726 17092 43732
rect 16948 43444 17000 43450
rect 16948 43386 17000 43392
rect 16856 43308 16908 43314
rect 16856 43250 16908 43256
rect 15752 43240 15804 43246
rect 15752 43182 15804 43188
rect 15384 42628 15436 42634
rect 15384 42570 15436 42576
rect 15396 42294 15424 42570
rect 15764 42566 15792 43182
rect 16764 43172 16816 43178
rect 16764 43114 16816 43120
rect 16672 43104 16724 43110
rect 16672 43046 16724 43052
rect 16684 42770 16712 43046
rect 16672 42764 16724 42770
rect 16672 42706 16724 42712
rect 15752 42560 15804 42566
rect 15752 42502 15804 42508
rect 15764 42362 15792 42502
rect 16684 42362 16712 42706
rect 16776 42702 16804 43114
rect 16868 42906 16896 43250
rect 16856 42900 16908 42906
rect 16856 42842 16908 42848
rect 16764 42696 16816 42702
rect 16764 42638 16816 42644
rect 15752 42356 15804 42362
rect 15752 42298 15804 42304
rect 16672 42356 16724 42362
rect 16672 42298 16724 42304
rect 15384 42288 15436 42294
rect 15384 42230 15436 42236
rect 16212 42288 16264 42294
rect 16212 42230 16264 42236
rect 16224 42106 16252 42230
rect 16040 42090 16252 42106
rect 16028 42084 16252 42090
rect 16080 42078 16252 42084
rect 16028 42026 16080 42032
rect 16960 41818 16988 43386
rect 17052 43314 17080 43726
rect 17040 43308 17092 43314
rect 17144 43296 17172 44134
rect 17236 43858 17264 44950
rect 17224 43852 17276 43858
rect 17224 43794 17276 43800
rect 17328 43382 17356 45018
rect 17512 44878 17540 45766
rect 18696 45484 18748 45490
rect 18696 45426 18748 45432
rect 17776 45416 17828 45422
rect 17776 45358 17828 45364
rect 17788 45082 17816 45358
rect 18052 45280 18104 45286
rect 18052 45222 18104 45228
rect 17776 45076 17828 45082
rect 17776 45018 17828 45024
rect 17500 44872 17552 44878
rect 17500 44814 17552 44820
rect 17592 44736 17644 44742
rect 17592 44678 17644 44684
rect 17868 44736 17920 44742
rect 17868 44678 17920 44684
rect 17500 44396 17552 44402
rect 17500 44338 17552 44344
rect 17512 43926 17540 44338
rect 17500 43920 17552 43926
rect 17500 43862 17552 43868
rect 17408 43648 17460 43654
rect 17408 43590 17460 43596
rect 17316 43376 17368 43382
rect 17316 43318 17368 43324
rect 17224 43308 17276 43314
rect 17144 43268 17224 43296
rect 17040 43250 17092 43256
rect 17224 43250 17276 43256
rect 17052 42226 17080 43250
rect 17132 42764 17184 42770
rect 17132 42706 17184 42712
rect 17144 42362 17172 42706
rect 17236 42702 17264 43250
rect 17224 42696 17276 42702
rect 17224 42638 17276 42644
rect 17316 42560 17368 42566
rect 17316 42502 17368 42508
rect 17132 42356 17184 42362
rect 17132 42298 17184 42304
rect 17040 42220 17092 42226
rect 17040 42162 17092 42168
rect 16948 41812 17000 41818
rect 16948 41754 17000 41760
rect 17132 41540 17184 41546
rect 17132 41482 17184 41488
rect 16028 41472 16080 41478
rect 16028 41414 16080 41420
rect 16040 41274 16068 41414
rect 16028 41268 16080 41274
rect 16028 41210 16080 41216
rect 16040 40730 16068 41210
rect 16948 40996 17000 41002
rect 16948 40938 17000 40944
rect 16672 40928 16724 40934
rect 16672 40870 16724 40876
rect 16028 40724 16080 40730
rect 16028 40666 16080 40672
rect 16580 40724 16632 40730
rect 16580 40666 16632 40672
rect 16040 40390 16068 40666
rect 16028 40384 16080 40390
rect 16028 40326 16080 40332
rect 15476 39500 15528 39506
rect 15476 39442 15528 39448
rect 15488 39302 15516 39442
rect 16304 39364 16356 39370
rect 16304 39306 16356 39312
rect 15476 39296 15528 39302
rect 15476 39238 15528 39244
rect 15936 39296 15988 39302
rect 15936 39238 15988 39244
rect 15384 38752 15436 38758
rect 15384 38694 15436 38700
rect 15396 32026 15424 38694
rect 15488 38350 15516 39238
rect 15948 39098 15976 39238
rect 15936 39092 15988 39098
rect 15936 39034 15988 39040
rect 15948 38962 15976 39034
rect 15936 38956 15988 38962
rect 15936 38898 15988 38904
rect 15476 38344 15528 38350
rect 15476 38286 15528 38292
rect 16316 38282 16344 39306
rect 16304 38276 16356 38282
rect 16304 38218 16356 38224
rect 16488 38276 16540 38282
rect 16488 38218 16540 38224
rect 16316 38010 16344 38218
rect 16396 38208 16448 38214
rect 16396 38150 16448 38156
rect 16304 38004 16356 38010
rect 16304 37946 16356 37952
rect 16028 37664 16080 37670
rect 16028 37606 16080 37612
rect 16040 37330 16068 37606
rect 16028 37324 16080 37330
rect 16028 37266 16080 37272
rect 15476 36032 15528 36038
rect 15476 35974 15528 35980
rect 15488 34746 15516 35974
rect 15936 35488 15988 35494
rect 15936 35430 15988 35436
rect 15948 34950 15976 35430
rect 15936 34944 15988 34950
rect 15936 34886 15988 34892
rect 15476 34740 15528 34746
rect 15476 34682 15528 34688
rect 15488 34474 15516 34682
rect 15476 34468 15528 34474
rect 15476 34410 15528 34416
rect 15384 32020 15436 32026
rect 15384 31962 15436 31968
rect 15948 4622 15976 34886
rect 16040 32434 16068 37266
rect 16028 32428 16080 32434
rect 16028 32370 16080 32376
rect 16028 31884 16080 31890
rect 16028 31826 16080 31832
rect 16040 31482 16068 31826
rect 16028 31476 16080 31482
rect 16028 31418 16080 31424
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 14280 2576 14332 2582
rect 14280 2518 14332 2524
rect 15016 2576 15068 2582
rect 15016 2518 15068 2524
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 12912 800 12940 2246
rect 14844 800 14872 2382
rect 16316 2378 16344 37946
rect 16408 37466 16436 38150
rect 16396 37460 16448 37466
rect 16396 37402 16448 37408
rect 16396 36100 16448 36106
rect 16396 36042 16448 36048
rect 16408 35494 16436 36042
rect 16396 35488 16448 35494
rect 16396 35430 16448 35436
rect 16396 34468 16448 34474
rect 16396 34410 16448 34416
rect 16408 33522 16436 34410
rect 16396 33516 16448 33522
rect 16396 33458 16448 33464
rect 16396 31952 16448 31958
rect 16396 31894 16448 31900
rect 16408 31822 16436 31894
rect 16396 31816 16448 31822
rect 16396 31758 16448 31764
rect 16500 25158 16528 38218
rect 16592 27402 16620 40666
rect 16684 40662 16712 40870
rect 16960 40662 16988 40938
rect 17144 40730 17172 41482
rect 17132 40724 17184 40730
rect 17132 40666 17184 40672
rect 16672 40656 16724 40662
rect 16672 40598 16724 40604
rect 16948 40656 17000 40662
rect 16948 40598 17000 40604
rect 16764 40180 16816 40186
rect 16764 40122 16816 40128
rect 16776 39438 16804 40122
rect 16948 40112 17000 40118
rect 16948 40054 17000 40060
rect 16960 39438 16988 40054
rect 17328 39846 17356 42502
rect 17420 42226 17448 43590
rect 17512 43246 17540 43862
rect 17604 43790 17632 44678
rect 17684 44192 17736 44198
rect 17684 44134 17736 44140
rect 17696 43858 17724 44134
rect 17684 43852 17736 43858
rect 17684 43794 17736 43800
rect 17592 43784 17644 43790
rect 17592 43726 17644 43732
rect 17604 43450 17632 43726
rect 17592 43444 17644 43450
rect 17592 43386 17644 43392
rect 17696 43382 17724 43794
rect 17880 43722 17908 44678
rect 18064 44334 18092 45222
rect 18328 44804 18380 44810
rect 18328 44746 18380 44752
rect 18052 44328 18104 44334
rect 18052 44270 18104 44276
rect 17868 43716 17920 43722
rect 17868 43658 17920 43664
rect 17776 43648 17828 43654
rect 17776 43590 17828 43596
rect 17684 43376 17736 43382
rect 17684 43318 17736 43324
rect 17500 43240 17552 43246
rect 17500 43182 17552 43188
rect 17592 43172 17644 43178
rect 17592 43114 17644 43120
rect 17604 42634 17632 43114
rect 17696 42906 17724 43318
rect 17684 42900 17736 42906
rect 17684 42842 17736 42848
rect 17788 42786 17816 43590
rect 17696 42758 17816 42786
rect 17880 43296 17908 43658
rect 17960 43308 18012 43314
rect 17880 43268 17960 43296
rect 17592 42628 17644 42634
rect 17592 42570 17644 42576
rect 17408 42220 17460 42226
rect 17408 42162 17460 42168
rect 17696 42090 17724 42758
rect 17776 42696 17828 42702
rect 17776 42638 17828 42644
rect 17788 42362 17816 42638
rect 17776 42356 17828 42362
rect 17776 42298 17828 42304
rect 17684 42084 17736 42090
rect 17684 42026 17736 42032
rect 17592 41812 17644 41818
rect 17592 41754 17644 41760
rect 17604 41070 17632 41754
rect 17788 41614 17816 42298
rect 17880 42226 17908 43268
rect 17960 43250 18012 43256
rect 18064 43246 18092 44270
rect 18052 43240 18104 43246
rect 18052 43182 18104 43188
rect 18340 42906 18368 44746
rect 18420 44396 18472 44402
rect 18420 44338 18472 44344
rect 18512 44396 18564 44402
rect 18512 44338 18564 44344
rect 18432 43994 18460 44338
rect 18524 44198 18552 44338
rect 18604 44328 18656 44334
rect 18604 44270 18656 44276
rect 18512 44192 18564 44198
rect 18512 44134 18564 44140
rect 18420 43988 18472 43994
rect 18420 43930 18472 43936
rect 18524 43450 18552 44134
rect 18616 43994 18644 44270
rect 18708 44266 18736 45426
rect 18880 45280 18932 45286
rect 18880 45222 18932 45228
rect 18892 44334 18920 45222
rect 18880 44328 18932 44334
rect 18880 44270 18932 44276
rect 18696 44260 18748 44266
rect 18696 44202 18748 44208
rect 18604 43988 18656 43994
rect 18604 43930 18656 43936
rect 18604 43716 18656 43722
rect 18604 43658 18656 43664
rect 18512 43444 18564 43450
rect 18512 43386 18564 43392
rect 18616 43314 18644 43658
rect 18604 43308 18656 43314
rect 18604 43250 18656 43256
rect 18328 42900 18380 42906
rect 18328 42842 18380 42848
rect 18052 42560 18104 42566
rect 18052 42502 18104 42508
rect 17868 42220 17920 42226
rect 17868 42162 17920 42168
rect 17776 41608 17828 41614
rect 17776 41550 17828 41556
rect 17960 41608 18012 41614
rect 17960 41550 18012 41556
rect 17788 41414 17816 41550
rect 17696 41386 17816 41414
rect 17592 41064 17644 41070
rect 17592 41006 17644 41012
rect 17500 40928 17552 40934
rect 17500 40870 17552 40876
rect 17512 40118 17540 40870
rect 17696 40458 17724 41386
rect 17972 41274 18000 41550
rect 17960 41268 18012 41274
rect 17960 41210 18012 41216
rect 18064 41206 18092 42502
rect 18340 41818 18368 42842
rect 18892 42294 18920 44270
rect 18984 42770 19012 51046
rect 22204 51046 22416 51074
rect 22008 50720 22060 50726
rect 22008 50662 22060 50668
rect 22020 50318 22048 50662
rect 22008 50312 22060 50318
rect 22008 50254 22060 50260
rect 21640 50176 21692 50182
rect 21640 50118 21692 50124
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 21652 49842 21680 50118
rect 21640 49836 21692 49842
rect 21640 49778 21692 49784
rect 21652 49745 21680 49778
rect 22020 49774 22048 50254
rect 22008 49768 22060 49774
rect 21638 49736 21694 49745
rect 22008 49710 22060 49716
rect 21638 49671 21694 49680
rect 22020 49094 22048 49710
rect 22008 49088 22060 49094
rect 22008 49030 22060 49036
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 20168 48136 20220 48142
rect 20168 48078 20220 48084
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 20180 47666 20208 48078
rect 22020 48006 22048 49030
rect 20720 48000 20772 48006
rect 20720 47942 20772 47948
rect 22008 48000 22060 48006
rect 22008 47942 22060 47948
rect 20168 47660 20220 47666
rect 20168 47602 20220 47608
rect 20180 47462 20208 47602
rect 20732 47598 20760 47942
rect 22020 47734 22048 47942
rect 21548 47728 21600 47734
rect 21548 47670 21600 47676
rect 22008 47728 22060 47734
rect 22008 47670 22060 47676
rect 20720 47592 20772 47598
rect 20720 47534 20772 47540
rect 20732 47462 20760 47534
rect 21560 47462 21588 47670
rect 20168 47456 20220 47462
rect 20720 47456 20772 47462
rect 20168 47398 20220 47404
rect 20718 47424 20720 47433
rect 21548 47456 21600 47462
rect 20772 47424 20774 47433
rect 20180 47054 20208 47398
rect 21548 47398 21600 47404
rect 20718 47359 20774 47368
rect 20168 47048 20220 47054
rect 20168 46990 20220 46996
rect 20628 46980 20680 46986
rect 20628 46922 20680 46928
rect 19340 46912 19392 46918
rect 19340 46854 19392 46860
rect 19352 46374 19380 46854
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 19340 46368 19392 46374
rect 19340 46310 19392 46316
rect 19352 46170 19380 46310
rect 19340 46164 19392 46170
rect 19340 46106 19392 46112
rect 19248 46028 19300 46034
rect 19248 45970 19300 45976
rect 19260 45354 19288 45970
rect 19248 45348 19300 45354
rect 19248 45290 19300 45296
rect 19260 45082 19288 45290
rect 19248 45076 19300 45082
rect 19248 45018 19300 45024
rect 19260 44470 19288 45018
rect 19352 45014 19380 46106
rect 19984 45960 20036 45966
rect 19984 45902 20036 45908
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 19996 45490 20024 45902
rect 20076 45824 20128 45830
rect 20076 45766 20128 45772
rect 19984 45484 20036 45490
rect 19984 45426 20036 45432
rect 19432 45416 19484 45422
rect 19432 45358 19484 45364
rect 19444 45082 19472 45358
rect 19432 45076 19484 45082
rect 19432 45018 19484 45024
rect 19340 45008 19392 45014
rect 19340 44950 19392 44956
rect 19996 44878 20024 45426
rect 19984 44872 20036 44878
rect 19984 44814 20036 44820
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19248 44464 19300 44470
rect 19248 44406 19300 44412
rect 19996 43926 20024 44814
rect 20088 44810 20116 45766
rect 20076 44804 20128 44810
rect 20076 44746 20128 44752
rect 20088 44470 20116 44746
rect 20260 44736 20312 44742
rect 20260 44678 20312 44684
rect 20272 44470 20300 44678
rect 20076 44464 20128 44470
rect 20076 44406 20128 44412
rect 20260 44464 20312 44470
rect 20260 44406 20312 44412
rect 19984 43920 20036 43926
rect 19984 43862 20036 43868
rect 20088 43790 20116 44406
rect 20352 43920 20404 43926
rect 20352 43862 20404 43868
rect 19432 43784 19484 43790
rect 19432 43726 19484 43732
rect 20076 43784 20128 43790
rect 20076 43726 20128 43732
rect 19340 43648 19392 43654
rect 19340 43590 19392 43596
rect 19352 43450 19380 43590
rect 19340 43444 19392 43450
rect 19340 43386 19392 43392
rect 19444 43110 19472 43726
rect 19984 43716 20036 43722
rect 19984 43658 20036 43664
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19996 43382 20024 43658
rect 20076 43648 20128 43654
rect 20076 43590 20128 43596
rect 19984 43376 20036 43382
rect 19984 43318 20036 43324
rect 19432 43104 19484 43110
rect 19432 43046 19484 43052
rect 19984 43104 20036 43110
rect 19984 43046 20036 43052
rect 18972 42764 19024 42770
rect 18972 42706 19024 42712
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 18880 42288 18932 42294
rect 18880 42230 18932 42236
rect 19432 42288 19484 42294
rect 19432 42230 19484 42236
rect 18512 42016 18564 42022
rect 18512 41958 18564 41964
rect 18328 41812 18380 41818
rect 18328 41754 18380 41760
rect 18236 41608 18288 41614
rect 18236 41550 18288 41556
rect 18144 41268 18196 41274
rect 18144 41210 18196 41216
rect 18052 41200 18104 41206
rect 18052 41142 18104 41148
rect 17960 40996 18012 41002
rect 17960 40938 18012 40944
rect 17684 40452 17736 40458
rect 17684 40394 17736 40400
rect 17972 40118 18000 40938
rect 18156 40594 18184 41210
rect 18248 41138 18276 41550
rect 18236 41132 18288 41138
rect 18236 41074 18288 41080
rect 18144 40588 18196 40594
rect 18144 40530 18196 40536
rect 18052 40520 18104 40526
rect 18052 40462 18104 40468
rect 17500 40112 17552 40118
rect 17500 40054 17552 40060
rect 17960 40112 18012 40118
rect 17960 40054 18012 40060
rect 18064 39982 18092 40462
rect 18248 40458 18276 41074
rect 18524 40594 18552 41958
rect 19444 41546 19472 42230
rect 19996 42158 20024 43046
rect 20088 42702 20116 43590
rect 20364 42702 20392 43862
rect 20640 43738 20668 46922
rect 20996 46368 21048 46374
rect 20996 46310 21048 46316
rect 21008 46170 21036 46310
rect 20996 46164 21048 46170
rect 20996 46106 21048 46112
rect 20996 45960 21048 45966
rect 20996 45902 21048 45908
rect 21008 45626 21036 45902
rect 20996 45620 21048 45626
rect 20996 45562 21048 45568
rect 20720 45348 20772 45354
rect 20720 45290 20772 45296
rect 20732 43790 20760 45290
rect 21008 44946 21036 45562
rect 21364 45552 21416 45558
rect 21364 45494 21416 45500
rect 21180 45416 21232 45422
rect 21180 45358 21232 45364
rect 21088 45280 21140 45286
rect 21088 45222 21140 45228
rect 20904 44940 20956 44946
rect 20904 44882 20956 44888
rect 20996 44940 21048 44946
rect 20996 44882 21048 44888
rect 20812 44872 20864 44878
rect 20812 44814 20864 44820
rect 20824 44198 20852 44814
rect 20812 44192 20864 44198
rect 20812 44134 20864 44140
rect 20548 43710 20668 43738
rect 20720 43784 20772 43790
rect 20720 43726 20772 43732
rect 20076 42696 20128 42702
rect 20076 42638 20128 42644
rect 20352 42696 20404 42702
rect 20352 42638 20404 42644
rect 20088 42226 20116 42638
rect 20260 42628 20312 42634
rect 20260 42570 20312 42576
rect 20168 42560 20220 42566
rect 20168 42502 20220 42508
rect 20076 42220 20128 42226
rect 20076 42162 20128 42168
rect 19984 42152 20036 42158
rect 19984 42094 20036 42100
rect 20180 41682 20208 42502
rect 20272 42362 20300 42570
rect 20260 42356 20312 42362
rect 20260 42298 20312 42304
rect 20444 42356 20496 42362
rect 20444 42298 20496 42304
rect 20272 41698 20300 42298
rect 20456 42226 20484 42298
rect 20444 42220 20496 42226
rect 20444 42162 20496 42168
rect 20444 42016 20496 42022
rect 20444 41958 20496 41964
rect 20168 41676 20220 41682
rect 20272 41670 20392 41698
rect 20168 41618 20220 41624
rect 20260 41608 20312 41614
rect 20260 41550 20312 41556
rect 19432 41540 19484 41546
rect 19432 41482 19484 41488
rect 19340 41472 19392 41478
rect 19340 41414 19392 41420
rect 18604 41132 18656 41138
rect 18604 41074 18656 41080
rect 18616 40730 18644 41074
rect 18786 41032 18842 41041
rect 18786 40967 18788 40976
rect 18840 40967 18842 40976
rect 18788 40938 18840 40944
rect 18604 40724 18656 40730
rect 18604 40666 18656 40672
rect 18972 40656 19024 40662
rect 18972 40598 19024 40604
rect 18512 40588 18564 40594
rect 18512 40530 18564 40536
rect 18788 40520 18840 40526
rect 18788 40462 18840 40468
rect 18236 40452 18288 40458
rect 18236 40394 18288 40400
rect 18696 40384 18748 40390
rect 18696 40326 18748 40332
rect 18052 39976 18104 39982
rect 18052 39918 18104 39924
rect 17316 39840 17368 39846
rect 17500 39840 17552 39846
rect 17316 39782 17368 39788
rect 17420 39800 17500 39828
rect 17328 39438 17356 39782
rect 16764 39432 16816 39438
rect 16764 39374 16816 39380
rect 16948 39432 17000 39438
rect 16948 39374 17000 39380
rect 17316 39432 17368 39438
rect 17316 39374 17368 39380
rect 16776 39030 16804 39374
rect 16764 39024 16816 39030
rect 16764 38966 16816 38972
rect 16672 38956 16724 38962
rect 16672 38898 16724 38904
rect 16684 38554 16712 38898
rect 16672 38548 16724 38554
rect 16672 38490 16724 38496
rect 16960 38282 16988 39374
rect 17224 38344 17276 38350
rect 17328 38332 17356 39374
rect 17420 39370 17448 39800
rect 17500 39782 17552 39788
rect 18064 39506 18092 39918
rect 18052 39500 18104 39506
rect 18052 39442 18104 39448
rect 17776 39432 17828 39438
rect 17776 39374 17828 39380
rect 17408 39364 17460 39370
rect 17408 39306 17460 39312
rect 17420 38962 17448 39306
rect 17500 39296 17552 39302
rect 17500 39238 17552 39244
rect 17408 38956 17460 38962
rect 17408 38898 17460 38904
rect 17512 38842 17540 39238
rect 17788 39098 17816 39374
rect 17776 39092 17828 39098
rect 17776 39034 17828 39040
rect 18708 39030 18736 40326
rect 18800 39846 18828 40462
rect 18880 40452 18932 40458
rect 18880 40394 18932 40400
rect 18788 39840 18840 39846
rect 18788 39782 18840 39788
rect 18800 39506 18828 39782
rect 18788 39500 18840 39506
rect 18788 39442 18840 39448
rect 18696 39024 18748 39030
rect 18340 38972 18696 38978
rect 18340 38966 18748 38972
rect 18340 38962 18736 38966
rect 18328 38956 18736 38962
rect 18380 38950 18736 38956
rect 18328 38898 18380 38904
rect 17276 38304 17356 38332
rect 17420 38814 17540 38842
rect 17224 38286 17276 38292
rect 16948 38276 17000 38282
rect 16948 38218 17000 38224
rect 16960 37126 16988 38218
rect 17236 37262 17264 38286
rect 17420 37874 17448 38814
rect 17500 38752 17552 38758
rect 17500 38694 17552 38700
rect 17512 38350 17540 38694
rect 17500 38344 17552 38350
rect 17500 38286 17552 38292
rect 18144 38344 18196 38350
rect 18144 38286 18196 38292
rect 18328 38344 18380 38350
rect 18328 38286 18380 38292
rect 17408 37868 17460 37874
rect 17408 37810 17460 37816
rect 17316 37392 17368 37398
rect 17316 37334 17368 37340
rect 17224 37256 17276 37262
rect 17224 37198 17276 37204
rect 16948 37120 17000 37126
rect 16948 37062 17000 37068
rect 17328 36786 17356 37334
rect 17420 36802 17448 37810
rect 17512 37466 17540 38286
rect 17684 38208 17736 38214
rect 17684 38150 17736 38156
rect 17776 38208 17828 38214
rect 17776 38150 17828 38156
rect 17696 38010 17724 38150
rect 17684 38004 17736 38010
rect 17684 37946 17736 37952
rect 17500 37460 17552 37466
rect 17500 37402 17552 37408
rect 17696 36922 17724 37946
rect 17788 37874 17816 38150
rect 17776 37868 17828 37874
rect 17776 37810 17828 37816
rect 17788 37398 17816 37810
rect 17776 37392 17828 37398
rect 17776 37334 17828 37340
rect 17868 37324 17920 37330
rect 17868 37266 17920 37272
rect 17684 36916 17736 36922
rect 17684 36858 17736 36864
rect 17420 36786 17632 36802
rect 17316 36780 17368 36786
rect 17420 36780 17644 36786
rect 17420 36774 17592 36780
rect 17316 36722 17368 36728
rect 17592 36722 17644 36728
rect 17328 36174 17356 36722
rect 17604 36310 17632 36722
rect 17592 36304 17644 36310
rect 17592 36246 17644 36252
rect 17316 36168 17368 36174
rect 17316 36110 17368 36116
rect 16948 36032 17000 36038
rect 16948 35974 17000 35980
rect 17592 36032 17644 36038
rect 17592 35974 17644 35980
rect 16856 35488 16908 35494
rect 16856 35430 16908 35436
rect 16764 35080 16816 35086
rect 16764 35022 16816 35028
rect 16776 34542 16804 35022
rect 16868 34678 16896 35430
rect 16960 35154 16988 35974
rect 16948 35148 17000 35154
rect 16948 35090 17000 35096
rect 17408 35148 17460 35154
rect 17408 35090 17460 35096
rect 16960 34746 16988 35090
rect 16948 34740 17000 34746
rect 16948 34682 17000 34688
rect 16856 34672 16908 34678
rect 16856 34614 16908 34620
rect 16764 34536 16816 34542
rect 16764 34478 16816 34484
rect 16776 33862 16804 34478
rect 16868 34202 16896 34614
rect 17420 34406 17448 35090
rect 17604 35086 17632 35974
rect 17880 35154 17908 37266
rect 18156 36922 18184 38286
rect 18236 37460 18288 37466
rect 18236 37402 18288 37408
rect 18144 36916 18196 36922
rect 18144 36858 18196 36864
rect 17960 36304 18012 36310
rect 17960 36246 18012 36252
rect 17972 36038 18000 36246
rect 18156 36242 18184 36858
rect 18248 36802 18276 37402
rect 18340 37398 18368 38286
rect 18512 37936 18564 37942
rect 18432 37884 18512 37890
rect 18432 37878 18564 37884
rect 18432 37862 18552 37878
rect 18328 37392 18380 37398
rect 18328 37334 18380 37340
rect 18432 37262 18460 37862
rect 18696 37800 18748 37806
rect 18696 37742 18748 37748
rect 18512 37664 18564 37670
rect 18512 37606 18564 37612
rect 18420 37256 18472 37262
rect 18420 37198 18472 37204
rect 18248 36786 18368 36802
rect 18248 36780 18380 36786
rect 18248 36774 18328 36780
rect 18248 36310 18276 36774
rect 18328 36722 18380 36728
rect 18432 36650 18460 37198
rect 18524 37126 18552 37606
rect 18708 37262 18736 37742
rect 18696 37256 18748 37262
rect 18696 37198 18748 37204
rect 18512 37120 18564 37126
rect 18512 37062 18564 37068
rect 18524 36854 18552 37062
rect 18512 36848 18564 36854
rect 18512 36790 18564 36796
rect 18420 36644 18472 36650
rect 18420 36586 18472 36592
rect 18236 36304 18288 36310
rect 18236 36246 18288 36252
rect 18144 36236 18196 36242
rect 18144 36178 18196 36184
rect 18052 36168 18104 36174
rect 18052 36110 18104 36116
rect 17960 36032 18012 36038
rect 17960 35974 18012 35980
rect 17972 35766 18000 35974
rect 18064 35834 18092 36110
rect 18052 35828 18104 35834
rect 18052 35770 18104 35776
rect 17960 35760 18012 35766
rect 17960 35702 18012 35708
rect 18156 35494 18184 36178
rect 18524 36174 18552 36790
rect 18604 36576 18656 36582
rect 18604 36518 18656 36524
rect 18236 36168 18288 36174
rect 18236 36110 18288 36116
rect 18512 36168 18564 36174
rect 18512 36110 18564 36116
rect 18248 35630 18276 36110
rect 18616 35834 18644 36518
rect 18696 36100 18748 36106
rect 18696 36042 18748 36048
rect 18604 35828 18656 35834
rect 18604 35770 18656 35776
rect 18708 35630 18736 36042
rect 18892 35894 18920 40394
rect 18800 35866 18920 35894
rect 18236 35624 18288 35630
rect 18236 35566 18288 35572
rect 18696 35624 18748 35630
rect 18696 35566 18748 35572
rect 18144 35488 18196 35494
rect 18144 35430 18196 35436
rect 18248 35290 18276 35566
rect 18236 35284 18288 35290
rect 18236 35226 18288 35232
rect 17868 35148 17920 35154
rect 17868 35090 17920 35096
rect 17960 35148 18012 35154
rect 17960 35090 18012 35096
rect 17592 35080 17644 35086
rect 17592 35022 17644 35028
rect 17604 34610 17632 35022
rect 17592 34604 17644 34610
rect 17592 34546 17644 34552
rect 17408 34400 17460 34406
rect 17408 34342 17460 34348
rect 16856 34196 16908 34202
rect 16856 34138 16908 34144
rect 16764 33856 16816 33862
rect 16764 33798 16816 33804
rect 16580 27396 16632 27402
rect 16580 27338 16632 27344
rect 16776 26234 16804 33798
rect 17972 33114 18000 35090
rect 18052 35080 18104 35086
rect 18052 35022 18104 35028
rect 18512 35080 18564 35086
rect 18512 35022 18564 35028
rect 18064 34678 18092 35022
rect 18524 34746 18552 35022
rect 18512 34740 18564 34746
rect 18512 34682 18564 34688
rect 18052 34672 18104 34678
rect 18052 34614 18104 34620
rect 18234 34640 18290 34649
rect 18064 34202 18092 34614
rect 18234 34575 18236 34584
rect 18288 34575 18290 34584
rect 18236 34546 18288 34552
rect 18144 34400 18196 34406
rect 18144 34342 18196 34348
rect 18052 34196 18104 34202
rect 18052 34138 18104 34144
rect 18156 33998 18184 34342
rect 18248 34066 18276 34546
rect 18420 34536 18472 34542
rect 18420 34478 18472 34484
rect 18432 34134 18460 34478
rect 18420 34128 18472 34134
rect 18420 34070 18472 34076
rect 18236 34060 18288 34066
rect 18236 34002 18288 34008
rect 18144 33992 18196 33998
rect 18144 33934 18196 33940
rect 17960 33108 18012 33114
rect 17960 33050 18012 33056
rect 17972 32910 18000 33050
rect 17960 32904 18012 32910
rect 17960 32846 18012 32852
rect 16856 32768 16908 32774
rect 16856 32710 16908 32716
rect 16868 31822 16896 32710
rect 17684 32496 17736 32502
rect 17684 32438 17736 32444
rect 17696 32366 17724 32438
rect 17684 32360 17736 32366
rect 17684 32302 17736 32308
rect 17972 32230 18000 32846
rect 18156 32774 18184 33934
rect 18248 33522 18276 34002
rect 18328 33924 18380 33930
rect 18328 33866 18380 33872
rect 18340 33658 18368 33866
rect 18328 33652 18380 33658
rect 18328 33594 18380 33600
rect 18236 33516 18288 33522
rect 18236 33458 18288 33464
rect 18420 32972 18472 32978
rect 18420 32914 18472 32920
rect 18144 32768 18196 32774
rect 18144 32710 18196 32716
rect 18328 32768 18380 32774
rect 18328 32710 18380 32716
rect 18156 32586 18184 32710
rect 18064 32570 18184 32586
rect 18052 32564 18184 32570
rect 18104 32558 18184 32564
rect 18052 32506 18104 32512
rect 18052 32428 18104 32434
rect 18052 32370 18104 32376
rect 17960 32224 18012 32230
rect 17960 32166 18012 32172
rect 18064 31822 18092 32370
rect 18156 32026 18184 32558
rect 18144 32020 18196 32026
rect 18144 31962 18196 31968
rect 16856 31816 16908 31822
rect 16856 31758 16908 31764
rect 18052 31816 18104 31822
rect 18052 31758 18104 31764
rect 17960 31748 18012 31754
rect 17960 31690 18012 31696
rect 16948 31680 17000 31686
rect 16948 31622 17000 31628
rect 17224 31680 17276 31686
rect 17224 31622 17276 31628
rect 17592 31680 17644 31686
rect 17592 31622 17644 31628
rect 16960 31346 16988 31622
rect 17236 31346 17264 31622
rect 17604 31346 17632 31622
rect 17972 31346 18000 31690
rect 18064 31482 18092 31758
rect 18052 31476 18104 31482
rect 18052 31418 18104 31424
rect 16948 31340 17000 31346
rect 16948 31282 17000 31288
rect 17224 31340 17276 31346
rect 17224 31282 17276 31288
rect 17592 31340 17644 31346
rect 17592 31282 17644 31288
rect 17960 31340 18012 31346
rect 17960 31282 18012 31288
rect 16948 31136 17000 31142
rect 16948 31078 17000 31084
rect 16960 30734 16988 31078
rect 16948 30728 17000 30734
rect 16948 30670 17000 30676
rect 17236 28558 17264 31282
rect 17604 30598 17632 31282
rect 17592 30592 17644 30598
rect 17592 30534 17644 30540
rect 17972 30054 18000 31282
rect 18340 30802 18368 32710
rect 18432 32434 18460 32914
rect 18512 32904 18564 32910
rect 18512 32846 18564 32852
rect 18604 32904 18656 32910
rect 18604 32846 18656 32852
rect 18420 32428 18472 32434
rect 18420 32370 18472 32376
rect 18432 31958 18460 32370
rect 18524 32026 18552 32846
rect 18616 32570 18644 32846
rect 18604 32564 18656 32570
rect 18604 32506 18656 32512
rect 18696 32224 18748 32230
rect 18696 32166 18748 32172
rect 18512 32020 18564 32026
rect 18512 31962 18564 31968
rect 18420 31952 18472 31958
rect 18420 31894 18472 31900
rect 18432 31482 18460 31894
rect 18420 31476 18472 31482
rect 18420 31418 18472 31424
rect 18524 31346 18552 31962
rect 18708 31346 18736 32166
rect 18512 31340 18564 31346
rect 18512 31282 18564 31288
rect 18696 31340 18748 31346
rect 18696 31282 18748 31288
rect 18328 30796 18380 30802
rect 18328 30738 18380 30744
rect 17960 30048 18012 30054
rect 17960 29990 18012 29996
rect 17224 28552 17276 28558
rect 17224 28494 17276 28500
rect 16776 26206 16896 26234
rect 16488 25152 16540 25158
rect 16488 25094 16540 25100
rect 16868 2514 16896 26206
rect 17972 7206 18000 29990
rect 18144 29504 18196 29510
rect 18144 29446 18196 29452
rect 18156 29238 18184 29446
rect 18144 29232 18196 29238
rect 18144 29174 18196 29180
rect 18800 28694 18828 35866
rect 18880 35692 18932 35698
rect 18880 35634 18932 35640
rect 18892 34746 18920 35634
rect 18880 34740 18932 34746
rect 18880 34682 18932 34688
rect 18984 33658 19012 40598
rect 19352 40458 19380 41414
rect 19444 41138 19472 41482
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19432 41132 19484 41138
rect 19432 41074 19484 41080
rect 20272 40730 20300 41550
rect 20364 41546 20392 41670
rect 20456 41614 20484 41958
rect 20444 41608 20496 41614
rect 20444 41550 20496 41556
rect 20352 41540 20404 41546
rect 20352 41482 20404 41488
rect 20260 40724 20312 40730
rect 20260 40666 20312 40672
rect 19982 40624 20038 40633
rect 19432 40588 19484 40594
rect 20548 40610 20576 43710
rect 20824 43382 20852 44134
rect 20916 43994 20944 44882
rect 20996 44736 21048 44742
rect 20996 44678 21048 44684
rect 20904 43988 20956 43994
rect 20904 43930 20956 43936
rect 20812 43376 20864 43382
rect 20812 43318 20864 43324
rect 20720 42220 20772 42226
rect 20720 42162 20772 42168
rect 20628 41472 20680 41478
rect 20628 41414 20680 41420
rect 19982 40559 20038 40568
rect 20272 40582 20576 40610
rect 19432 40530 19484 40536
rect 19340 40452 19392 40458
rect 19340 40394 19392 40400
rect 19444 40050 19472 40530
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19996 40050 20024 40559
rect 19432 40044 19484 40050
rect 19432 39986 19484 39992
rect 19984 40044 20036 40050
rect 19984 39986 20036 39992
rect 19340 39432 19392 39438
rect 19340 39374 19392 39380
rect 19352 39098 19380 39374
rect 19432 39296 19484 39302
rect 19432 39238 19484 39244
rect 19340 39092 19392 39098
rect 19340 39034 19392 39040
rect 19444 38826 19472 39238
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 20168 39092 20220 39098
rect 20168 39034 20220 39040
rect 19524 38888 19576 38894
rect 19524 38830 19576 38836
rect 19432 38820 19484 38826
rect 19432 38762 19484 38768
rect 19536 38350 19564 38830
rect 20180 38350 20208 39034
rect 19248 38344 19300 38350
rect 19524 38344 19576 38350
rect 19248 38286 19300 38292
rect 19444 38304 19524 38332
rect 19260 37194 19288 38286
rect 19444 38010 19472 38304
rect 19524 38286 19576 38292
rect 20168 38344 20220 38350
rect 20168 38286 20220 38292
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19432 38004 19484 38010
rect 19432 37946 19484 37952
rect 19444 37330 19472 37946
rect 20180 37874 20208 38286
rect 20076 37868 20128 37874
rect 20076 37810 20128 37816
rect 20168 37868 20220 37874
rect 20168 37810 20220 37816
rect 19708 37664 19760 37670
rect 19708 37606 19760 37612
rect 19720 37466 19748 37606
rect 19708 37460 19760 37466
rect 19708 37402 19760 37408
rect 19432 37324 19484 37330
rect 19432 37266 19484 37272
rect 20088 37262 20116 37810
rect 20076 37256 20128 37262
rect 20076 37198 20128 37204
rect 19248 37188 19300 37194
rect 19248 37130 19300 37136
rect 19984 37188 20036 37194
rect 19984 37130 20036 37136
rect 19064 36780 19116 36786
rect 19064 36722 19116 36728
rect 19076 35222 19104 36722
rect 19260 36582 19288 37130
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19996 36922 20024 37130
rect 19984 36916 20036 36922
rect 19984 36858 20036 36864
rect 20168 36712 20220 36718
rect 20168 36654 20220 36660
rect 19248 36576 19300 36582
rect 19248 36518 19300 36524
rect 20180 36242 20208 36654
rect 20168 36236 20220 36242
rect 20168 36178 20220 36184
rect 19984 36032 20036 36038
rect 19984 35974 20036 35980
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19996 35834 20024 35974
rect 20180 35834 20208 36178
rect 19248 35828 19300 35834
rect 19248 35770 19300 35776
rect 19984 35828 20036 35834
rect 19984 35770 20036 35776
rect 20168 35828 20220 35834
rect 20168 35770 20220 35776
rect 19156 35624 19208 35630
rect 19156 35566 19208 35572
rect 19064 35216 19116 35222
rect 19064 35158 19116 35164
rect 19076 34678 19104 35158
rect 19168 34950 19196 35566
rect 19260 35494 19288 35770
rect 19248 35488 19300 35494
rect 19248 35430 19300 35436
rect 19260 35154 19288 35430
rect 19248 35148 19300 35154
rect 19248 35090 19300 35096
rect 19996 35086 20024 35770
rect 19432 35080 19484 35086
rect 19432 35022 19484 35028
rect 19984 35080 20036 35086
rect 19984 35022 20036 35028
rect 19340 35012 19392 35018
rect 19340 34954 19392 34960
rect 19156 34944 19208 34950
rect 19156 34886 19208 34892
rect 19064 34672 19116 34678
rect 19064 34614 19116 34620
rect 19352 34542 19380 34954
rect 19444 34610 19472 35022
rect 20076 34944 20128 34950
rect 20076 34886 20128 34892
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19432 34604 19484 34610
rect 19432 34546 19484 34552
rect 19340 34536 19392 34542
rect 19340 34478 19392 34484
rect 19444 34202 19472 34546
rect 19800 34536 19852 34542
rect 19800 34478 19852 34484
rect 19812 34202 19840 34478
rect 19432 34196 19484 34202
rect 19432 34138 19484 34144
rect 19800 34196 19852 34202
rect 19800 34138 19852 34144
rect 19444 33998 19472 34138
rect 20088 34066 20116 34886
rect 20076 34060 20128 34066
rect 20076 34002 20128 34008
rect 19432 33992 19484 33998
rect 19432 33934 19484 33940
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 18972 33652 19024 33658
rect 18972 33594 19024 33600
rect 18984 32978 19012 33594
rect 19340 33312 19392 33318
rect 19340 33254 19392 33260
rect 18972 32972 19024 32978
rect 18972 32914 19024 32920
rect 18984 32502 19012 32914
rect 19248 32768 19300 32774
rect 19248 32710 19300 32716
rect 19260 32502 19288 32710
rect 18972 32496 19024 32502
rect 18972 32438 19024 32444
rect 19248 32496 19300 32502
rect 19248 32438 19300 32444
rect 19352 31822 19380 33254
rect 20272 32994 20300 40582
rect 20444 39432 20496 39438
rect 20444 39374 20496 39380
rect 20456 39098 20484 39374
rect 20640 39098 20668 41414
rect 20732 41138 20760 42162
rect 21008 41614 21036 44678
rect 21100 44538 21128 45222
rect 21088 44532 21140 44538
rect 21088 44474 21140 44480
rect 21100 43722 21128 44474
rect 21192 44266 21220 45358
rect 21376 44402 21404 45494
rect 21456 45484 21508 45490
rect 21456 45426 21508 45432
rect 21468 44470 21496 45426
rect 21456 44464 21508 44470
rect 21456 44406 21508 44412
rect 21364 44396 21416 44402
rect 21364 44338 21416 44344
rect 21180 44260 21232 44266
rect 21180 44202 21232 44208
rect 21192 43790 21220 44202
rect 21180 43784 21232 43790
rect 21180 43726 21232 43732
rect 21088 43716 21140 43722
rect 21088 43658 21140 43664
rect 21376 43654 21404 44338
rect 21468 43790 21496 44406
rect 21456 43784 21508 43790
rect 21456 43726 21508 43732
rect 21364 43648 21416 43654
rect 21364 43590 21416 43596
rect 21088 43104 21140 43110
rect 21088 43046 21140 43052
rect 20996 41608 21048 41614
rect 20996 41550 21048 41556
rect 20720 41132 20772 41138
rect 20720 41074 20772 41080
rect 20732 40526 20760 41074
rect 20904 40996 20956 41002
rect 20904 40938 20956 40944
rect 20916 40526 20944 40938
rect 20720 40520 20772 40526
rect 20720 40462 20772 40468
rect 20904 40520 20956 40526
rect 20904 40462 20956 40468
rect 20732 40186 20760 40462
rect 20812 40452 20864 40458
rect 20812 40394 20864 40400
rect 20720 40180 20772 40186
rect 20720 40122 20772 40128
rect 20824 40050 20852 40394
rect 20812 40044 20864 40050
rect 20812 39986 20864 39992
rect 20824 39370 20852 39986
rect 20812 39364 20864 39370
rect 20812 39306 20864 39312
rect 20720 39296 20772 39302
rect 20720 39238 20772 39244
rect 20444 39092 20496 39098
rect 20444 39034 20496 39040
rect 20628 39092 20680 39098
rect 20628 39034 20680 39040
rect 20640 35834 20668 39034
rect 20732 39030 20760 39238
rect 20720 39024 20772 39030
rect 20720 38966 20772 38972
rect 20732 38214 20760 38966
rect 20824 38962 20852 39306
rect 21100 38962 21128 43046
rect 21376 42090 21404 43590
rect 21364 42084 21416 42090
rect 21364 42026 21416 42032
rect 21180 41608 21232 41614
rect 21180 41550 21232 41556
rect 21192 41070 21220 41550
rect 21272 41132 21324 41138
rect 21272 41074 21324 41080
rect 21180 41064 21232 41070
rect 21180 41006 21232 41012
rect 21284 40050 21312 41074
rect 21272 40044 21324 40050
rect 21272 39986 21324 39992
rect 21180 39840 21232 39846
rect 21180 39782 21232 39788
rect 21192 39642 21220 39782
rect 21180 39636 21232 39642
rect 21180 39578 21232 39584
rect 20812 38956 20864 38962
rect 20812 38898 20864 38904
rect 21088 38956 21140 38962
rect 21088 38898 21140 38904
rect 20996 38888 21048 38894
rect 20996 38830 21048 38836
rect 21272 38888 21324 38894
rect 21272 38830 21324 38836
rect 21008 38758 21036 38830
rect 20996 38752 21048 38758
rect 20996 38694 21048 38700
rect 21284 38418 21312 38830
rect 21468 38758 21496 43726
rect 21456 38752 21508 38758
rect 21456 38694 21508 38700
rect 21272 38412 21324 38418
rect 21272 38354 21324 38360
rect 20904 38344 20956 38350
rect 20904 38286 20956 38292
rect 21180 38344 21232 38350
rect 21180 38286 21232 38292
rect 20720 38208 20772 38214
rect 20720 38150 20772 38156
rect 20732 37890 20760 38150
rect 20916 37942 20944 38286
rect 21088 38276 21140 38282
rect 21088 38218 21140 38224
rect 20996 38208 21048 38214
rect 20996 38150 21048 38156
rect 20904 37936 20956 37942
rect 20732 37862 20852 37890
rect 20904 37878 20956 37884
rect 20720 37800 20772 37806
rect 20720 37742 20772 37748
rect 20628 35828 20680 35834
rect 20628 35770 20680 35776
rect 20628 35692 20680 35698
rect 20628 35634 20680 35640
rect 20640 35290 20668 35634
rect 20628 35284 20680 35290
rect 20628 35226 20680 35232
rect 20732 35154 20760 37742
rect 20824 37466 20852 37862
rect 21008 37754 21036 38150
rect 21100 37874 21128 38218
rect 21192 38010 21220 38286
rect 21180 38004 21232 38010
rect 21180 37946 21232 37952
rect 21088 37868 21140 37874
rect 21088 37810 21140 37816
rect 21284 37806 21312 38354
rect 21364 38208 21416 38214
rect 21364 38150 21416 38156
rect 21376 37942 21404 38150
rect 21364 37936 21416 37942
rect 21364 37878 21416 37884
rect 21272 37800 21324 37806
rect 20916 37738 21128 37754
rect 21272 37742 21324 37748
rect 20916 37732 21140 37738
rect 20916 37726 21088 37732
rect 20812 37460 20864 37466
rect 20812 37402 20864 37408
rect 20916 37262 20944 37726
rect 21088 37674 21140 37680
rect 21456 37664 21508 37670
rect 21456 37606 21508 37612
rect 20904 37256 20956 37262
rect 20904 37198 20956 37204
rect 20996 37120 21048 37126
rect 20996 37062 21048 37068
rect 20904 36032 20956 36038
rect 20904 35974 20956 35980
rect 20812 35692 20864 35698
rect 20812 35634 20864 35640
rect 20720 35148 20772 35154
rect 20720 35090 20772 35096
rect 20628 35080 20680 35086
rect 20628 35022 20680 35028
rect 20640 34610 20668 35022
rect 20628 34604 20680 34610
rect 20628 34546 20680 34552
rect 20824 34202 20852 35634
rect 20916 35630 20944 35974
rect 21008 35816 21036 37062
rect 21364 36780 21416 36786
rect 21364 36722 21416 36728
rect 21088 36644 21140 36650
rect 21088 36586 21140 36592
rect 21100 36378 21128 36586
rect 21088 36372 21140 36378
rect 21088 36314 21140 36320
rect 21100 35894 21128 36314
rect 21376 36106 21404 36722
rect 21468 36174 21496 37606
rect 21456 36168 21508 36174
rect 21456 36110 21508 36116
rect 21364 36100 21416 36106
rect 21364 36042 21416 36048
rect 21272 36032 21324 36038
rect 21272 35974 21324 35980
rect 21100 35866 21220 35894
rect 21008 35788 21128 35816
rect 20904 35624 20956 35630
rect 20904 35566 20956 35572
rect 21100 35562 21128 35788
rect 21088 35556 21140 35562
rect 21088 35498 21140 35504
rect 21192 35494 21220 35866
rect 20904 35488 20956 35494
rect 20904 35430 20956 35436
rect 21180 35488 21232 35494
rect 21180 35430 21232 35436
rect 20916 35290 20944 35430
rect 21284 35290 21312 35974
rect 20904 35284 20956 35290
rect 20904 35226 20956 35232
rect 21088 35284 21140 35290
rect 21088 35226 21140 35232
rect 21272 35284 21324 35290
rect 21272 35226 21324 35232
rect 21100 34610 21128 35226
rect 21376 35034 21404 36042
rect 21468 35630 21496 36110
rect 21456 35624 21508 35630
rect 21456 35566 21508 35572
rect 21284 35018 21404 35034
rect 21272 35012 21404 35018
rect 21324 35006 21404 35012
rect 21272 34954 21324 34960
rect 21088 34604 21140 34610
rect 21088 34546 21140 34552
rect 21284 34542 21312 34954
rect 21272 34536 21324 34542
rect 21272 34478 21324 34484
rect 20812 34196 20864 34202
rect 20812 34138 20864 34144
rect 21456 33856 21508 33862
rect 21456 33798 21508 33804
rect 21272 33448 21324 33454
rect 21272 33390 21324 33396
rect 20812 33312 20864 33318
rect 20812 33254 20864 33260
rect 20824 33130 20852 33254
rect 20180 32966 20300 32994
rect 20548 33102 20852 33130
rect 20076 32904 20128 32910
rect 20076 32846 20128 32852
rect 19432 32768 19484 32774
rect 19432 32710 19484 32716
rect 19444 32450 19472 32710
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19444 32434 19564 32450
rect 19444 32428 19576 32434
rect 19444 32422 19524 32428
rect 19524 32370 19576 32376
rect 20088 32298 20116 32846
rect 20076 32292 20128 32298
rect 20076 32234 20128 32240
rect 19340 31816 19392 31822
rect 19340 31758 19392 31764
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19524 31340 19576 31346
rect 19524 31282 19576 31288
rect 18880 31136 18932 31142
rect 18880 31078 18932 31084
rect 18892 28762 18920 31078
rect 19536 30666 19564 31282
rect 19616 31272 19668 31278
rect 19616 31214 19668 31220
rect 19628 30870 19656 31214
rect 19616 30864 19668 30870
rect 19616 30806 19668 30812
rect 19524 30660 19576 30666
rect 19444 30620 19524 30648
rect 19444 30326 19472 30620
rect 19524 30602 19576 30608
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19432 30320 19484 30326
rect 19432 30262 19484 30268
rect 19248 29640 19300 29646
rect 19248 29582 19300 29588
rect 19984 29640 20036 29646
rect 19984 29582 20036 29588
rect 19260 29306 19288 29582
rect 19340 29504 19392 29510
rect 19340 29446 19392 29452
rect 19248 29300 19300 29306
rect 19248 29242 19300 29248
rect 18880 28756 18932 28762
rect 18880 28698 18932 28704
rect 18788 28688 18840 28694
rect 18788 28630 18840 28636
rect 18892 27674 18920 28698
rect 19352 28626 19380 29446
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19800 28960 19852 28966
rect 19800 28902 19852 28908
rect 19432 28756 19484 28762
rect 19432 28698 19484 28704
rect 19444 28642 19472 28698
rect 19340 28620 19392 28626
rect 19444 28614 19656 28642
rect 19340 28562 19392 28568
rect 19352 28506 19380 28562
rect 19628 28558 19656 28614
rect 19812 28558 19840 28902
rect 19996 28694 20024 29582
rect 20180 29578 20208 32966
rect 20260 32904 20312 32910
rect 20260 32846 20312 32852
rect 20272 32570 20300 32846
rect 20260 32564 20312 32570
rect 20260 32506 20312 32512
rect 20272 31822 20300 32506
rect 20260 31816 20312 31822
rect 20260 31758 20312 31764
rect 20272 30734 20300 31758
rect 20548 31754 20576 33102
rect 20720 32768 20772 32774
rect 20720 32710 20772 32716
rect 20732 32366 20760 32710
rect 20812 32428 20864 32434
rect 20812 32370 20864 32376
rect 20720 32360 20772 32366
rect 20720 32302 20772 32308
rect 20732 31822 20760 32302
rect 20720 31816 20772 31822
rect 20720 31758 20772 31764
rect 20824 31754 20852 32370
rect 20996 31816 21048 31822
rect 20996 31758 21048 31764
rect 20536 31748 20588 31754
rect 20536 31690 20588 31696
rect 20812 31748 20864 31754
rect 20812 31690 20864 31696
rect 20444 31680 20496 31686
rect 20444 31622 20496 31628
rect 20456 31278 20484 31622
rect 20720 31340 20772 31346
rect 20720 31282 20772 31288
rect 20444 31272 20496 31278
rect 20444 31214 20496 31220
rect 20260 30728 20312 30734
rect 20260 30670 20312 30676
rect 20732 30258 20760 31282
rect 20824 30682 20852 31690
rect 20824 30654 20944 30682
rect 20812 30592 20864 30598
rect 20812 30534 20864 30540
rect 20720 30252 20772 30258
rect 20720 30194 20772 30200
rect 20260 30184 20312 30190
rect 20260 30126 20312 30132
rect 20168 29572 20220 29578
rect 20168 29514 20220 29520
rect 20168 29232 20220 29238
rect 20168 29174 20220 29180
rect 19984 28688 20036 28694
rect 19984 28630 20036 28636
rect 19616 28552 19668 28558
rect 19352 28478 19472 28506
rect 19616 28494 19668 28500
rect 19800 28552 19852 28558
rect 19800 28494 19852 28500
rect 19340 28416 19392 28422
rect 19340 28358 19392 28364
rect 18880 27668 18932 27674
rect 18880 27610 18932 27616
rect 19352 26450 19380 28358
rect 19444 27470 19472 28478
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19996 28218 20024 28630
rect 20076 28620 20128 28626
rect 20076 28562 20128 28568
rect 19984 28212 20036 28218
rect 19984 28154 20036 28160
rect 20088 27470 20116 28562
rect 20180 28082 20208 29174
rect 20272 29170 20300 30126
rect 20352 30048 20404 30054
rect 20352 29990 20404 29996
rect 20364 29782 20392 29990
rect 20352 29776 20404 29782
rect 20352 29718 20404 29724
rect 20260 29164 20312 29170
rect 20260 29106 20312 29112
rect 20168 28076 20220 28082
rect 20168 28018 20220 28024
rect 19432 27464 19484 27470
rect 19432 27406 19484 27412
rect 20076 27464 20128 27470
rect 20076 27406 20128 27412
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 20180 27130 20208 28018
rect 20272 28014 20300 29106
rect 20364 29034 20392 29718
rect 20824 29714 20852 30534
rect 20916 30326 20944 30654
rect 20904 30320 20956 30326
rect 20904 30262 20956 30268
rect 21008 30258 21036 31758
rect 21284 31754 21312 33390
rect 21364 33380 21416 33386
rect 21364 33322 21416 33328
rect 21376 32774 21404 33322
rect 21468 33318 21496 33798
rect 21456 33312 21508 33318
rect 21456 33254 21508 33260
rect 21468 32910 21496 33254
rect 21456 32904 21508 32910
rect 21456 32846 21508 32852
rect 21364 32768 21416 32774
rect 21364 32710 21416 32716
rect 21376 31890 21404 32710
rect 21364 31884 21416 31890
rect 21364 31826 21416 31832
rect 21272 31748 21324 31754
rect 21272 31690 21324 31696
rect 21284 30666 21312 31690
rect 21376 30734 21404 31826
rect 21364 30728 21416 30734
rect 21364 30670 21416 30676
rect 21272 30660 21324 30666
rect 21272 30602 21324 30608
rect 21456 30320 21508 30326
rect 21456 30262 21508 30268
rect 20996 30252 21048 30258
rect 20996 30194 21048 30200
rect 20904 29776 20956 29782
rect 20904 29718 20956 29724
rect 20812 29708 20864 29714
rect 20812 29650 20864 29656
rect 20812 29300 20864 29306
rect 20812 29242 20864 29248
rect 20352 29028 20404 29034
rect 20352 28970 20404 28976
rect 20720 29028 20772 29034
rect 20720 28970 20772 28976
rect 20364 28150 20392 28970
rect 20732 28150 20760 28970
rect 20824 28422 20852 29242
rect 20916 29170 20944 29718
rect 21272 29708 21324 29714
rect 21272 29650 21324 29656
rect 20904 29164 20956 29170
rect 20904 29106 20956 29112
rect 20904 28960 20956 28966
rect 20904 28902 20956 28908
rect 20916 28558 20944 28902
rect 21284 28762 21312 29650
rect 21468 29646 21496 30262
rect 21456 29640 21508 29646
rect 21456 29582 21508 29588
rect 21272 28756 21324 28762
rect 21272 28698 21324 28704
rect 20904 28552 20956 28558
rect 20904 28494 20956 28500
rect 21272 28552 21324 28558
rect 21272 28494 21324 28500
rect 20812 28416 20864 28422
rect 20812 28358 20864 28364
rect 20352 28144 20404 28150
rect 20352 28086 20404 28092
rect 20720 28144 20772 28150
rect 20720 28086 20772 28092
rect 20260 28008 20312 28014
rect 20260 27950 20312 27956
rect 20168 27124 20220 27130
rect 20168 27066 20220 27072
rect 20272 27062 20300 27950
rect 20732 27606 20760 28086
rect 20824 27878 20852 28358
rect 21284 28234 21312 28494
rect 21284 28206 21404 28234
rect 20812 27872 20864 27878
rect 20812 27814 20864 27820
rect 21272 27872 21324 27878
rect 21272 27814 21324 27820
rect 20720 27600 20772 27606
rect 20720 27542 20772 27548
rect 21088 27464 21140 27470
rect 21088 27406 21140 27412
rect 20260 27056 20312 27062
rect 20260 26998 20312 27004
rect 20996 26988 21048 26994
rect 21100 26976 21128 27406
rect 21048 26948 21128 26976
rect 20996 26930 21048 26936
rect 19340 26444 19392 26450
rect 19340 26386 19392 26392
rect 20168 26444 20220 26450
rect 20168 26386 20220 26392
rect 20076 26376 20128 26382
rect 20076 26318 20128 26324
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 20088 26042 20116 26318
rect 20076 26036 20128 26042
rect 20076 25978 20128 25984
rect 19340 25968 19392 25974
rect 20180 25922 20208 26386
rect 21100 26246 21128 26948
rect 21284 26926 21312 27814
rect 21376 27674 21404 28206
rect 21456 28008 21508 28014
rect 21456 27950 21508 27956
rect 21364 27668 21416 27674
rect 21364 27610 21416 27616
rect 21468 27538 21496 27950
rect 21456 27532 21508 27538
rect 21456 27474 21508 27480
rect 21468 26994 21496 27474
rect 21456 26988 21508 26994
rect 21456 26930 21508 26936
rect 21272 26920 21324 26926
rect 21272 26862 21324 26868
rect 21468 26518 21496 26930
rect 21456 26512 21508 26518
rect 21456 26454 21508 26460
rect 21088 26240 21140 26246
rect 21088 26182 21140 26188
rect 19340 25910 19392 25916
rect 19352 25702 19380 25910
rect 19984 25900 20036 25906
rect 19984 25842 20036 25848
rect 20088 25894 20208 25922
rect 19340 25696 19392 25702
rect 19340 25638 19392 25644
rect 19352 24614 19380 25638
rect 19996 25294 20024 25842
rect 20088 25430 20116 25894
rect 21100 25702 21128 26182
rect 20168 25696 20220 25702
rect 20168 25638 20220 25644
rect 21088 25696 21140 25702
rect 21088 25638 21140 25644
rect 20076 25424 20128 25430
rect 20076 25366 20128 25372
rect 20180 25362 20208 25638
rect 20168 25356 20220 25362
rect 20168 25298 20220 25304
rect 20904 25356 20956 25362
rect 20904 25298 20956 25304
rect 19984 25288 20036 25294
rect 19984 25230 20036 25236
rect 20812 25288 20864 25294
rect 20812 25230 20864 25236
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19996 24954 20024 25230
rect 20824 24954 20852 25230
rect 19984 24948 20036 24954
rect 19984 24890 20036 24896
rect 20812 24948 20864 24954
rect 20812 24890 20864 24896
rect 20720 24880 20772 24886
rect 20720 24822 20772 24828
rect 19340 24608 19392 24614
rect 19340 24550 19392 24556
rect 19352 16574 19380 24550
rect 20732 24410 20760 24822
rect 20916 24818 20944 25298
rect 20904 24812 20956 24818
rect 20904 24754 20956 24760
rect 20720 24404 20772 24410
rect 20720 24346 20772 24352
rect 20536 24132 20588 24138
rect 20536 24074 20588 24080
rect 20812 24132 20864 24138
rect 20812 24074 20864 24080
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 20548 23730 20576 24074
rect 20824 23730 20852 24074
rect 20536 23724 20588 23730
rect 20536 23666 20588 23672
rect 20812 23724 20864 23730
rect 20812 23666 20864 23672
rect 19984 23520 20036 23526
rect 19984 23462 20036 23468
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19352 16546 19472 16574
rect 17960 7200 18012 7206
rect 17960 7142 18012 7148
rect 19340 2848 19392 2854
rect 19340 2790 19392 2796
rect 16856 2508 16908 2514
rect 16856 2450 16908 2456
rect 19352 2446 19380 2790
rect 19444 2582 19472 16546
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19432 2576 19484 2582
rect 19432 2518 19484 2524
rect 19996 2514 20024 23462
rect 20824 23322 20852 23666
rect 20812 23316 20864 23322
rect 20812 23258 20864 23264
rect 21100 13938 21128 25638
rect 21272 24812 21324 24818
rect 21272 24754 21324 24760
rect 21284 23866 21312 24754
rect 21364 24744 21416 24750
rect 21364 24686 21416 24692
rect 21376 24410 21404 24686
rect 21364 24404 21416 24410
rect 21364 24346 21416 24352
rect 21272 23860 21324 23866
rect 21272 23802 21324 23808
rect 21088 13932 21140 13938
rect 21088 13874 21140 13880
rect 21272 2848 21324 2854
rect 21272 2790 21324 2796
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 16304 2372 16356 2378
rect 16304 2314 16356 2320
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 16776 800 16804 2246
rect 17696 1970 17724 2246
rect 17684 1964 17736 1970
rect 17684 1906 17736 1912
rect 19352 800 19380 2382
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 21284 800 21312 2790
rect 21560 2650 21588 47398
rect 21824 46912 21876 46918
rect 21824 46854 21876 46860
rect 21836 46510 21864 46854
rect 22100 46708 22152 46714
rect 22100 46650 22152 46656
rect 21824 46504 21876 46510
rect 21824 46446 21876 46452
rect 21824 45892 21876 45898
rect 21824 45834 21876 45840
rect 21640 45348 21692 45354
rect 21640 45290 21692 45296
rect 21652 44878 21680 45290
rect 21640 44872 21692 44878
rect 21640 44814 21692 44820
rect 21836 44470 21864 45834
rect 22112 45540 22140 46650
rect 22020 45512 22140 45540
rect 22020 45370 22048 45512
rect 22112 45422 22140 45453
rect 22100 45416 22152 45422
rect 22020 45364 22100 45370
rect 22020 45358 22152 45364
rect 22020 45342 22140 45358
rect 22112 45286 22140 45342
rect 22100 45280 22152 45286
rect 22100 45222 22152 45228
rect 22008 44872 22060 44878
rect 22008 44814 22060 44820
rect 21824 44464 21876 44470
rect 21824 44406 21876 44412
rect 21836 43874 21864 44406
rect 21836 43846 21956 43874
rect 21824 42288 21876 42294
rect 21824 42230 21876 42236
rect 21640 41744 21692 41750
rect 21638 41712 21640 41721
rect 21692 41712 21694 41721
rect 21638 41647 21694 41656
rect 21836 41614 21864 42230
rect 21824 41608 21876 41614
rect 21824 41550 21876 41556
rect 21928 40390 21956 43846
rect 22020 43790 22048 44814
rect 22100 44328 22152 44334
rect 22100 44270 22152 44276
rect 22112 43790 22140 44270
rect 22008 43784 22060 43790
rect 22008 43726 22060 43732
rect 22100 43784 22152 43790
rect 22100 43726 22152 43732
rect 22100 43308 22152 43314
rect 22100 43250 22152 43256
rect 22112 42770 22140 43250
rect 22008 42764 22060 42770
rect 22008 42706 22060 42712
rect 22100 42764 22152 42770
rect 22100 42706 22152 42712
rect 22020 42022 22048 42706
rect 22008 42016 22060 42022
rect 22008 41958 22060 41964
rect 21916 40384 21968 40390
rect 21916 40326 21968 40332
rect 21824 38956 21876 38962
rect 21824 38898 21876 38904
rect 21640 38344 21692 38350
rect 21640 38286 21692 38292
rect 21652 36922 21680 38286
rect 21836 38214 21864 38898
rect 21928 38729 21956 40326
rect 22204 39642 22232 51046
rect 22572 50930 22600 51274
rect 22560 50924 22612 50930
rect 22560 50866 22612 50872
rect 22572 50522 22600 50866
rect 22560 50516 22612 50522
rect 22560 50458 22612 50464
rect 22664 50318 22692 51546
rect 23584 51542 23612 51954
rect 23572 51536 23624 51542
rect 23572 51478 23624 51484
rect 23676 51338 23704 51954
rect 23768 51406 23796 52022
rect 23860 52018 23888 52294
rect 23848 52012 23900 52018
rect 23848 51954 23900 51960
rect 23848 51536 23900 51542
rect 23848 51478 23900 51484
rect 23756 51400 23808 51406
rect 23756 51342 23808 51348
rect 23664 51332 23716 51338
rect 23664 51274 23716 51280
rect 23676 51074 23704 51274
rect 23584 51046 23704 51074
rect 22744 50924 22796 50930
rect 22744 50866 22796 50872
rect 23204 50924 23256 50930
rect 23204 50866 23256 50872
rect 22652 50312 22704 50318
rect 22652 50254 22704 50260
rect 22664 49842 22692 50254
rect 22756 49978 22784 50866
rect 23216 50318 23244 50866
rect 23480 50720 23532 50726
rect 23480 50662 23532 50668
rect 23492 50454 23520 50662
rect 23480 50448 23532 50454
rect 23480 50390 23532 50396
rect 23204 50312 23256 50318
rect 23204 50254 23256 50260
rect 23584 50250 23612 51046
rect 23768 50726 23796 51342
rect 23860 51066 23888 51478
rect 24044 51074 24072 52566
rect 24504 52494 24532 53178
rect 25596 52556 25648 52562
rect 25596 52498 25648 52504
rect 24492 52488 24544 52494
rect 24492 52430 24544 52436
rect 24504 51474 24532 52430
rect 25608 52154 25636 52498
rect 25596 52148 25648 52154
rect 25596 52090 25648 52096
rect 24860 51536 24912 51542
rect 24860 51478 24912 51484
rect 24492 51468 24544 51474
rect 24492 51410 24544 51416
rect 23848 51060 23900 51066
rect 23848 51002 23900 51008
rect 23952 51046 24072 51074
rect 23952 50930 23980 51046
rect 24504 50998 24532 51410
rect 24872 51074 24900 51478
rect 24952 51400 25004 51406
rect 24952 51342 25004 51348
rect 25596 51400 25648 51406
rect 25596 51342 25648 51348
rect 24780 51046 24900 51074
rect 24492 50992 24544 50998
rect 24492 50934 24544 50940
rect 23940 50924 23992 50930
rect 23940 50866 23992 50872
rect 23756 50720 23808 50726
rect 23756 50662 23808 50668
rect 23572 50244 23624 50250
rect 23572 50186 23624 50192
rect 22744 49972 22796 49978
rect 22744 49914 22796 49920
rect 22652 49836 22704 49842
rect 22652 49778 22704 49784
rect 23480 49632 23532 49638
rect 23480 49574 23532 49580
rect 23492 49230 23520 49574
rect 23480 49224 23532 49230
rect 23480 49166 23532 49172
rect 23584 48890 23612 50186
rect 23848 49700 23900 49706
rect 23848 49642 23900 49648
rect 23664 49292 23716 49298
rect 23664 49234 23716 49240
rect 23572 48884 23624 48890
rect 23572 48826 23624 48832
rect 23676 48686 23704 49234
rect 23756 49156 23808 49162
rect 23756 49098 23808 49104
rect 23664 48680 23716 48686
rect 23664 48622 23716 48628
rect 22928 48612 22980 48618
rect 22928 48554 22980 48560
rect 23572 48612 23624 48618
rect 23572 48554 23624 48560
rect 22940 48142 22968 48554
rect 23584 48521 23612 48554
rect 23570 48512 23626 48521
rect 23570 48447 23626 48456
rect 22928 48136 22980 48142
rect 22928 48078 22980 48084
rect 23112 48000 23164 48006
rect 23112 47942 23164 47948
rect 22284 47660 22336 47666
rect 22284 47602 22336 47608
rect 22296 47530 22324 47602
rect 22284 47524 22336 47530
rect 22284 47466 22336 47472
rect 22468 46980 22520 46986
rect 22468 46922 22520 46928
rect 22376 46912 22428 46918
rect 22376 46854 22428 46860
rect 22388 46714 22416 46854
rect 22376 46708 22428 46714
rect 22376 46650 22428 46656
rect 22284 46504 22336 46510
rect 22284 46446 22336 46452
rect 22296 44402 22324 46446
rect 22376 46368 22428 46374
rect 22376 46310 22428 46316
rect 22388 45626 22416 46310
rect 22376 45620 22428 45626
rect 22376 45562 22428 45568
rect 22376 45416 22428 45422
rect 22376 45358 22428 45364
rect 22284 44396 22336 44402
rect 22284 44338 22336 44344
rect 22296 43858 22324 44338
rect 22284 43852 22336 43858
rect 22284 43794 22336 43800
rect 22388 43314 22416 45358
rect 22480 44878 22508 46922
rect 22836 45960 22888 45966
rect 22836 45902 22888 45908
rect 22744 45484 22796 45490
rect 22744 45426 22796 45432
rect 22560 45348 22612 45354
rect 22560 45290 22612 45296
rect 22572 45082 22600 45290
rect 22756 45082 22784 45426
rect 22560 45076 22612 45082
rect 22560 45018 22612 45024
rect 22744 45076 22796 45082
rect 22744 45018 22796 45024
rect 22468 44872 22520 44878
rect 22468 44814 22520 44820
rect 22480 44334 22508 44814
rect 22848 44402 22876 45902
rect 23020 45824 23072 45830
rect 23020 45766 23072 45772
rect 22928 45008 22980 45014
rect 22928 44950 22980 44956
rect 22940 44810 22968 44950
rect 22928 44804 22980 44810
rect 22928 44746 22980 44752
rect 23032 44742 23060 45766
rect 23124 45082 23152 47942
rect 23388 47592 23440 47598
rect 23388 47534 23440 47540
rect 23400 47122 23428 47534
rect 23676 47530 23704 48622
rect 23664 47524 23716 47530
rect 23664 47466 23716 47472
rect 23388 47116 23440 47122
rect 23388 47058 23440 47064
rect 23400 46578 23428 47058
rect 23572 47048 23624 47054
rect 23572 46990 23624 46996
rect 23584 46578 23612 46990
rect 23768 46714 23796 49098
rect 23860 48754 23888 49642
rect 23952 49298 23980 50866
rect 24032 50720 24084 50726
rect 24032 50662 24084 50668
rect 24044 50182 24072 50662
rect 24032 50176 24084 50182
rect 24032 50118 24084 50124
rect 24676 50176 24728 50182
rect 24676 50118 24728 50124
rect 24044 49842 24072 50118
rect 24492 49972 24544 49978
rect 24492 49914 24544 49920
rect 24504 49842 24532 49914
rect 24032 49836 24084 49842
rect 24032 49778 24084 49784
rect 24308 49836 24360 49842
rect 24308 49778 24360 49784
rect 24492 49836 24544 49842
rect 24492 49778 24544 49784
rect 23940 49292 23992 49298
rect 23940 49234 23992 49240
rect 23848 48748 23900 48754
rect 23848 48690 23900 48696
rect 23860 48074 23888 48690
rect 23940 48680 23992 48686
rect 23940 48622 23992 48628
rect 23848 48068 23900 48074
rect 23848 48010 23900 48016
rect 23952 47802 23980 48622
rect 24044 48618 24072 49778
rect 24032 48612 24084 48618
rect 24032 48554 24084 48560
rect 24032 48272 24084 48278
rect 24032 48214 24084 48220
rect 24044 47802 24072 48214
rect 24320 48210 24348 49778
rect 24492 49632 24544 49638
rect 24492 49574 24544 49580
rect 24504 49230 24532 49574
rect 24400 49224 24452 49230
rect 24400 49166 24452 49172
rect 24492 49224 24544 49230
rect 24492 49166 24544 49172
rect 24308 48204 24360 48210
rect 24308 48146 24360 48152
rect 23940 47796 23992 47802
rect 23940 47738 23992 47744
rect 24032 47796 24084 47802
rect 24032 47738 24084 47744
rect 24412 47190 24440 49166
rect 24504 48822 24532 49166
rect 24492 48816 24544 48822
rect 24492 48758 24544 48764
rect 24400 47184 24452 47190
rect 24400 47126 24452 47132
rect 23756 46708 23808 46714
rect 23756 46650 23808 46656
rect 24412 46578 24440 47126
rect 23388 46572 23440 46578
rect 23388 46514 23440 46520
rect 23572 46572 23624 46578
rect 23572 46514 23624 46520
rect 24400 46572 24452 46578
rect 24400 46514 24452 46520
rect 24504 46510 24532 48758
rect 24688 47258 24716 50118
rect 24780 49910 24808 51046
rect 24964 50862 24992 51342
rect 25608 50930 25636 51342
rect 25136 50924 25188 50930
rect 25136 50866 25188 50872
rect 25596 50924 25648 50930
rect 25596 50866 25648 50872
rect 25872 50924 25924 50930
rect 25872 50866 25924 50872
rect 24952 50856 25004 50862
rect 24952 50798 25004 50804
rect 24964 50522 24992 50798
rect 24952 50516 25004 50522
rect 24952 50458 25004 50464
rect 24860 50244 24912 50250
rect 24860 50186 24912 50192
rect 24768 49904 24820 49910
rect 24768 49846 24820 49852
rect 24872 49842 24900 50186
rect 24860 49836 24912 49842
rect 24860 49778 24912 49784
rect 24872 49366 24900 49778
rect 24860 49360 24912 49366
rect 24860 49302 24912 49308
rect 25044 49156 25096 49162
rect 25044 49098 25096 49104
rect 24860 48748 24912 48754
rect 24860 48690 24912 48696
rect 24872 48346 24900 48690
rect 25056 48618 25084 49098
rect 25148 48822 25176 50866
rect 25780 50788 25832 50794
rect 25780 50730 25832 50736
rect 25792 50386 25820 50730
rect 25780 50380 25832 50386
rect 25780 50322 25832 50328
rect 25884 50318 25912 50866
rect 25872 50312 25924 50318
rect 25872 50254 25924 50260
rect 25504 50244 25556 50250
rect 25504 50186 25556 50192
rect 25516 49842 25544 50186
rect 25504 49836 25556 49842
rect 25504 49778 25556 49784
rect 25884 49774 25912 50254
rect 25872 49768 25924 49774
rect 25872 49710 25924 49716
rect 25412 49428 25464 49434
rect 25412 49370 25464 49376
rect 25320 49088 25372 49094
rect 25320 49030 25372 49036
rect 25136 48816 25188 48822
rect 25136 48758 25188 48764
rect 25044 48612 25096 48618
rect 25044 48554 25096 48560
rect 24860 48340 24912 48346
rect 24860 48282 24912 48288
rect 25056 48278 25084 48554
rect 25044 48272 25096 48278
rect 24964 48232 25044 48260
rect 24860 48136 24912 48142
rect 24860 48078 24912 48084
rect 24676 47252 24728 47258
rect 24676 47194 24728 47200
rect 24584 47116 24636 47122
rect 24584 47058 24636 47064
rect 24596 46900 24624 47058
rect 24688 47054 24716 47194
rect 24676 47048 24728 47054
rect 24676 46990 24728 46996
rect 24596 46872 24716 46900
rect 24492 46504 24544 46510
rect 24492 46446 24544 46452
rect 23204 46436 23256 46442
rect 23204 46378 23256 46384
rect 23216 46170 23244 46378
rect 23204 46164 23256 46170
rect 23204 46106 23256 46112
rect 23112 45076 23164 45082
rect 23112 45018 23164 45024
rect 23020 44736 23072 44742
rect 23020 44678 23072 44684
rect 22836 44396 22888 44402
rect 22836 44338 22888 44344
rect 22468 44328 22520 44334
rect 22468 44270 22520 44276
rect 22848 43790 22876 44338
rect 22836 43784 22888 43790
rect 22836 43726 22888 43732
rect 22376 43308 22428 43314
rect 22376 43250 22428 43256
rect 22376 43172 22428 43178
rect 22376 43114 22428 43120
rect 22388 42362 22416 43114
rect 22376 42356 22428 42362
rect 22376 42298 22428 42304
rect 22744 41608 22796 41614
rect 22744 41550 22796 41556
rect 22756 41002 22784 41550
rect 23032 41414 23060 44678
rect 23216 43450 23244 46106
rect 24400 45892 24452 45898
rect 24400 45834 24452 45840
rect 24412 45626 24440 45834
rect 24492 45824 24544 45830
rect 24492 45766 24544 45772
rect 24400 45620 24452 45626
rect 24400 45562 24452 45568
rect 23756 45484 23808 45490
rect 23756 45426 23808 45432
rect 23388 45280 23440 45286
rect 23388 45222 23440 45228
rect 23400 44946 23428 45222
rect 23388 44940 23440 44946
rect 23388 44882 23440 44888
rect 23400 44538 23428 44882
rect 23768 44878 23796 45426
rect 23940 45416 23992 45422
rect 23940 45358 23992 45364
rect 23756 44872 23808 44878
rect 23756 44814 23808 44820
rect 23388 44532 23440 44538
rect 23388 44474 23440 44480
rect 23572 44464 23624 44470
rect 23572 44406 23624 44412
rect 23480 44396 23532 44402
rect 23480 44338 23532 44344
rect 23492 43722 23520 44338
rect 23584 43790 23612 44406
rect 23768 43994 23796 44814
rect 23848 44396 23900 44402
rect 23848 44338 23900 44344
rect 23756 43988 23808 43994
rect 23756 43930 23808 43936
rect 23572 43784 23624 43790
rect 23572 43726 23624 43732
rect 23860 43722 23888 44338
rect 23952 43926 23980 45358
rect 24412 45286 24440 45562
rect 24216 45280 24268 45286
rect 24216 45222 24268 45228
rect 24400 45280 24452 45286
rect 24400 45222 24452 45228
rect 24228 44334 24256 45222
rect 24412 44878 24440 45222
rect 24400 44872 24452 44878
rect 24400 44814 24452 44820
rect 24216 44328 24268 44334
rect 24216 44270 24268 44276
rect 23940 43920 23992 43926
rect 23940 43862 23992 43868
rect 23480 43716 23532 43722
rect 23480 43658 23532 43664
rect 23848 43716 23900 43722
rect 23848 43658 23900 43664
rect 23204 43444 23256 43450
rect 23204 43386 23256 43392
rect 23216 43330 23244 43386
rect 23124 43302 23244 43330
rect 23388 43308 23440 43314
rect 23124 42702 23152 43302
rect 23388 43250 23440 43256
rect 23204 43104 23256 43110
rect 23204 43046 23256 43052
rect 23112 42696 23164 42702
rect 23112 42638 23164 42644
rect 23124 42158 23152 42638
rect 23216 42226 23244 43046
rect 23296 42288 23348 42294
rect 23296 42230 23348 42236
rect 23204 42220 23256 42226
rect 23204 42162 23256 42168
rect 23112 42152 23164 42158
rect 23112 42094 23164 42100
rect 23308 41614 23336 42230
rect 23400 42226 23428 43250
rect 23492 42702 23520 43658
rect 23572 43648 23624 43654
rect 23572 43590 23624 43596
rect 23584 43314 23612 43590
rect 23860 43382 23888 43658
rect 23848 43376 23900 43382
rect 23848 43318 23900 43324
rect 23572 43308 23624 43314
rect 23572 43250 23624 43256
rect 23664 43172 23716 43178
rect 23664 43114 23716 43120
rect 23676 42770 23704 43114
rect 23664 42764 23716 42770
rect 23664 42706 23716 42712
rect 23480 42696 23532 42702
rect 23480 42638 23532 42644
rect 23860 42362 23888 43318
rect 23952 43314 23980 43862
rect 24032 43852 24084 43858
rect 24032 43794 24084 43800
rect 24044 43722 24072 43794
rect 24032 43716 24084 43722
rect 24032 43658 24084 43664
rect 23940 43308 23992 43314
rect 23940 43250 23992 43256
rect 24044 42838 24072 43658
rect 24400 43648 24452 43654
rect 24400 43590 24452 43596
rect 24308 43104 24360 43110
rect 24308 43046 24360 43052
rect 24032 42832 24084 42838
rect 24032 42774 24084 42780
rect 24216 42560 24268 42566
rect 24216 42502 24268 42508
rect 23848 42356 23900 42362
rect 23848 42298 23900 42304
rect 24228 42226 24256 42502
rect 23388 42220 23440 42226
rect 23388 42162 23440 42168
rect 24216 42220 24268 42226
rect 24216 42162 24268 42168
rect 23296 41608 23348 41614
rect 23296 41550 23348 41556
rect 23846 41576 23902 41585
rect 23846 41511 23848 41520
rect 23900 41511 23902 41520
rect 23848 41482 23900 41488
rect 23032 41386 23152 41414
rect 22744 40996 22796 41002
rect 22744 40938 22796 40944
rect 22468 40384 22520 40390
rect 22468 40326 22520 40332
rect 22376 40044 22428 40050
rect 22376 39986 22428 39992
rect 22388 39642 22416 39986
rect 22480 39642 22508 40326
rect 22192 39636 22244 39642
rect 22192 39578 22244 39584
rect 22376 39636 22428 39642
rect 22376 39578 22428 39584
rect 22468 39636 22520 39642
rect 22468 39578 22520 39584
rect 22204 38978 22232 39578
rect 22376 39432 22428 39438
rect 22376 39374 22428 39380
rect 22388 39098 22416 39374
rect 22756 39370 22784 40938
rect 23124 40934 23152 41386
rect 23860 41138 23888 41482
rect 23664 41132 23716 41138
rect 23664 41074 23716 41080
rect 23848 41132 23900 41138
rect 23848 41074 23900 41080
rect 24032 41132 24084 41138
rect 24032 41074 24084 41080
rect 23388 41064 23440 41070
rect 23388 41006 23440 41012
rect 23112 40928 23164 40934
rect 23112 40870 23164 40876
rect 22836 39976 22888 39982
rect 22836 39918 22888 39924
rect 22560 39364 22612 39370
rect 22560 39306 22612 39312
rect 22744 39364 22796 39370
rect 22744 39306 22796 39312
rect 22468 39296 22520 39302
rect 22468 39238 22520 39244
rect 22376 39092 22428 39098
rect 22376 39034 22428 39040
rect 22008 38956 22060 38962
rect 22204 38950 22324 38978
rect 22008 38898 22060 38904
rect 21914 38720 21970 38729
rect 21914 38655 21970 38664
rect 22020 38418 22048 38898
rect 22192 38888 22244 38894
rect 22192 38830 22244 38836
rect 22204 38758 22232 38830
rect 22192 38752 22244 38758
rect 22192 38694 22244 38700
rect 22008 38412 22060 38418
rect 22008 38354 22060 38360
rect 22204 38350 22232 38694
rect 22192 38344 22244 38350
rect 22192 38286 22244 38292
rect 21824 38208 21876 38214
rect 21824 38150 21876 38156
rect 22100 38208 22152 38214
rect 22100 38150 22152 38156
rect 21824 37800 21876 37806
rect 21824 37742 21876 37748
rect 21836 36922 21864 37742
rect 21640 36916 21692 36922
rect 21640 36858 21692 36864
rect 21824 36916 21876 36922
rect 21824 36858 21876 36864
rect 21732 36644 21784 36650
rect 21732 36586 21784 36592
rect 21640 36236 21692 36242
rect 21640 36178 21692 36184
rect 21652 35698 21680 36178
rect 21744 36174 21772 36586
rect 21916 36304 21968 36310
rect 21916 36246 21968 36252
rect 21732 36168 21784 36174
rect 21732 36110 21784 36116
rect 21640 35692 21692 35698
rect 21640 35634 21692 35640
rect 21824 35488 21876 35494
rect 21824 35430 21876 35436
rect 21836 30258 21864 35430
rect 21928 35154 21956 36246
rect 21916 35148 21968 35154
rect 21916 35090 21968 35096
rect 22008 34468 22060 34474
rect 22008 34410 22060 34416
rect 22020 33998 22048 34410
rect 22008 33992 22060 33998
rect 22008 33934 22060 33940
rect 21916 33584 21968 33590
rect 21916 33526 21968 33532
rect 21928 32842 21956 33526
rect 22008 32904 22060 32910
rect 22008 32846 22060 32852
rect 21916 32836 21968 32842
rect 21916 32778 21968 32784
rect 21928 32434 21956 32778
rect 22020 32502 22048 32846
rect 22008 32496 22060 32502
rect 22008 32438 22060 32444
rect 21916 32428 21968 32434
rect 21916 32370 21968 32376
rect 22008 31136 22060 31142
rect 22008 31078 22060 31084
rect 22020 30802 22048 31078
rect 22008 30796 22060 30802
rect 22008 30738 22060 30744
rect 22112 30258 22140 38150
rect 22296 37330 22324 38950
rect 22480 37806 22508 39238
rect 22572 38962 22600 39306
rect 22848 39098 22876 39918
rect 23124 39370 23152 40870
rect 23296 40588 23348 40594
rect 23296 40530 23348 40536
rect 23308 40050 23336 40530
rect 23400 40526 23428 41006
rect 23676 40662 23704 41074
rect 23756 40928 23808 40934
rect 23756 40870 23808 40876
rect 23664 40656 23716 40662
rect 23664 40598 23716 40604
rect 23676 40526 23704 40598
rect 23388 40520 23440 40526
rect 23388 40462 23440 40468
rect 23664 40520 23716 40526
rect 23664 40462 23716 40468
rect 23296 40044 23348 40050
rect 23296 39986 23348 39992
rect 23480 39840 23532 39846
rect 23480 39782 23532 39788
rect 23492 39506 23520 39782
rect 23664 39636 23716 39642
rect 23664 39578 23716 39584
rect 23480 39500 23532 39506
rect 23480 39442 23532 39448
rect 23676 39438 23704 39578
rect 23768 39438 23796 40870
rect 23940 40180 23992 40186
rect 23940 40122 23992 40128
rect 23952 40050 23980 40122
rect 23940 40044 23992 40050
rect 23940 39986 23992 39992
rect 23664 39432 23716 39438
rect 23664 39374 23716 39380
rect 23756 39432 23808 39438
rect 23756 39374 23808 39380
rect 23112 39364 23164 39370
rect 23112 39306 23164 39312
rect 22836 39092 22888 39098
rect 22836 39034 22888 39040
rect 22560 38956 22612 38962
rect 22560 38898 22612 38904
rect 22558 38720 22614 38729
rect 22558 38655 22614 38664
rect 22468 37800 22520 37806
rect 22468 37742 22520 37748
rect 22376 37392 22428 37398
rect 22376 37334 22428 37340
rect 22192 37324 22244 37330
rect 22192 37266 22244 37272
rect 22284 37324 22336 37330
rect 22284 37266 22336 37272
rect 22204 34626 22232 37266
rect 22296 36582 22324 37266
rect 22388 36854 22416 37334
rect 22480 37194 22508 37742
rect 22468 37188 22520 37194
rect 22468 37130 22520 37136
rect 22572 36922 22600 38655
rect 22836 38344 22888 38350
rect 22836 38286 22888 38292
rect 22848 37874 22876 38286
rect 22836 37868 22888 37874
rect 22836 37810 22888 37816
rect 22560 36916 22612 36922
rect 22560 36858 22612 36864
rect 22376 36848 22428 36854
rect 22376 36790 22428 36796
rect 22284 36576 22336 36582
rect 22284 36518 22336 36524
rect 22572 35680 22600 36858
rect 23020 36780 23072 36786
rect 23020 36722 23072 36728
rect 23032 36378 23060 36722
rect 23020 36372 23072 36378
rect 23020 36314 23072 36320
rect 22744 35692 22796 35698
rect 22572 35652 22744 35680
rect 22744 35634 22796 35640
rect 22756 35154 22784 35634
rect 22744 35148 22796 35154
rect 22744 35090 22796 35096
rect 22560 35080 22612 35086
rect 22560 35022 22612 35028
rect 22928 35080 22980 35086
rect 22928 35022 22980 35028
rect 22572 34746 22600 35022
rect 22940 34746 22968 35022
rect 22560 34740 22612 34746
rect 22560 34682 22612 34688
rect 22928 34740 22980 34746
rect 22928 34682 22980 34688
rect 22284 34672 22336 34678
rect 22204 34620 22284 34626
rect 23124 34626 23152 39306
rect 23296 39296 23348 39302
rect 23296 39238 23348 39244
rect 23308 38962 23336 39238
rect 23296 38956 23348 38962
rect 23296 38898 23348 38904
rect 23676 38654 23704 39374
rect 23768 39098 23796 39374
rect 23756 39092 23808 39098
rect 23756 39034 23808 39040
rect 23952 38962 23980 39986
rect 24044 39794 24072 41074
rect 24320 41070 24348 43046
rect 24412 41585 24440 43590
rect 24504 42702 24532 45766
rect 24688 45014 24716 46872
rect 24872 46714 24900 48078
rect 24964 47054 24992 48232
rect 25044 48214 25096 48220
rect 25148 47666 25176 48758
rect 25136 47660 25188 47666
rect 25136 47602 25188 47608
rect 24952 47048 25004 47054
rect 24952 46990 25004 46996
rect 25044 47048 25096 47054
rect 25044 46990 25096 46996
rect 24860 46708 24912 46714
rect 24860 46650 24912 46656
rect 25056 46170 25084 46990
rect 25044 46164 25096 46170
rect 25044 46106 25096 46112
rect 25148 45966 25176 47602
rect 25332 47598 25360 49030
rect 25424 48686 25452 49370
rect 25504 49224 25556 49230
rect 25504 49166 25556 49172
rect 25412 48680 25464 48686
rect 25412 48622 25464 48628
rect 25320 47592 25372 47598
rect 25320 47534 25372 47540
rect 25228 47184 25280 47190
rect 25228 47126 25280 47132
rect 25240 46714 25268 47126
rect 25228 46708 25280 46714
rect 25228 46650 25280 46656
rect 25424 46442 25452 48622
rect 25516 47734 25544 49166
rect 25688 47796 25740 47802
rect 25688 47738 25740 47744
rect 25504 47728 25556 47734
rect 25504 47670 25556 47676
rect 25516 47190 25544 47670
rect 25504 47184 25556 47190
rect 25504 47126 25556 47132
rect 25516 46510 25544 47126
rect 25700 46578 25728 47738
rect 25872 47592 25924 47598
rect 25872 47534 25924 47540
rect 25780 47048 25832 47054
rect 25780 46990 25832 46996
rect 25688 46572 25740 46578
rect 25688 46514 25740 46520
rect 25504 46504 25556 46510
rect 25504 46446 25556 46452
rect 25412 46436 25464 46442
rect 25412 46378 25464 46384
rect 25136 45960 25188 45966
rect 25136 45902 25188 45908
rect 25148 45626 25176 45902
rect 25136 45620 25188 45626
rect 25136 45562 25188 45568
rect 25424 45286 25452 46378
rect 25792 45558 25820 46990
rect 25884 46578 25912 47534
rect 25872 46572 25924 46578
rect 25872 46514 25924 46520
rect 25780 45552 25832 45558
rect 25780 45494 25832 45500
rect 25412 45280 25464 45286
rect 25412 45222 25464 45228
rect 24676 45008 24728 45014
rect 24676 44950 24728 44956
rect 25320 45008 25372 45014
rect 25320 44950 25372 44956
rect 24688 44878 24716 44950
rect 24676 44872 24728 44878
rect 24676 44814 24728 44820
rect 24688 44742 24716 44814
rect 24676 44736 24728 44742
rect 24676 44678 24728 44684
rect 25044 44736 25096 44742
rect 25044 44678 25096 44684
rect 25056 44198 25084 44678
rect 25044 44192 25096 44198
rect 25044 44134 25096 44140
rect 24584 43988 24636 43994
rect 24584 43930 24636 43936
rect 24596 43246 24624 43930
rect 25056 43858 25084 44134
rect 25044 43852 25096 43858
rect 25044 43794 25096 43800
rect 25056 43246 25084 43794
rect 25332 43790 25360 44950
rect 25424 44810 25452 45222
rect 25688 44872 25740 44878
rect 25688 44814 25740 44820
rect 25412 44804 25464 44810
rect 25412 44746 25464 44752
rect 25424 44470 25452 44746
rect 25412 44464 25464 44470
rect 25412 44406 25464 44412
rect 25504 44396 25556 44402
rect 25504 44338 25556 44344
rect 25596 44396 25648 44402
rect 25596 44338 25648 44344
rect 25320 43784 25372 43790
rect 25320 43726 25372 43732
rect 25516 43314 25544 44338
rect 25608 43722 25636 44338
rect 25700 43994 25728 44814
rect 25688 43988 25740 43994
rect 25688 43930 25740 43936
rect 25596 43716 25648 43722
rect 25596 43658 25648 43664
rect 25700 43450 25728 43930
rect 25792 43790 25820 45494
rect 25780 43784 25832 43790
rect 25780 43726 25832 43732
rect 25688 43444 25740 43450
rect 25688 43386 25740 43392
rect 25320 43308 25372 43314
rect 25320 43250 25372 43256
rect 25504 43308 25556 43314
rect 25556 43268 25636 43296
rect 25504 43250 25556 43256
rect 24584 43240 24636 43246
rect 24584 43182 24636 43188
rect 25044 43240 25096 43246
rect 25044 43182 25096 43188
rect 25044 43104 25096 43110
rect 25044 43046 25096 43052
rect 24492 42696 24544 42702
rect 24492 42638 24544 42644
rect 24504 42226 24532 42638
rect 24492 42220 24544 42226
rect 24492 42162 24544 42168
rect 24504 41818 24532 42162
rect 24492 41812 24544 41818
rect 24492 41754 24544 41760
rect 24398 41576 24454 41585
rect 24398 41511 24454 41520
rect 24676 41540 24728 41546
rect 24676 41482 24728 41488
rect 24688 41138 24716 41482
rect 24676 41132 24728 41138
rect 24676 41074 24728 41080
rect 24308 41064 24360 41070
rect 24308 41006 24360 41012
rect 24124 40452 24176 40458
rect 24124 40394 24176 40400
rect 24136 39982 24164 40394
rect 24216 40384 24268 40390
rect 24216 40326 24268 40332
rect 24228 40050 24256 40326
rect 24216 40044 24268 40050
rect 24216 39986 24268 39992
rect 24124 39976 24176 39982
rect 24124 39918 24176 39924
rect 24228 39914 24256 39986
rect 24216 39908 24268 39914
rect 24216 39850 24268 39856
rect 24044 39766 24164 39794
rect 23940 38956 23992 38962
rect 23940 38898 23992 38904
rect 23676 38626 23796 38654
rect 23388 37868 23440 37874
rect 23388 37810 23440 37816
rect 23400 37330 23428 37810
rect 23664 37392 23716 37398
rect 23664 37334 23716 37340
rect 23388 37324 23440 37330
rect 23388 37266 23440 37272
rect 23676 36786 23704 37334
rect 23664 36780 23716 36786
rect 23664 36722 23716 36728
rect 23676 36106 23704 36722
rect 23768 36718 23796 38626
rect 24032 38276 24084 38282
rect 24032 38218 24084 38224
rect 24044 37670 24072 38218
rect 23848 37664 23900 37670
rect 23848 37606 23900 37612
rect 24032 37664 24084 37670
rect 24032 37606 24084 37612
rect 23860 36786 23888 37606
rect 23940 37460 23992 37466
rect 23940 37402 23992 37408
rect 23848 36780 23900 36786
rect 23848 36722 23900 36728
rect 23756 36712 23808 36718
rect 23756 36654 23808 36660
rect 23860 36106 23888 36722
rect 23952 36650 23980 37402
rect 24044 37330 24072 37606
rect 24032 37324 24084 37330
rect 24032 37266 24084 37272
rect 24032 36712 24084 36718
rect 24032 36654 24084 36660
rect 23940 36644 23992 36650
rect 23940 36586 23992 36592
rect 23664 36100 23716 36106
rect 23664 36042 23716 36048
rect 23848 36100 23900 36106
rect 23848 36042 23900 36048
rect 23388 35488 23440 35494
rect 23388 35430 23440 35436
rect 23572 35488 23624 35494
rect 23572 35430 23624 35436
rect 23400 35290 23428 35430
rect 23388 35284 23440 35290
rect 23388 35226 23440 35232
rect 22204 34614 22336 34620
rect 22204 34598 22324 34614
rect 22940 34598 23152 34626
rect 22204 34134 22232 34598
rect 22652 34400 22704 34406
rect 22652 34342 22704 34348
rect 22192 34128 22244 34134
rect 22192 34070 22244 34076
rect 22204 33998 22232 34070
rect 22664 33998 22692 34342
rect 22192 33992 22244 33998
rect 22192 33934 22244 33940
rect 22652 33992 22704 33998
rect 22652 33934 22704 33940
rect 22560 33516 22612 33522
rect 22560 33458 22612 33464
rect 22652 33516 22704 33522
rect 22652 33458 22704 33464
rect 22572 32910 22600 33458
rect 22560 32904 22612 32910
rect 22560 32846 22612 32852
rect 22572 32434 22600 32846
rect 22664 32774 22692 33458
rect 22652 32768 22704 32774
rect 22652 32710 22704 32716
rect 22560 32428 22612 32434
rect 22560 32370 22612 32376
rect 22652 32224 22704 32230
rect 22652 32166 22704 32172
rect 22664 31822 22692 32166
rect 22192 31816 22244 31822
rect 22192 31758 22244 31764
rect 22652 31816 22704 31822
rect 22652 31758 22704 31764
rect 22204 31278 22232 31758
rect 22560 31680 22612 31686
rect 22560 31622 22612 31628
rect 22572 31346 22600 31622
rect 22664 31414 22692 31758
rect 22652 31408 22704 31414
rect 22652 31350 22704 31356
rect 22560 31340 22612 31346
rect 22560 31282 22612 31288
rect 22192 31272 22244 31278
rect 22192 31214 22244 31220
rect 22204 30938 22232 31214
rect 22192 30932 22244 30938
rect 22192 30874 22244 30880
rect 21824 30252 21876 30258
rect 21824 30194 21876 30200
rect 22100 30252 22152 30258
rect 22100 30194 22152 30200
rect 21836 30138 21864 30194
rect 21744 30110 21864 30138
rect 21744 29170 21772 30110
rect 22008 30048 22060 30054
rect 22008 29990 22060 29996
rect 22020 29646 22048 29990
rect 22008 29640 22060 29646
rect 22008 29582 22060 29588
rect 21732 29164 21784 29170
rect 21732 29106 21784 29112
rect 22020 29034 22048 29582
rect 22112 29306 22140 30194
rect 22940 29850 22968 34598
rect 23584 34066 23612 35430
rect 23676 34678 23704 36042
rect 23860 35290 23888 36042
rect 24044 36038 24072 36654
rect 24032 36032 24084 36038
rect 24032 35974 24084 35980
rect 23848 35284 23900 35290
rect 23848 35226 23900 35232
rect 23860 35086 23888 35226
rect 23848 35080 23900 35086
rect 23848 35022 23900 35028
rect 23664 34672 23716 34678
rect 23664 34614 23716 34620
rect 23572 34060 23624 34066
rect 23572 34002 23624 34008
rect 23296 33992 23348 33998
rect 23296 33934 23348 33940
rect 23308 33522 23336 33934
rect 23296 33516 23348 33522
rect 23296 33458 23348 33464
rect 23388 33516 23440 33522
rect 23388 33458 23440 33464
rect 23112 33312 23164 33318
rect 23112 33254 23164 33260
rect 23124 32892 23152 33254
rect 23308 32978 23336 33458
rect 23296 32972 23348 32978
rect 23296 32914 23348 32920
rect 23204 32904 23256 32910
rect 23124 32864 23204 32892
rect 23020 32768 23072 32774
rect 23020 32710 23072 32716
rect 23032 32314 23060 32710
rect 23124 32434 23152 32864
rect 23204 32846 23256 32852
rect 23296 32768 23348 32774
rect 23296 32710 23348 32716
rect 23112 32428 23164 32434
rect 23112 32370 23164 32376
rect 23204 32428 23256 32434
rect 23204 32370 23256 32376
rect 23216 32314 23244 32370
rect 23032 32286 23244 32314
rect 23112 31748 23164 31754
rect 23112 31690 23164 31696
rect 23124 31498 23152 31690
rect 23216 31686 23244 32286
rect 23308 32230 23336 32710
rect 23400 32298 23428 33458
rect 23584 33318 23612 34002
rect 23756 33992 23808 33998
rect 23756 33934 23808 33940
rect 23768 33454 23796 33934
rect 23756 33448 23808 33454
rect 23756 33390 23808 33396
rect 23572 33312 23624 33318
rect 23572 33254 23624 33260
rect 23768 32502 23796 33390
rect 23848 33312 23900 33318
rect 23848 33254 23900 33260
rect 23756 32496 23808 32502
rect 23756 32438 23808 32444
rect 23664 32428 23716 32434
rect 23664 32370 23716 32376
rect 23388 32292 23440 32298
rect 23388 32234 23440 32240
rect 23296 32224 23348 32230
rect 23296 32166 23348 32172
rect 23572 31816 23624 31822
rect 23492 31776 23572 31804
rect 23204 31680 23256 31686
rect 23204 31622 23256 31628
rect 23124 31470 23244 31498
rect 23492 31482 23520 31776
rect 23572 31758 23624 31764
rect 23216 31346 23244 31470
rect 23480 31476 23532 31482
rect 23480 31418 23532 31424
rect 23204 31340 23256 31346
rect 23204 31282 23256 31288
rect 23216 30734 23244 31282
rect 23388 31272 23440 31278
rect 23388 31214 23440 31220
rect 23204 30728 23256 30734
rect 23204 30670 23256 30676
rect 23400 30394 23428 31214
rect 23676 30938 23704 32370
rect 23860 32230 23888 33254
rect 23940 32768 23992 32774
rect 23940 32710 23992 32716
rect 23756 32224 23808 32230
rect 23756 32166 23808 32172
rect 23848 32224 23900 32230
rect 23848 32166 23900 32172
rect 23768 31482 23796 32166
rect 23756 31476 23808 31482
rect 23756 31418 23808 31424
rect 23756 31340 23808 31346
rect 23756 31282 23808 31288
rect 23664 30932 23716 30938
rect 23664 30874 23716 30880
rect 23572 30728 23624 30734
rect 23572 30670 23624 30676
rect 23388 30388 23440 30394
rect 23388 30330 23440 30336
rect 23480 30320 23532 30326
rect 23480 30262 23532 30268
rect 23388 30252 23440 30258
rect 23388 30194 23440 30200
rect 22928 29844 22980 29850
rect 22928 29786 22980 29792
rect 23204 29844 23256 29850
rect 23204 29786 23256 29792
rect 23112 29640 23164 29646
rect 23112 29582 23164 29588
rect 22284 29572 22336 29578
rect 22284 29514 22336 29520
rect 22100 29300 22152 29306
rect 22100 29242 22152 29248
rect 22100 29164 22152 29170
rect 22100 29106 22152 29112
rect 22008 29028 22060 29034
rect 22008 28970 22060 28976
rect 22112 28558 22140 29106
rect 22296 28558 22324 29514
rect 22836 29504 22888 29510
rect 22836 29446 22888 29452
rect 22848 29170 22876 29446
rect 23124 29170 23152 29582
rect 23216 29578 23244 29786
rect 23296 29776 23348 29782
rect 23296 29718 23348 29724
rect 23204 29572 23256 29578
rect 23204 29514 23256 29520
rect 22836 29164 22888 29170
rect 22836 29106 22888 29112
rect 23112 29164 23164 29170
rect 23112 29106 23164 29112
rect 22376 28960 22428 28966
rect 22376 28902 22428 28908
rect 22560 28960 22612 28966
rect 22560 28902 22612 28908
rect 22100 28552 22152 28558
rect 22100 28494 22152 28500
rect 22284 28552 22336 28558
rect 22284 28494 22336 28500
rect 22008 28484 22060 28490
rect 22008 28426 22060 28432
rect 22020 28218 22048 28426
rect 22388 28218 22416 28902
rect 22008 28212 22060 28218
rect 22008 28154 22060 28160
rect 22376 28212 22428 28218
rect 22376 28154 22428 28160
rect 21916 28144 21968 28150
rect 21916 28086 21968 28092
rect 21928 27470 21956 28086
rect 22020 28082 22048 28154
rect 22008 28076 22060 28082
rect 22008 28018 22060 28024
rect 22388 27674 22416 28154
rect 22376 27668 22428 27674
rect 22376 27610 22428 27616
rect 22572 27470 22600 28902
rect 23112 28484 23164 28490
rect 23112 28426 23164 28432
rect 22652 28416 22704 28422
rect 22652 28358 22704 28364
rect 21916 27464 21968 27470
rect 21916 27406 21968 27412
rect 22560 27464 22612 27470
rect 22560 27406 22612 27412
rect 22192 27396 22244 27402
rect 22192 27338 22244 27344
rect 22204 26994 22232 27338
rect 22284 27328 22336 27334
rect 22284 27270 22336 27276
rect 22296 26994 22324 27270
rect 22572 26994 22600 27406
rect 22664 27402 22692 28358
rect 23124 28082 23152 28426
rect 23112 28076 23164 28082
rect 23216 28064 23244 29514
rect 23308 29102 23336 29718
rect 23400 29714 23428 30194
rect 23388 29708 23440 29714
rect 23388 29650 23440 29656
rect 23492 29306 23520 30262
rect 23584 30258 23612 30670
rect 23768 30666 23796 31282
rect 23756 30660 23808 30666
rect 23756 30602 23808 30608
rect 23768 30258 23796 30602
rect 23572 30252 23624 30258
rect 23572 30194 23624 30200
rect 23756 30252 23808 30258
rect 23756 30194 23808 30200
rect 23664 30184 23716 30190
rect 23664 30126 23716 30132
rect 23676 29730 23704 30126
rect 23768 29850 23796 30194
rect 23952 30190 23980 32710
rect 24044 31890 24072 35974
rect 24136 35698 24164 39766
rect 24320 39302 24348 41006
rect 25056 40934 25084 43046
rect 25332 42770 25360 43250
rect 25412 43240 25464 43246
rect 25412 43182 25464 43188
rect 25320 42764 25372 42770
rect 25320 42706 25372 42712
rect 25332 41614 25360 42706
rect 25424 42702 25452 43182
rect 25412 42696 25464 42702
rect 25412 42638 25464 42644
rect 25424 42362 25452 42638
rect 25412 42356 25464 42362
rect 25412 42298 25464 42304
rect 25608 41614 25636 43268
rect 25792 42362 25820 43726
rect 25780 42356 25832 42362
rect 25780 42298 25832 42304
rect 25320 41608 25372 41614
rect 25320 41550 25372 41556
rect 25504 41608 25556 41614
rect 25504 41550 25556 41556
rect 25596 41608 25648 41614
rect 25596 41550 25648 41556
rect 25332 41138 25360 41550
rect 25516 41274 25544 41550
rect 25976 41414 26004 53926
rect 26240 52896 26292 52902
rect 26240 52838 26292 52844
rect 26148 52556 26200 52562
rect 26068 52516 26148 52544
rect 26068 51066 26096 52516
rect 26148 52498 26200 52504
rect 26252 52426 26280 52838
rect 26240 52420 26292 52426
rect 26240 52362 26292 52368
rect 26252 51882 26280 52362
rect 26240 51876 26292 51882
rect 26240 51818 26292 51824
rect 26252 51610 26280 51818
rect 26240 51604 26292 51610
rect 26240 51546 26292 51552
rect 26148 51264 26200 51270
rect 26148 51206 26200 51212
rect 26056 51060 26108 51066
rect 26056 51002 26108 51008
rect 26160 50862 26188 51206
rect 26148 50856 26200 50862
rect 26148 50798 26200 50804
rect 26252 50726 26280 51546
rect 26988 51542 27016 53926
rect 27160 53508 27212 53514
rect 27160 53450 27212 53456
rect 26976 51536 27028 51542
rect 26976 51478 27028 51484
rect 26240 50720 26292 50726
rect 26240 50662 26292 50668
rect 26884 50720 26936 50726
rect 26884 50662 26936 50668
rect 26516 50380 26568 50386
rect 26516 50322 26568 50328
rect 26240 50176 26292 50182
rect 26240 50118 26292 50124
rect 26252 49842 26280 50118
rect 26240 49836 26292 49842
rect 26240 49778 26292 49784
rect 26056 49088 26108 49094
rect 26056 49030 26108 49036
rect 26240 49088 26292 49094
rect 26240 49030 26292 49036
rect 26068 47666 26096 49030
rect 26252 48754 26280 49030
rect 26240 48748 26292 48754
rect 26240 48690 26292 48696
rect 26332 48544 26384 48550
rect 26332 48486 26384 48492
rect 26344 48142 26372 48486
rect 26424 48204 26476 48210
rect 26424 48146 26476 48152
rect 26332 48136 26384 48142
rect 26332 48078 26384 48084
rect 26240 48000 26292 48006
rect 26240 47942 26292 47948
rect 26056 47660 26108 47666
rect 26056 47602 26108 47608
rect 26068 47462 26096 47602
rect 26056 47456 26108 47462
rect 26056 47398 26108 47404
rect 26252 47054 26280 47942
rect 26436 47802 26464 48146
rect 26424 47796 26476 47802
rect 26424 47738 26476 47744
rect 26424 47252 26476 47258
rect 26424 47194 26476 47200
rect 26436 47054 26464 47194
rect 26240 47048 26292 47054
rect 26240 46990 26292 46996
rect 26424 47048 26476 47054
rect 26424 46990 26476 46996
rect 26240 46912 26292 46918
rect 26240 46854 26292 46860
rect 26252 46646 26280 46854
rect 26240 46640 26292 46646
rect 26240 46582 26292 46588
rect 26528 46578 26556 50322
rect 26700 50312 26752 50318
rect 26700 50254 26752 50260
rect 26792 50312 26844 50318
rect 26792 50254 26844 50260
rect 26608 48680 26660 48686
rect 26608 48622 26660 48628
rect 26620 47530 26648 48622
rect 26608 47524 26660 47530
rect 26608 47466 26660 47472
rect 26516 46572 26568 46578
rect 26516 46514 26568 46520
rect 26712 46374 26740 50254
rect 26804 49978 26832 50254
rect 26792 49972 26844 49978
rect 26792 49914 26844 49920
rect 26896 49824 26924 50662
rect 27172 50522 27200 53450
rect 27712 52488 27764 52494
rect 27712 52430 27764 52436
rect 27344 52352 27396 52358
rect 27344 52294 27396 52300
rect 27356 51406 27384 52294
rect 27724 52154 27752 52430
rect 27712 52148 27764 52154
rect 27712 52090 27764 52096
rect 27620 51944 27672 51950
rect 27620 51886 27672 51892
rect 27632 51610 27660 51886
rect 27620 51604 27672 51610
rect 27620 51546 27672 51552
rect 27344 51400 27396 51406
rect 27344 51342 27396 51348
rect 27252 51332 27304 51338
rect 27252 51274 27304 51280
rect 27160 50516 27212 50522
rect 27160 50458 27212 50464
rect 26976 50312 27028 50318
rect 26976 50254 27028 50260
rect 26804 49796 26924 49824
rect 26804 49094 26832 49796
rect 26884 49156 26936 49162
rect 26884 49098 26936 49104
rect 26792 49088 26844 49094
rect 26792 49030 26844 49036
rect 26804 48686 26832 49030
rect 26896 48754 26924 49098
rect 26884 48748 26936 48754
rect 26884 48690 26936 48696
rect 26792 48680 26844 48686
rect 26792 48622 26844 48628
rect 26988 47258 27016 50254
rect 27264 48278 27292 51274
rect 27528 51264 27580 51270
rect 27528 51206 27580 51212
rect 27540 50386 27568 51206
rect 27908 51074 27936 54606
rect 28080 53984 28132 53990
rect 28080 53926 28132 53932
rect 28092 53582 28120 53926
rect 28080 53576 28132 53582
rect 28080 53518 28132 53524
rect 28092 53038 28120 53518
rect 28184 53446 28212 54606
rect 30104 54528 30156 54534
rect 30104 54470 30156 54476
rect 28264 54188 28316 54194
rect 28264 54130 28316 54136
rect 29460 54188 29512 54194
rect 29460 54130 29512 54136
rect 28172 53440 28224 53446
rect 28172 53382 28224 53388
rect 27988 53032 28040 53038
rect 27988 52974 28040 52980
rect 28080 53032 28132 53038
rect 28080 52974 28132 52980
rect 28000 52630 28028 52974
rect 27988 52624 28040 52630
rect 27988 52566 28040 52572
rect 27988 52012 28040 52018
rect 28092 52000 28120 52974
rect 28040 51972 28120 52000
rect 27988 51954 28040 51960
rect 27816 51046 27936 51074
rect 27528 50380 27580 50386
rect 27528 50322 27580 50328
rect 27620 49768 27672 49774
rect 27620 49710 27672 49716
rect 27528 48612 27580 48618
rect 27528 48554 27580 48560
rect 27252 48272 27304 48278
rect 27252 48214 27304 48220
rect 27540 48142 27568 48554
rect 27528 48136 27580 48142
rect 27528 48078 27580 48084
rect 27160 47660 27212 47666
rect 27160 47602 27212 47608
rect 27436 47660 27488 47666
rect 27436 47602 27488 47608
rect 26976 47252 27028 47258
rect 26976 47194 27028 47200
rect 27172 47054 27200 47602
rect 27448 47054 27476 47602
rect 27160 47048 27212 47054
rect 27160 46990 27212 46996
rect 27436 47048 27488 47054
rect 27436 46990 27488 46996
rect 27632 46986 27660 49710
rect 27712 48680 27764 48686
rect 27712 48622 27764 48628
rect 27724 47122 27752 48622
rect 27712 47116 27764 47122
rect 27712 47058 27764 47064
rect 27620 46980 27672 46986
rect 27620 46922 27672 46928
rect 27528 46640 27580 46646
rect 27528 46582 27580 46588
rect 26424 46368 26476 46374
rect 26424 46310 26476 46316
rect 26700 46368 26752 46374
rect 26700 46310 26752 46316
rect 27436 46368 27488 46374
rect 27436 46310 27488 46316
rect 26332 45960 26384 45966
rect 26332 45902 26384 45908
rect 26344 45558 26372 45902
rect 26332 45552 26384 45558
rect 26332 45494 26384 45500
rect 26436 44810 26464 46310
rect 27448 45966 27476 46310
rect 27436 45960 27488 45966
rect 27436 45902 27488 45908
rect 26700 45824 26752 45830
rect 26700 45766 26752 45772
rect 26712 45490 26740 45766
rect 27540 45626 27568 46582
rect 27528 45620 27580 45626
rect 27528 45562 27580 45568
rect 26700 45484 26752 45490
rect 26700 45426 26752 45432
rect 26424 44804 26476 44810
rect 26424 44746 26476 44752
rect 26148 44260 26200 44266
rect 26148 44202 26200 44208
rect 26160 43926 26188 44202
rect 26240 44192 26292 44198
rect 26240 44134 26292 44140
rect 26148 43920 26200 43926
rect 26148 43862 26200 43868
rect 26252 42566 26280 44134
rect 26436 43330 26464 44746
rect 26436 43302 26556 43330
rect 26424 43240 26476 43246
rect 26424 43182 26476 43188
rect 26240 42560 26292 42566
rect 26240 42502 26292 42508
rect 26252 42158 26280 42502
rect 26332 42356 26384 42362
rect 26332 42298 26384 42304
rect 26240 42152 26292 42158
rect 26240 42094 26292 42100
rect 25976 41386 26188 41414
rect 25504 41268 25556 41274
rect 25504 41210 25556 41216
rect 26056 41200 26108 41206
rect 26056 41142 26108 41148
rect 25320 41132 25372 41138
rect 25320 41074 25372 41080
rect 24400 40928 24452 40934
rect 24400 40870 24452 40876
rect 25044 40928 25096 40934
rect 25044 40870 25096 40876
rect 24412 40594 24440 40870
rect 24400 40588 24452 40594
rect 24400 40530 24452 40536
rect 24584 40520 24636 40526
rect 24584 40462 24636 40468
rect 24596 40050 24624 40462
rect 24584 40044 24636 40050
rect 24584 39986 24636 39992
rect 24952 39976 25004 39982
rect 24952 39918 25004 39924
rect 24964 39846 24992 39918
rect 24492 39840 24544 39846
rect 24492 39782 24544 39788
rect 24952 39840 25004 39846
rect 24952 39782 25004 39788
rect 24504 39438 24532 39782
rect 24964 39522 24992 39782
rect 24872 39494 24992 39522
rect 24872 39438 24900 39494
rect 24492 39432 24544 39438
rect 24492 39374 24544 39380
rect 24860 39432 24912 39438
rect 24860 39374 24912 39380
rect 24952 39432 25004 39438
rect 24952 39374 25004 39380
rect 24308 39296 24360 39302
rect 24308 39238 24360 39244
rect 24400 38752 24452 38758
rect 24400 38694 24452 38700
rect 24412 38350 24440 38694
rect 24400 38344 24452 38350
rect 24400 38286 24452 38292
rect 24308 37868 24360 37874
rect 24308 37810 24360 37816
rect 24320 37398 24348 37810
rect 24308 37392 24360 37398
rect 24308 37334 24360 37340
rect 24320 37194 24348 37334
rect 24504 37262 24532 39374
rect 24872 38962 24900 39374
rect 24964 39030 24992 39374
rect 24952 39024 25004 39030
rect 24952 38966 25004 38972
rect 24860 38956 24912 38962
rect 24860 38898 24912 38904
rect 24676 38752 24728 38758
rect 24676 38694 24728 38700
rect 24688 38282 24716 38694
rect 24676 38276 24728 38282
rect 24676 38218 24728 38224
rect 24688 37806 24716 38218
rect 24768 38208 24820 38214
rect 24768 38150 24820 38156
rect 24780 37874 24808 38150
rect 24768 37868 24820 37874
rect 24768 37810 24820 37816
rect 24676 37800 24728 37806
rect 24676 37742 24728 37748
rect 24676 37664 24728 37670
rect 24676 37606 24728 37612
rect 24688 37262 24716 37606
rect 24492 37256 24544 37262
rect 24492 37198 24544 37204
rect 24676 37256 24728 37262
rect 24676 37198 24728 37204
rect 24308 37188 24360 37194
rect 24308 37130 24360 37136
rect 24216 37120 24268 37126
rect 24216 37062 24268 37068
rect 24228 35698 24256 37062
rect 24320 36786 24348 37130
rect 24400 37120 24452 37126
rect 24400 37062 24452 37068
rect 24584 37120 24636 37126
rect 24584 37062 24636 37068
rect 24308 36780 24360 36786
rect 24308 36722 24360 36728
rect 24124 35692 24176 35698
rect 24124 35634 24176 35640
rect 24216 35692 24268 35698
rect 24216 35634 24268 35640
rect 24136 35222 24164 35634
rect 24412 35290 24440 37062
rect 24596 36174 24624 37062
rect 24780 36786 24808 37810
rect 24860 37256 24912 37262
rect 24860 37198 24912 37204
rect 24872 36922 24900 37198
rect 24860 36916 24912 36922
rect 24860 36858 24912 36864
rect 24768 36780 24820 36786
rect 24768 36722 24820 36728
rect 24768 36576 24820 36582
rect 24768 36518 24820 36524
rect 24780 36174 24808 36518
rect 24584 36168 24636 36174
rect 24584 36110 24636 36116
rect 24768 36168 24820 36174
rect 24768 36110 24820 36116
rect 24768 35692 24820 35698
rect 24768 35634 24820 35640
rect 24584 35488 24636 35494
rect 24584 35430 24636 35436
rect 24400 35284 24452 35290
rect 24400 35226 24452 35232
rect 24124 35216 24176 35222
rect 24124 35158 24176 35164
rect 24596 34932 24624 35430
rect 24780 35290 24808 35634
rect 25056 35562 25084 40870
rect 26068 40526 26096 41142
rect 26056 40520 26108 40526
rect 26056 40462 26108 40468
rect 25780 40384 25832 40390
rect 25780 40326 25832 40332
rect 25792 40186 25820 40326
rect 25780 40180 25832 40186
rect 25780 40122 25832 40128
rect 25504 39840 25556 39846
rect 25504 39782 25556 39788
rect 25516 39574 25544 39782
rect 25504 39568 25556 39574
rect 25504 39510 25556 39516
rect 25136 39296 25188 39302
rect 25136 39238 25188 39244
rect 25148 37194 25176 39238
rect 25228 38956 25280 38962
rect 25228 38898 25280 38904
rect 25240 38826 25268 38898
rect 25228 38820 25280 38826
rect 25228 38762 25280 38768
rect 25320 38480 25372 38486
rect 25320 38422 25372 38428
rect 25228 38208 25280 38214
rect 25228 38150 25280 38156
rect 25240 38010 25268 38150
rect 25228 38004 25280 38010
rect 25228 37946 25280 37952
rect 25332 37806 25360 38422
rect 26056 38344 26108 38350
rect 26056 38286 26108 38292
rect 26068 38010 26096 38286
rect 26056 38004 26108 38010
rect 26056 37946 26108 37952
rect 25412 37868 25464 37874
rect 25412 37810 25464 37816
rect 25320 37800 25372 37806
rect 25320 37742 25372 37748
rect 25136 37188 25188 37194
rect 25136 37130 25188 37136
rect 25228 37188 25280 37194
rect 25228 37130 25280 37136
rect 25240 36718 25268 37130
rect 25228 36712 25280 36718
rect 25228 36654 25280 36660
rect 25332 35834 25360 37742
rect 25424 37262 25452 37810
rect 25412 37256 25464 37262
rect 25412 37198 25464 37204
rect 26160 36922 26188 41386
rect 26344 41206 26372 42298
rect 26332 41200 26384 41206
rect 26332 41142 26384 41148
rect 26240 40996 26292 41002
rect 26240 40938 26292 40944
rect 26252 40390 26280 40938
rect 26332 40928 26384 40934
rect 26332 40870 26384 40876
rect 26344 40594 26372 40870
rect 26332 40588 26384 40594
rect 26332 40530 26384 40536
rect 26240 40384 26292 40390
rect 26240 40326 26292 40332
rect 26344 40050 26372 40530
rect 26332 40044 26384 40050
rect 26252 40004 26332 40032
rect 26252 39098 26280 40004
rect 26332 39986 26384 39992
rect 26436 39370 26464 43182
rect 26528 43178 26556 43302
rect 26516 43172 26568 43178
rect 26516 43114 26568 43120
rect 26608 41472 26660 41478
rect 26608 41414 26660 41420
rect 26516 41200 26568 41206
rect 26516 41142 26568 41148
rect 26528 40934 26556 41142
rect 26516 40928 26568 40934
rect 26516 40870 26568 40876
rect 26620 40594 26648 41414
rect 26608 40588 26660 40594
rect 26608 40530 26660 40536
rect 26516 40384 26568 40390
rect 26516 40326 26568 40332
rect 26528 39370 26556 40326
rect 26608 40112 26660 40118
rect 26608 40054 26660 40060
rect 26424 39364 26476 39370
rect 26424 39306 26476 39312
rect 26516 39364 26568 39370
rect 26516 39306 26568 39312
rect 26332 39296 26384 39302
rect 26332 39238 26384 39244
rect 26344 39098 26372 39238
rect 26240 39092 26292 39098
rect 26240 39034 26292 39040
rect 26332 39092 26384 39098
rect 26332 39034 26384 39040
rect 26332 38752 26384 38758
rect 26332 38694 26384 38700
rect 26148 36916 26200 36922
rect 26148 36858 26200 36864
rect 25412 36712 25464 36718
rect 25412 36654 25464 36660
rect 25424 36378 25452 36654
rect 26240 36644 26292 36650
rect 26240 36586 26292 36592
rect 25872 36576 25924 36582
rect 25872 36518 25924 36524
rect 25412 36372 25464 36378
rect 25412 36314 25464 36320
rect 25884 36242 25912 36518
rect 25872 36236 25924 36242
rect 25872 36178 25924 36184
rect 26252 35834 26280 36586
rect 26344 36582 26372 38694
rect 26436 37874 26464 39306
rect 26528 39030 26556 39306
rect 26516 39024 26568 39030
rect 26516 38966 26568 38972
rect 26528 38554 26556 38966
rect 26516 38548 26568 38554
rect 26516 38490 26568 38496
rect 26620 38400 26648 40054
rect 26712 38570 26740 45426
rect 26884 45416 26936 45422
rect 26884 45358 26936 45364
rect 26896 44810 26924 45358
rect 27816 45354 27844 51046
rect 27896 49224 27948 49230
rect 27896 49166 27948 49172
rect 27908 47734 27936 49166
rect 27896 47728 27948 47734
rect 27896 47670 27948 47676
rect 28000 46034 28028 51954
rect 28184 50250 28212 53382
rect 28172 50244 28224 50250
rect 28172 50186 28224 50192
rect 28080 49768 28132 49774
rect 28080 49710 28132 49716
rect 28092 49094 28120 49710
rect 28080 49088 28132 49094
rect 28132 49048 28212 49076
rect 28080 49030 28132 49036
rect 28184 48142 28212 49048
rect 28276 48890 28304 54130
rect 28908 53984 28960 53990
rect 28908 53926 28960 53932
rect 28816 53440 28868 53446
rect 28816 53382 28868 53388
rect 28828 53106 28856 53382
rect 28816 53100 28868 53106
rect 28816 53042 28868 53048
rect 28724 52896 28776 52902
rect 28724 52838 28776 52844
rect 28736 52494 28764 52838
rect 28724 52488 28776 52494
rect 28724 52430 28776 52436
rect 28816 52488 28868 52494
rect 28920 52442 28948 53926
rect 29472 53650 29500 54130
rect 30116 54126 30144 54470
rect 30104 54120 30156 54126
rect 30104 54062 30156 54068
rect 29552 53984 29604 53990
rect 29552 53926 29604 53932
rect 29460 53644 29512 53650
rect 29460 53586 29512 53592
rect 29368 53508 29420 53514
rect 29368 53450 29420 53456
rect 29000 53032 29052 53038
rect 29000 52974 29052 52980
rect 29012 52698 29040 52974
rect 29000 52692 29052 52698
rect 29000 52634 29052 52640
rect 29380 52494 29408 53450
rect 28868 52436 28948 52442
rect 28816 52430 28948 52436
rect 29368 52488 29420 52494
rect 29368 52430 29420 52436
rect 28828 52414 28948 52430
rect 29000 52420 29052 52426
rect 28724 51808 28776 51814
rect 28724 51750 28776 51756
rect 28736 50794 28764 51750
rect 28828 51610 28856 52414
rect 29000 52362 29052 52368
rect 28816 51604 28868 51610
rect 28816 51546 28868 51552
rect 28828 51406 28856 51546
rect 28816 51400 28868 51406
rect 28816 51342 28868 51348
rect 28724 50788 28776 50794
rect 28724 50730 28776 50736
rect 28908 50720 28960 50726
rect 28908 50662 28960 50668
rect 28920 50182 28948 50662
rect 28908 50176 28960 50182
rect 28908 50118 28960 50124
rect 28540 49224 28592 49230
rect 28540 49166 28592 49172
rect 28448 49088 28500 49094
rect 28448 49030 28500 49036
rect 28264 48884 28316 48890
rect 28264 48826 28316 48832
rect 28356 48748 28408 48754
rect 28356 48690 28408 48696
rect 28368 48142 28396 48690
rect 28460 48686 28488 49030
rect 28448 48680 28500 48686
rect 28448 48622 28500 48628
rect 28552 48142 28580 49166
rect 28816 49088 28868 49094
rect 28816 49030 28868 49036
rect 28828 48754 28856 49030
rect 28816 48748 28868 48754
rect 28816 48690 28868 48696
rect 28920 48210 28948 50118
rect 28908 48204 28960 48210
rect 28908 48146 28960 48152
rect 28172 48136 28224 48142
rect 28356 48136 28408 48142
rect 28224 48084 28304 48090
rect 28172 48078 28304 48084
rect 28356 48078 28408 48084
rect 28540 48136 28592 48142
rect 28540 48078 28592 48084
rect 28632 48136 28684 48142
rect 28632 48078 28684 48084
rect 28184 48062 28304 48078
rect 28276 46374 28304 48062
rect 28644 47734 28672 48078
rect 28632 47728 28684 47734
rect 28632 47670 28684 47676
rect 28920 47598 28948 48146
rect 29012 47802 29040 52362
rect 29472 52086 29500 53586
rect 29564 53514 29592 53926
rect 30012 53644 30064 53650
rect 30012 53586 30064 53592
rect 29552 53508 29604 53514
rect 29552 53450 29604 53456
rect 29564 52562 29592 53450
rect 29552 52556 29604 52562
rect 29552 52498 29604 52504
rect 29828 52488 29880 52494
rect 29828 52430 29880 52436
rect 29840 52154 29868 52430
rect 29828 52148 29880 52154
rect 29828 52090 29880 52096
rect 29460 52080 29512 52086
rect 29460 52022 29512 52028
rect 30024 52018 30052 53586
rect 30116 52902 30144 54062
rect 30104 52896 30156 52902
rect 30104 52838 30156 52844
rect 30116 52086 30144 52838
rect 30288 52488 30340 52494
rect 30288 52430 30340 52436
rect 30104 52080 30156 52086
rect 30104 52022 30156 52028
rect 30012 52012 30064 52018
rect 30012 51954 30064 51960
rect 30012 51332 30064 51338
rect 30012 51274 30064 51280
rect 29828 51264 29880 51270
rect 29828 51206 29880 51212
rect 29276 50720 29328 50726
rect 29276 50662 29328 50668
rect 29288 50386 29316 50662
rect 29276 50380 29328 50386
rect 29276 50322 29328 50328
rect 29288 48822 29316 50322
rect 29736 49836 29788 49842
rect 29736 49778 29788 49784
rect 29368 49632 29420 49638
rect 29368 49574 29420 49580
rect 29276 48816 29328 48822
rect 29276 48758 29328 48764
rect 29184 48612 29236 48618
rect 29184 48554 29236 48560
rect 29000 47796 29052 47802
rect 29000 47738 29052 47744
rect 29196 47666 29224 48554
rect 29288 48142 29316 48758
rect 29380 48550 29408 49574
rect 29748 49434 29776 49778
rect 29736 49428 29788 49434
rect 29736 49370 29788 49376
rect 29840 49314 29868 51206
rect 30024 50998 30052 51274
rect 30012 50992 30064 50998
rect 30012 50934 30064 50940
rect 30300 50930 30328 52430
rect 30380 50992 30432 50998
rect 30380 50934 30432 50940
rect 30288 50924 30340 50930
rect 30288 50866 30340 50872
rect 30104 50720 30156 50726
rect 30104 50662 30156 50668
rect 30116 50318 30144 50662
rect 30300 50522 30328 50866
rect 30288 50516 30340 50522
rect 30288 50458 30340 50464
rect 30104 50312 30156 50318
rect 30104 50254 30156 50260
rect 29920 50176 29972 50182
rect 29920 50118 29972 50124
rect 29932 49366 29960 50118
rect 30300 49842 30328 50458
rect 30392 50386 30420 50934
rect 30380 50380 30432 50386
rect 30380 50322 30432 50328
rect 30288 49836 30340 49842
rect 30288 49778 30340 49784
rect 30012 49768 30064 49774
rect 30012 49710 30064 49716
rect 29748 49286 29868 49314
rect 29920 49360 29972 49366
rect 29920 49302 29972 49308
rect 29748 49230 29776 49286
rect 29552 49224 29604 49230
rect 29552 49166 29604 49172
rect 29736 49224 29788 49230
rect 29736 49166 29788 49172
rect 29828 49224 29880 49230
rect 29828 49166 29880 49172
rect 29564 49094 29592 49166
rect 29552 49088 29604 49094
rect 29552 49030 29604 49036
rect 29564 48754 29592 49030
rect 29552 48748 29604 48754
rect 29552 48690 29604 48696
rect 29748 48686 29776 49166
rect 29736 48680 29788 48686
rect 29736 48622 29788 48628
rect 29368 48544 29420 48550
rect 29368 48486 29420 48492
rect 29380 48314 29408 48486
rect 29840 48346 29868 49166
rect 29920 48544 29972 48550
rect 29920 48486 29972 48492
rect 29828 48340 29880 48346
rect 29380 48286 29500 48314
rect 29276 48136 29328 48142
rect 29472 48113 29500 48286
rect 29828 48282 29880 48288
rect 29932 48210 29960 48486
rect 29920 48204 29972 48210
rect 29920 48146 29972 48152
rect 29276 48078 29328 48084
rect 29458 48104 29514 48113
rect 29288 47734 29316 48078
rect 29458 48039 29514 48048
rect 29276 47728 29328 47734
rect 29276 47670 29328 47676
rect 29184 47660 29236 47666
rect 29184 47602 29236 47608
rect 29368 47660 29420 47666
rect 29368 47602 29420 47608
rect 28908 47592 28960 47598
rect 28908 47534 28960 47540
rect 28540 47456 28592 47462
rect 28540 47398 28592 47404
rect 28552 47122 28580 47398
rect 28920 47190 28948 47534
rect 29380 47258 29408 47602
rect 29368 47252 29420 47258
rect 29368 47194 29420 47200
rect 28908 47184 28960 47190
rect 28908 47126 28960 47132
rect 28540 47116 28592 47122
rect 28540 47058 28592 47064
rect 28448 46980 28500 46986
rect 28448 46922 28500 46928
rect 28264 46368 28316 46374
rect 28264 46310 28316 46316
rect 27988 46028 28040 46034
rect 27988 45970 28040 45976
rect 27804 45348 27856 45354
rect 27804 45290 27856 45296
rect 27528 45280 27580 45286
rect 27528 45222 27580 45228
rect 27540 45082 27568 45222
rect 27528 45076 27580 45082
rect 27528 45018 27580 45024
rect 26884 44804 26936 44810
rect 26884 44746 26936 44752
rect 26792 44396 26844 44402
rect 26792 44338 26844 44344
rect 26804 42702 26832 44338
rect 26792 42696 26844 42702
rect 26792 42638 26844 42644
rect 26792 42084 26844 42090
rect 26792 42026 26844 42032
rect 26804 41138 26832 42026
rect 26896 41596 26924 44746
rect 27160 44736 27212 44742
rect 27160 44678 27212 44684
rect 27172 44538 27200 44678
rect 27160 44532 27212 44538
rect 27160 44474 27212 44480
rect 27540 44402 27568 45018
rect 27712 44872 27764 44878
rect 27712 44814 27764 44820
rect 27528 44396 27580 44402
rect 27528 44338 27580 44344
rect 27068 43308 27120 43314
rect 27068 43250 27120 43256
rect 27080 42906 27108 43250
rect 27252 43104 27304 43110
rect 27252 43046 27304 43052
rect 27344 43104 27396 43110
rect 27344 43046 27396 43052
rect 27068 42900 27120 42906
rect 27068 42842 27120 42848
rect 27264 42838 27292 43046
rect 27252 42832 27304 42838
rect 27252 42774 27304 42780
rect 27252 42696 27304 42702
rect 27252 42638 27304 42644
rect 27066 41712 27122 41721
rect 27066 41647 27122 41656
rect 26896 41568 27016 41596
rect 26884 41472 26936 41478
rect 26884 41414 26936 41420
rect 26896 41274 26924 41414
rect 26884 41268 26936 41274
rect 26884 41210 26936 41216
rect 26988 41154 27016 41568
rect 27080 41478 27108 41647
rect 27068 41472 27120 41478
rect 27068 41414 27120 41420
rect 27264 41426 27292 42638
rect 27356 42362 27384 43046
rect 27540 42838 27568 44338
rect 27724 43450 27752 44814
rect 28000 44470 28028 45970
rect 28080 45552 28132 45558
rect 28080 45494 28132 45500
rect 27988 44464 28040 44470
rect 27988 44406 28040 44412
rect 28092 44334 28120 45494
rect 28276 45082 28304 46310
rect 28356 45824 28408 45830
rect 28356 45766 28408 45772
rect 28368 45286 28396 45766
rect 28460 45286 28488 46922
rect 28920 45558 28948 47126
rect 29472 47122 29500 48039
rect 29920 48000 29972 48006
rect 29920 47942 29972 47948
rect 29000 47116 29052 47122
rect 29000 47058 29052 47064
rect 29460 47116 29512 47122
rect 29460 47058 29512 47064
rect 29012 46374 29040 47058
rect 29552 47048 29604 47054
rect 29552 46990 29604 46996
rect 29184 46980 29236 46986
rect 29184 46922 29236 46928
rect 29196 46714 29224 46922
rect 29184 46708 29236 46714
rect 29184 46650 29236 46656
rect 29460 46640 29512 46646
rect 29460 46582 29512 46588
rect 29000 46368 29052 46374
rect 29000 46310 29052 46316
rect 29472 45898 29500 46582
rect 29564 46170 29592 46990
rect 29932 46646 29960 47942
rect 29920 46640 29972 46646
rect 29920 46582 29972 46588
rect 29736 46572 29788 46578
rect 29736 46514 29788 46520
rect 29828 46572 29880 46578
rect 29828 46514 29880 46520
rect 29552 46164 29604 46170
rect 29552 46106 29604 46112
rect 29748 45966 29776 46514
rect 29840 46374 29868 46514
rect 29828 46368 29880 46374
rect 29828 46310 29880 46316
rect 29840 45966 29868 46310
rect 29736 45960 29788 45966
rect 29736 45902 29788 45908
rect 29828 45960 29880 45966
rect 29828 45902 29880 45908
rect 29460 45892 29512 45898
rect 29460 45834 29512 45840
rect 28908 45552 28960 45558
rect 28908 45494 28960 45500
rect 28356 45280 28408 45286
rect 28356 45222 28408 45228
rect 28448 45280 28500 45286
rect 28448 45222 28500 45228
rect 29000 45280 29052 45286
rect 29000 45222 29052 45228
rect 28264 45076 28316 45082
rect 28264 45018 28316 45024
rect 28276 44810 28304 45018
rect 28264 44804 28316 44810
rect 28264 44746 28316 44752
rect 28172 44736 28224 44742
rect 28172 44678 28224 44684
rect 28080 44328 28132 44334
rect 28080 44270 28132 44276
rect 27712 43444 27764 43450
rect 27712 43386 27764 43392
rect 28092 42838 28120 44270
rect 27528 42832 27580 42838
rect 27528 42774 27580 42780
rect 28080 42832 28132 42838
rect 28080 42774 28132 42780
rect 27436 42696 27488 42702
rect 27436 42638 27488 42644
rect 27344 42356 27396 42362
rect 27344 42298 27396 42304
rect 27356 42226 27384 42298
rect 27344 42220 27396 42226
rect 27344 42162 27396 42168
rect 27448 41750 27476 42638
rect 27540 42226 27568 42774
rect 27712 42560 27764 42566
rect 27712 42502 27764 42508
rect 27724 42294 27752 42502
rect 27712 42288 27764 42294
rect 27712 42230 27764 42236
rect 27528 42220 27580 42226
rect 27528 42162 27580 42168
rect 27896 42016 27948 42022
rect 27896 41958 27948 41964
rect 27436 41744 27488 41750
rect 27436 41686 27488 41692
rect 27342 41440 27398 41449
rect 27264 41398 27342 41426
rect 27342 41375 27398 41384
rect 26792 41132 26844 41138
rect 26792 41074 26844 41080
rect 26896 41126 27016 41154
rect 26804 40526 26832 41074
rect 26896 41002 26924 41126
rect 26976 41064 27028 41070
rect 26976 41006 27028 41012
rect 27252 41064 27304 41070
rect 27252 41006 27304 41012
rect 26884 40996 26936 41002
rect 26884 40938 26936 40944
rect 26792 40520 26844 40526
rect 26792 40462 26844 40468
rect 26884 40452 26936 40458
rect 26884 40394 26936 40400
rect 26896 39642 26924 40394
rect 26884 39636 26936 39642
rect 26884 39578 26936 39584
rect 26988 39506 27016 41006
rect 27160 40928 27212 40934
rect 27160 40870 27212 40876
rect 27068 40180 27120 40186
rect 27068 40122 27120 40128
rect 27080 39982 27108 40122
rect 27172 40118 27200 40870
rect 27264 40730 27292 41006
rect 27252 40724 27304 40730
rect 27252 40666 27304 40672
rect 27356 40458 27384 41375
rect 27344 40452 27396 40458
rect 27344 40394 27396 40400
rect 27160 40112 27212 40118
rect 27160 40054 27212 40060
rect 27344 40044 27396 40050
rect 27264 40004 27344 40032
rect 27068 39976 27120 39982
rect 27068 39918 27120 39924
rect 27160 39840 27212 39846
rect 27160 39782 27212 39788
rect 26976 39500 27028 39506
rect 26976 39442 27028 39448
rect 26712 38542 26832 38570
rect 26700 38480 26752 38486
rect 26700 38422 26752 38428
rect 26528 38372 26648 38400
rect 26424 37868 26476 37874
rect 26424 37810 26476 37816
rect 26436 37330 26464 37810
rect 26424 37324 26476 37330
rect 26424 37266 26476 37272
rect 26528 36718 26556 38372
rect 26608 38276 26660 38282
rect 26608 38218 26660 38224
rect 26620 37738 26648 38218
rect 26712 37806 26740 38422
rect 26700 37800 26752 37806
rect 26700 37742 26752 37748
rect 26608 37732 26660 37738
rect 26608 37674 26660 37680
rect 26620 37466 26648 37674
rect 26700 37664 26752 37670
rect 26700 37606 26752 37612
rect 26608 37460 26660 37466
rect 26608 37402 26660 37408
rect 26712 37398 26740 37606
rect 26700 37392 26752 37398
rect 26700 37334 26752 37340
rect 26516 36712 26568 36718
rect 26516 36654 26568 36660
rect 26332 36576 26384 36582
rect 26332 36518 26384 36524
rect 26344 36174 26372 36518
rect 26332 36168 26384 36174
rect 26332 36110 26384 36116
rect 25320 35828 25372 35834
rect 25320 35770 25372 35776
rect 26240 35828 26292 35834
rect 26240 35770 26292 35776
rect 25044 35556 25096 35562
rect 25044 35498 25096 35504
rect 24768 35284 24820 35290
rect 24768 35226 24820 35232
rect 25044 35012 25096 35018
rect 25044 34954 25096 34960
rect 24596 34904 24716 34932
rect 24688 34610 24716 34904
rect 25056 34678 25084 34954
rect 25332 34746 25360 35770
rect 25872 35216 25924 35222
rect 25872 35158 25924 35164
rect 25780 34944 25832 34950
rect 25780 34886 25832 34892
rect 25320 34740 25372 34746
rect 25320 34682 25372 34688
rect 25044 34672 25096 34678
rect 25044 34614 25096 34620
rect 24676 34604 24728 34610
rect 24676 34546 24728 34552
rect 24860 34604 24912 34610
rect 24860 34546 24912 34552
rect 24688 34406 24716 34546
rect 24676 34400 24728 34406
rect 24676 34342 24728 34348
rect 24688 34066 24716 34342
rect 24872 34134 24900 34546
rect 24860 34128 24912 34134
rect 24860 34070 24912 34076
rect 24676 34060 24728 34066
rect 24676 34002 24728 34008
rect 24492 33856 24544 33862
rect 24492 33798 24544 33804
rect 24504 33590 24532 33798
rect 24688 33658 24716 34002
rect 24676 33652 24728 33658
rect 24676 33594 24728 33600
rect 24492 33584 24544 33590
rect 24492 33526 24544 33532
rect 24492 33380 24544 33386
rect 24492 33322 24544 33328
rect 24504 32978 24532 33322
rect 24492 32972 24544 32978
rect 24492 32914 24544 32920
rect 24400 32428 24452 32434
rect 24504 32416 24532 32914
rect 24452 32388 24532 32416
rect 24400 32370 24452 32376
rect 24676 32224 24728 32230
rect 24676 32166 24728 32172
rect 24032 31884 24084 31890
rect 24032 31826 24084 31832
rect 24688 31414 24716 32166
rect 24676 31408 24728 31414
rect 24676 31350 24728 31356
rect 24216 31136 24268 31142
rect 24216 31078 24268 31084
rect 24584 31136 24636 31142
rect 24584 31078 24636 31084
rect 23940 30184 23992 30190
rect 23940 30126 23992 30132
rect 23756 29844 23808 29850
rect 23756 29786 23808 29792
rect 23676 29702 23796 29730
rect 23768 29578 23796 29702
rect 23848 29640 23900 29646
rect 23848 29582 23900 29588
rect 23756 29572 23808 29578
rect 23756 29514 23808 29520
rect 23480 29300 23532 29306
rect 23480 29242 23532 29248
rect 23296 29096 23348 29102
rect 23296 29038 23348 29044
rect 23664 28688 23716 28694
rect 23664 28630 23716 28636
rect 23388 28484 23440 28490
rect 23388 28426 23440 28432
rect 23400 28218 23428 28426
rect 23388 28212 23440 28218
rect 23388 28154 23440 28160
rect 23676 28150 23704 28630
rect 23664 28144 23716 28150
rect 23664 28086 23716 28092
rect 23388 28076 23440 28082
rect 23216 28036 23388 28064
rect 23112 28018 23164 28024
rect 23388 28018 23440 28024
rect 23204 27872 23256 27878
rect 23204 27814 23256 27820
rect 22652 27396 22704 27402
rect 22652 27338 22704 27344
rect 22192 26988 22244 26994
rect 22192 26930 22244 26936
rect 22284 26988 22336 26994
rect 22284 26930 22336 26936
rect 22560 26988 22612 26994
rect 22560 26930 22612 26936
rect 22204 26586 22232 26930
rect 22664 26926 22692 27338
rect 23216 27062 23244 27814
rect 23400 27674 23428 28018
rect 23388 27668 23440 27674
rect 23388 27610 23440 27616
rect 23676 27538 23704 28086
rect 23664 27532 23716 27538
rect 23664 27474 23716 27480
rect 23204 27056 23256 27062
rect 23204 26998 23256 27004
rect 22652 26920 22704 26926
rect 22652 26862 22704 26868
rect 22192 26580 22244 26586
rect 22192 26522 22244 26528
rect 21732 26444 21784 26450
rect 21732 26386 21784 26392
rect 21744 25498 21772 26386
rect 22468 26308 22520 26314
rect 22468 26250 22520 26256
rect 22192 25900 22244 25906
rect 22192 25842 22244 25848
rect 21732 25492 21784 25498
rect 21732 25434 21784 25440
rect 22204 25158 22232 25842
rect 22480 25702 22508 26250
rect 23676 25906 23704 27474
rect 23768 26314 23796 29514
rect 23860 29306 23888 29582
rect 23848 29300 23900 29306
rect 23848 29242 23900 29248
rect 23940 28416 23992 28422
rect 23940 28358 23992 28364
rect 24124 28416 24176 28422
rect 24124 28358 24176 28364
rect 23952 28218 23980 28358
rect 23940 28212 23992 28218
rect 23940 28154 23992 28160
rect 24136 28150 24164 28358
rect 24124 28144 24176 28150
rect 24124 28086 24176 28092
rect 24124 27464 24176 27470
rect 24124 27406 24176 27412
rect 24136 27130 24164 27406
rect 24124 27124 24176 27130
rect 24124 27066 24176 27072
rect 24228 26994 24256 31078
rect 24596 30734 24624 31078
rect 24952 30796 25004 30802
rect 24952 30738 25004 30744
rect 24584 30728 24636 30734
rect 24584 30670 24636 30676
rect 24768 30728 24820 30734
rect 24768 30670 24820 30676
rect 24400 30592 24452 30598
rect 24400 30534 24452 30540
rect 24412 30258 24440 30534
rect 24780 30394 24808 30670
rect 24768 30388 24820 30394
rect 24768 30330 24820 30336
rect 24400 30252 24452 30258
rect 24400 30194 24452 30200
rect 24860 30252 24912 30258
rect 24860 30194 24912 30200
rect 24872 29850 24900 30194
rect 24860 29844 24912 29850
rect 24860 29786 24912 29792
rect 24964 29714 24992 30738
rect 24952 29708 25004 29714
rect 24952 29650 25004 29656
rect 24860 29028 24912 29034
rect 24860 28970 24912 28976
rect 24584 28076 24636 28082
rect 24584 28018 24636 28024
rect 24216 26988 24268 26994
rect 24216 26930 24268 26936
rect 24492 26988 24544 26994
rect 24492 26930 24544 26936
rect 24504 26586 24532 26930
rect 24492 26580 24544 26586
rect 24492 26522 24544 26528
rect 24400 26376 24452 26382
rect 24400 26318 24452 26324
rect 23756 26308 23808 26314
rect 23756 26250 23808 26256
rect 23664 25900 23716 25906
rect 23664 25842 23716 25848
rect 22468 25696 22520 25702
rect 22468 25638 22520 25644
rect 22480 25158 22508 25638
rect 22192 25152 22244 25158
rect 22192 25094 22244 25100
rect 22468 25152 22520 25158
rect 22468 25094 22520 25100
rect 22204 24886 22232 25094
rect 22192 24880 22244 24886
rect 22192 24822 22244 24828
rect 22008 24812 22060 24818
rect 22008 24754 22060 24760
rect 22020 24342 22048 24754
rect 22008 24336 22060 24342
rect 22008 24278 22060 24284
rect 22204 2650 22232 24822
rect 22284 2848 22336 2854
rect 22284 2790 22336 2796
rect 21548 2644 21600 2650
rect 21548 2586 21600 2592
rect 22192 2644 22244 2650
rect 22192 2586 22244 2592
rect 22296 2446 22324 2790
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 22480 2038 22508 25094
rect 23768 2514 23796 26250
rect 24412 26042 24440 26318
rect 24400 26036 24452 26042
rect 24400 25978 24452 25984
rect 24596 25922 24624 28018
rect 24768 28008 24820 28014
rect 24872 27996 24900 28970
rect 24952 28960 25004 28966
rect 24952 28902 25004 28908
rect 24964 28082 24992 28902
rect 24952 28076 25004 28082
rect 24952 28018 25004 28024
rect 24820 27968 24900 27996
rect 24768 27950 24820 27956
rect 24964 27946 24992 28018
rect 24952 27940 25004 27946
rect 24952 27882 25004 27888
rect 24860 26376 24912 26382
rect 24860 26318 24912 26324
rect 24872 26042 24900 26318
rect 24860 26036 24912 26042
rect 24860 25978 24912 25984
rect 24504 25894 24624 25922
rect 24676 25900 24728 25906
rect 24504 25158 24532 25894
rect 24676 25842 24728 25848
rect 24584 25832 24636 25838
rect 24584 25774 24636 25780
rect 24492 25152 24544 25158
rect 24492 25094 24544 25100
rect 24596 24954 24624 25774
rect 24688 25498 24716 25842
rect 24676 25492 24728 25498
rect 24676 25434 24728 25440
rect 24584 24948 24636 24954
rect 24584 24890 24636 24896
rect 25056 22094 25084 34614
rect 25332 32502 25360 34682
rect 25792 34610 25820 34886
rect 25884 34678 25912 35158
rect 26424 34740 26476 34746
rect 26424 34682 26476 34688
rect 25872 34672 25924 34678
rect 25872 34614 25924 34620
rect 25504 34604 25556 34610
rect 25504 34546 25556 34552
rect 25780 34604 25832 34610
rect 25780 34546 25832 34552
rect 25516 34202 25544 34546
rect 26056 34536 26108 34542
rect 26056 34478 26108 34484
rect 26068 34202 26096 34478
rect 25504 34196 25556 34202
rect 25504 34138 25556 34144
rect 26056 34196 26108 34202
rect 26056 34138 26108 34144
rect 26240 34196 26292 34202
rect 26240 34138 26292 34144
rect 25780 33312 25832 33318
rect 25780 33254 25832 33260
rect 25792 32910 25820 33254
rect 25596 32904 25648 32910
rect 25596 32846 25648 32852
rect 25780 32904 25832 32910
rect 25780 32846 25832 32852
rect 25504 32768 25556 32774
rect 25504 32710 25556 32716
rect 25320 32496 25372 32502
rect 25320 32438 25372 32444
rect 25332 30870 25360 32438
rect 25516 32434 25544 32710
rect 25608 32570 25636 32846
rect 25792 32774 25820 32846
rect 25780 32768 25832 32774
rect 25780 32710 25832 32716
rect 25596 32564 25648 32570
rect 25596 32506 25648 32512
rect 25504 32428 25556 32434
rect 25504 32370 25556 32376
rect 25596 32224 25648 32230
rect 25596 32166 25648 32172
rect 25608 31754 25636 32166
rect 25872 31816 25924 31822
rect 25872 31758 25924 31764
rect 25596 31748 25648 31754
rect 25596 31690 25648 31696
rect 25504 31680 25556 31686
rect 25504 31622 25556 31628
rect 25516 31346 25544 31622
rect 25504 31340 25556 31346
rect 25504 31282 25556 31288
rect 25320 30864 25372 30870
rect 25320 30806 25372 30812
rect 25332 30190 25360 30806
rect 25320 30184 25372 30190
rect 25320 30126 25372 30132
rect 25516 30138 25544 31282
rect 25608 30258 25636 31690
rect 25884 31482 25912 31758
rect 25872 31476 25924 31482
rect 25872 31418 25924 31424
rect 25688 31340 25740 31346
rect 25688 31282 25740 31288
rect 25780 31340 25832 31346
rect 25780 31282 25832 31288
rect 25700 30938 25728 31282
rect 25688 30932 25740 30938
rect 25688 30874 25740 30880
rect 25792 30394 25820 31282
rect 26068 30938 26096 34138
rect 26252 33998 26280 34138
rect 26436 34134 26464 34682
rect 26424 34128 26476 34134
rect 26424 34070 26476 34076
rect 26240 33992 26292 33998
rect 26240 33934 26292 33940
rect 26252 33590 26280 33934
rect 26436 33930 26464 34070
rect 26424 33924 26476 33930
rect 26424 33866 26476 33872
rect 26528 33658 26556 36654
rect 26516 33652 26568 33658
rect 26516 33594 26568 33600
rect 26240 33584 26292 33590
rect 26240 33526 26292 33532
rect 26252 33046 26280 33526
rect 26424 33312 26476 33318
rect 26424 33254 26476 33260
rect 26240 33040 26292 33046
rect 26240 32982 26292 32988
rect 26436 32978 26464 33254
rect 26424 32972 26476 32978
rect 26424 32914 26476 32920
rect 26528 32910 26556 33594
rect 26516 32904 26568 32910
rect 26516 32846 26568 32852
rect 26148 32020 26200 32026
rect 26148 31962 26200 31968
rect 26160 31822 26188 31962
rect 26148 31816 26200 31822
rect 26148 31758 26200 31764
rect 26056 30932 26108 30938
rect 26056 30874 26108 30880
rect 25780 30388 25832 30394
rect 25780 30330 25832 30336
rect 25596 30252 25648 30258
rect 25596 30194 25648 30200
rect 25136 28960 25188 28966
rect 25136 28902 25188 28908
rect 25148 28694 25176 28902
rect 25332 28694 25360 30126
rect 25516 30110 25728 30138
rect 25504 29708 25556 29714
rect 25556 29668 25636 29696
rect 25504 29650 25556 29656
rect 25412 29504 25464 29510
rect 25412 29446 25464 29452
rect 25424 29238 25452 29446
rect 25412 29232 25464 29238
rect 25412 29174 25464 29180
rect 25504 28960 25556 28966
rect 25504 28902 25556 28908
rect 25136 28688 25188 28694
rect 25320 28688 25372 28694
rect 25136 28630 25188 28636
rect 25240 28636 25320 28642
rect 25240 28630 25372 28636
rect 25240 28614 25360 28630
rect 25136 28552 25188 28558
rect 25136 28494 25188 28500
rect 25148 27130 25176 28494
rect 25136 27124 25188 27130
rect 25136 27066 25188 27072
rect 25240 26926 25268 28614
rect 25320 28552 25372 28558
rect 25320 28494 25372 28500
rect 25332 28218 25360 28494
rect 25412 28484 25464 28490
rect 25412 28426 25464 28432
rect 25320 28212 25372 28218
rect 25320 28154 25372 28160
rect 25320 27872 25372 27878
rect 25320 27814 25372 27820
rect 25332 27470 25360 27814
rect 25320 27464 25372 27470
rect 25320 27406 25372 27412
rect 25424 27130 25452 28426
rect 25516 27878 25544 28902
rect 25608 28150 25636 29668
rect 25596 28144 25648 28150
rect 25596 28086 25648 28092
rect 25504 27872 25556 27878
rect 25504 27814 25556 27820
rect 25412 27124 25464 27130
rect 25412 27066 25464 27072
rect 25228 26920 25280 26926
rect 25228 26862 25280 26868
rect 25424 26382 25452 27066
rect 25608 27062 25636 28086
rect 25700 27674 25728 30110
rect 25792 29646 25820 30330
rect 26068 30326 26096 30874
rect 26148 30728 26200 30734
rect 26148 30670 26200 30676
rect 26056 30320 26108 30326
rect 26056 30262 26108 30268
rect 26160 30190 26188 30670
rect 26240 30252 26292 30258
rect 26240 30194 26292 30200
rect 26148 30184 26200 30190
rect 26148 30126 26200 30132
rect 26056 30048 26108 30054
rect 26056 29990 26108 29996
rect 25780 29640 25832 29646
rect 25780 29582 25832 29588
rect 25792 29170 25820 29582
rect 26068 29510 26096 29990
rect 26160 29850 26188 30126
rect 26148 29844 26200 29850
rect 26148 29786 26200 29792
rect 26056 29504 26108 29510
rect 26056 29446 26108 29452
rect 26068 29170 26096 29446
rect 25780 29164 25832 29170
rect 26056 29164 26108 29170
rect 25780 29106 25832 29112
rect 25976 29124 26056 29152
rect 25976 29016 26004 29124
rect 26056 29106 26108 29112
rect 26160 29102 26188 29786
rect 26252 29238 26280 30194
rect 26240 29232 26292 29238
rect 26240 29174 26292 29180
rect 26148 29096 26200 29102
rect 26148 29038 26200 29044
rect 26332 29096 26384 29102
rect 26332 29038 26384 29044
rect 25884 28988 26004 29016
rect 25884 28200 25912 28988
rect 26344 28422 26372 29038
rect 26332 28416 26384 28422
rect 26332 28358 26384 28364
rect 26344 28218 26372 28358
rect 26332 28212 26384 28218
rect 25884 28172 26004 28200
rect 25872 28076 25924 28082
rect 25872 28018 25924 28024
rect 25688 27668 25740 27674
rect 25688 27610 25740 27616
rect 25700 27470 25728 27610
rect 25884 27606 25912 28018
rect 25872 27600 25924 27606
rect 25872 27542 25924 27548
rect 25688 27464 25740 27470
rect 25688 27406 25740 27412
rect 25596 27056 25648 27062
rect 25596 26998 25648 27004
rect 25412 26376 25464 26382
rect 25412 26318 25464 26324
rect 25608 25498 25636 26998
rect 25700 25770 25728 27406
rect 25976 27334 26004 28172
rect 26332 28154 26384 28160
rect 26148 28144 26200 28150
rect 26148 28086 26200 28092
rect 26056 27940 26108 27946
rect 26056 27882 26108 27888
rect 26068 27470 26096 27882
rect 26056 27464 26108 27470
rect 26056 27406 26108 27412
rect 25964 27328 26016 27334
rect 25964 27270 26016 27276
rect 25976 26874 26004 27270
rect 26160 27130 26188 28086
rect 26608 27464 26660 27470
rect 26608 27406 26660 27412
rect 26148 27124 26200 27130
rect 26148 27066 26200 27072
rect 26240 26988 26292 26994
rect 26240 26930 26292 26936
rect 25884 26846 26004 26874
rect 26148 26920 26200 26926
rect 26148 26862 26200 26868
rect 25884 26450 25912 26846
rect 25964 26784 26016 26790
rect 25964 26726 26016 26732
rect 25976 26586 26004 26726
rect 25964 26580 26016 26586
rect 25964 26522 26016 26528
rect 26160 26450 26188 26862
rect 25872 26444 25924 26450
rect 25872 26386 25924 26392
rect 26148 26444 26200 26450
rect 26148 26386 26200 26392
rect 26056 26376 26108 26382
rect 26056 26318 26108 26324
rect 26068 25906 26096 26318
rect 26252 26042 26280 26930
rect 26424 26852 26476 26858
rect 26424 26794 26476 26800
rect 26436 26450 26464 26794
rect 26424 26444 26476 26450
rect 26424 26386 26476 26392
rect 26332 26376 26384 26382
rect 26332 26318 26384 26324
rect 26240 26036 26292 26042
rect 26240 25978 26292 25984
rect 26344 25906 26372 26318
rect 26056 25900 26108 25906
rect 26056 25842 26108 25848
rect 26332 25900 26384 25906
rect 26332 25842 26384 25848
rect 25688 25764 25740 25770
rect 25688 25706 25740 25712
rect 25596 25492 25648 25498
rect 25596 25434 25648 25440
rect 25700 24954 25728 25706
rect 26620 25362 26648 27406
rect 26608 25356 26660 25362
rect 26608 25298 26660 25304
rect 26332 25288 26384 25294
rect 26332 25230 26384 25236
rect 25688 24948 25740 24954
rect 25688 24890 25740 24896
rect 26344 24410 26372 25230
rect 26332 24404 26384 24410
rect 26332 24346 26384 24352
rect 24964 22066 25084 22094
rect 24584 2576 24636 2582
rect 24582 2544 24584 2553
rect 24636 2544 24638 2553
rect 23756 2508 23808 2514
rect 24582 2479 24638 2488
rect 23756 2450 23808 2456
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 22468 2032 22520 2038
rect 22468 1974 22520 1980
rect 23860 800 23888 2246
rect 24964 1902 24992 22066
rect 25780 2372 25832 2378
rect 25780 2314 25832 2320
rect 24952 1896 25004 1902
rect 24952 1838 25004 1844
rect 25792 800 25820 2314
rect 26804 1970 26832 38542
rect 26884 38344 26936 38350
rect 26884 38286 26936 38292
rect 26896 37194 26924 38286
rect 26884 37188 26936 37194
rect 26884 37130 26936 37136
rect 26884 36780 26936 36786
rect 26884 36722 26936 36728
rect 26896 36106 26924 36722
rect 26988 36650 27016 39442
rect 27172 38962 27200 39782
rect 27264 39302 27292 40004
rect 27344 39986 27396 39992
rect 27448 39982 27476 41686
rect 27908 41682 27936 41958
rect 27896 41676 27948 41682
rect 27896 41618 27948 41624
rect 27712 41608 27764 41614
rect 27712 41550 27764 41556
rect 27724 40662 27752 41550
rect 27712 40656 27764 40662
rect 27712 40598 27764 40604
rect 27528 40520 27580 40526
rect 27528 40462 27580 40468
rect 27540 40118 27568 40462
rect 28092 40186 28120 42774
rect 28184 42566 28212 44678
rect 28264 43648 28316 43654
rect 28264 43590 28316 43596
rect 28276 42906 28304 43590
rect 28460 43314 28488 45222
rect 28908 45008 28960 45014
rect 28908 44950 28960 44956
rect 28632 44464 28684 44470
rect 28632 44406 28684 44412
rect 28644 43858 28672 44406
rect 28632 43852 28684 43858
rect 28632 43794 28684 43800
rect 28920 43790 28948 44950
rect 29012 43994 29040 45222
rect 29000 43988 29052 43994
rect 29000 43930 29052 43936
rect 28908 43784 28960 43790
rect 28908 43726 28960 43732
rect 29012 43382 29040 43930
rect 29000 43376 29052 43382
rect 29000 43318 29052 43324
rect 28448 43308 28500 43314
rect 28448 43250 28500 43256
rect 28540 43240 28592 43246
rect 28540 43182 28592 43188
rect 28264 42900 28316 42906
rect 28264 42842 28316 42848
rect 28172 42560 28224 42566
rect 28172 42502 28224 42508
rect 28184 41274 28212 42502
rect 28552 42090 28580 43182
rect 28908 42628 28960 42634
rect 28908 42570 28960 42576
rect 28920 42362 28948 42570
rect 28908 42356 28960 42362
rect 28908 42298 28960 42304
rect 28920 42226 28948 42298
rect 28908 42220 28960 42226
rect 28908 42162 28960 42168
rect 28540 42084 28592 42090
rect 28540 42026 28592 42032
rect 28448 41812 28500 41818
rect 28448 41754 28500 41760
rect 28172 41268 28224 41274
rect 28172 41210 28224 41216
rect 28460 41002 28488 41754
rect 29000 41540 29052 41546
rect 29000 41482 29052 41488
rect 29012 41138 29040 41482
rect 29000 41132 29052 41138
rect 29000 41074 29052 41080
rect 28448 40996 28500 41002
rect 28448 40938 28500 40944
rect 28540 40928 28592 40934
rect 28540 40870 28592 40876
rect 28552 40662 28580 40870
rect 28906 40760 28962 40769
rect 28906 40695 28962 40704
rect 28540 40656 28592 40662
rect 28540 40598 28592 40604
rect 28920 40594 28948 40695
rect 28908 40588 28960 40594
rect 28908 40530 28960 40536
rect 28080 40180 28132 40186
rect 28080 40122 28132 40128
rect 27528 40112 27580 40118
rect 27528 40054 27580 40060
rect 27436 39976 27488 39982
rect 27436 39918 27488 39924
rect 27344 39908 27396 39914
rect 27344 39850 27396 39856
rect 27252 39296 27304 39302
rect 27252 39238 27304 39244
rect 27264 38962 27292 39238
rect 27160 38956 27212 38962
rect 27160 38898 27212 38904
rect 27252 38956 27304 38962
rect 27252 38898 27304 38904
rect 27264 38826 27292 38898
rect 27252 38820 27304 38826
rect 27252 38762 27304 38768
rect 27068 38276 27120 38282
rect 27068 38218 27120 38224
rect 27080 37874 27108 38218
rect 27160 38208 27212 38214
rect 27264 38196 27292 38762
rect 27356 38486 27384 39850
rect 27448 38962 27476 39918
rect 28092 39914 28120 40122
rect 28080 39908 28132 39914
rect 28080 39850 28132 39856
rect 27436 38956 27488 38962
rect 27436 38898 27488 38904
rect 27344 38480 27396 38486
rect 27344 38422 27396 38428
rect 27212 38168 27292 38196
rect 27160 38150 27212 38156
rect 27068 37868 27120 37874
rect 27068 37810 27120 37816
rect 27068 37392 27120 37398
rect 27068 37334 27120 37340
rect 27080 36786 27108 37334
rect 27172 37262 27200 38150
rect 27160 37256 27212 37262
rect 27160 37198 27212 37204
rect 27068 36780 27120 36786
rect 27068 36722 27120 36728
rect 27356 36718 27384 38422
rect 27448 38350 27476 38898
rect 27712 38548 27764 38554
rect 27712 38490 27764 38496
rect 27436 38344 27488 38350
rect 27436 38286 27488 38292
rect 27724 37262 27752 38490
rect 28356 37800 28408 37806
rect 28356 37742 28408 37748
rect 28368 37262 28396 37742
rect 27528 37256 27580 37262
rect 27528 37198 27580 37204
rect 27712 37256 27764 37262
rect 27712 37198 27764 37204
rect 28356 37256 28408 37262
rect 28356 37198 28408 37204
rect 28540 37256 28592 37262
rect 28540 37198 28592 37204
rect 27436 36780 27488 36786
rect 27436 36722 27488 36728
rect 27344 36712 27396 36718
rect 27344 36654 27396 36660
rect 26976 36644 27028 36650
rect 26976 36586 27028 36592
rect 26988 36242 27016 36586
rect 27160 36576 27212 36582
rect 27160 36518 27212 36524
rect 26976 36236 27028 36242
rect 26976 36178 27028 36184
rect 26884 36100 26936 36106
rect 26884 36042 26936 36048
rect 26896 35630 26924 36042
rect 26884 35624 26936 35630
rect 26884 35566 26936 35572
rect 26988 35154 27016 36178
rect 27068 35692 27120 35698
rect 27172 35680 27200 36518
rect 27120 35652 27200 35680
rect 27068 35634 27120 35640
rect 27068 35556 27120 35562
rect 27068 35498 27120 35504
rect 26976 35148 27028 35154
rect 26976 35090 27028 35096
rect 26884 34604 26936 34610
rect 26884 34546 26936 34552
rect 26896 34202 26924 34546
rect 26884 34196 26936 34202
rect 26884 34138 26936 34144
rect 26988 32910 27016 35090
rect 27080 33998 27108 35498
rect 27160 35080 27212 35086
rect 27160 35022 27212 35028
rect 27172 34746 27200 35022
rect 27160 34740 27212 34746
rect 27160 34682 27212 34688
rect 27068 33992 27120 33998
rect 27068 33934 27120 33940
rect 27172 33862 27200 34682
rect 27356 34474 27384 36654
rect 27448 35698 27476 36722
rect 27436 35692 27488 35698
rect 27436 35634 27488 35640
rect 27344 34468 27396 34474
rect 27344 34410 27396 34416
rect 27160 33856 27212 33862
rect 27160 33798 27212 33804
rect 27252 33856 27304 33862
rect 27252 33798 27304 33804
rect 27264 33522 27292 33798
rect 27252 33516 27304 33522
rect 27252 33458 27304 33464
rect 26976 32904 27028 32910
rect 26976 32846 27028 32852
rect 26988 31346 27016 32846
rect 27356 32570 27384 34410
rect 27436 34400 27488 34406
rect 27436 34342 27488 34348
rect 27448 33454 27476 34342
rect 27436 33448 27488 33454
rect 27436 33390 27488 33396
rect 27344 32564 27396 32570
rect 27344 32506 27396 32512
rect 27252 31952 27304 31958
rect 27252 31894 27304 31900
rect 27264 31346 27292 31894
rect 26976 31340 27028 31346
rect 26976 31282 27028 31288
rect 27252 31340 27304 31346
rect 27252 31282 27304 31288
rect 26988 30258 27016 31282
rect 27356 30938 27384 32506
rect 27344 30932 27396 30938
rect 27344 30874 27396 30880
rect 26976 30252 27028 30258
rect 26976 30194 27028 30200
rect 26988 29714 27016 30194
rect 26976 29708 27028 29714
rect 26976 29650 27028 29656
rect 27252 29640 27304 29646
rect 27252 29582 27304 29588
rect 26976 28960 27028 28966
rect 26976 28902 27028 28908
rect 26988 28558 27016 28902
rect 26976 28552 27028 28558
rect 26976 28494 27028 28500
rect 27264 27946 27292 29582
rect 27436 29028 27488 29034
rect 27436 28970 27488 28976
rect 27448 28082 27476 28970
rect 27436 28076 27488 28082
rect 27436 28018 27488 28024
rect 27252 27940 27304 27946
rect 27252 27882 27304 27888
rect 27344 26988 27396 26994
rect 27344 26930 27396 26936
rect 27160 26784 27212 26790
rect 27160 26726 27212 26732
rect 27172 26450 27200 26726
rect 27160 26444 27212 26450
rect 27160 26386 27212 26392
rect 27068 26376 27120 26382
rect 27068 26318 27120 26324
rect 27080 26042 27108 26318
rect 27068 26036 27120 26042
rect 27068 25978 27120 25984
rect 27172 25974 27200 26386
rect 27160 25968 27212 25974
rect 27160 25910 27212 25916
rect 27172 25498 27200 25910
rect 27356 25838 27384 26930
rect 27448 25906 27476 28018
rect 27436 25900 27488 25906
rect 27436 25842 27488 25848
rect 27344 25832 27396 25838
rect 27344 25774 27396 25780
rect 27160 25492 27212 25498
rect 27160 25434 27212 25440
rect 27356 25430 27384 25774
rect 27344 25424 27396 25430
rect 27344 25366 27396 25372
rect 27540 22094 27568 37198
rect 27724 36174 27752 37198
rect 27988 37120 28040 37126
rect 27988 37062 28040 37068
rect 27712 36168 27764 36174
rect 27712 36110 27764 36116
rect 27724 34950 27752 36110
rect 28000 35766 28028 37062
rect 28552 36378 28580 37198
rect 28920 37194 28948 40530
rect 28908 37188 28960 37194
rect 28908 37130 28960 37136
rect 28724 37120 28776 37126
rect 28724 37062 28776 37068
rect 28540 36372 28592 36378
rect 28540 36314 28592 36320
rect 28736 36242 28764 37062
rect 29184 36712 29236 36718
rect 29184 36654 29236 36660
rect 28724 36236 28776 36242
rect 28724 36178 28776 36184
rect 29000 36168 29052 36174
rect 29000 36110 29052 36116
rect 27988 35760 28040 35766
rect 27988 35702 28040 35708
rect 27712 34944 27764 34950
rect 27712 34886 27764 34892
rect 27724 32230 27752 34886
rect 27712 32224 27764 32230
rect 27712 32166 27764 32172
rect 27724 31754 27752 32166
rect 27712 31748 27764 31754
rect 27712 31690 27764 31696
rect 27724 30598 27752 31690
rect 28000 31210 28028 35702
rect 29012 35562 29040 36110
rect 29196 36038 29224 36654
rect 29184 36032 29236 36038
rect 29184 35974 29236 35980
rect 29000 35556 29052 35562
rect 29000 35498 29052 35504
rect 28356 35284 28408 35290
rect 28356 35226 28408 35232
rect 28172 34400 28224 34406
rect 28172 34342 28224 34348
rect 28184 33998 28212 34342
rect 28368 34066 28396 35226
rect 29092 35216 29144 35222
rect 29092 35158 29144 35164
rect 29104 34610 29132 35158
rect 29196 35154 29224 35974
rect 29184 35148 29236 35154
rect 29184 35090 29236 35096
rect 28816 34604 28868 34610
rect 28816 34546 28868 34552
rect 29092 34604 29144 34610
rect 29092 34546 29144 34552
rect 28828 34134 28856 34546
rect 29000 34536 29052 34542
rect 29000 34478 29052 34484
rect 29012 34134 29040 34478
rect 28816 34128 28868 34134
rect 28816 34070 28868 34076
rect 29000 34128 29052 34134
rect 29000 34070 29052 34076
rect 28264 34060 28316 34066
rect 28264 34002 28316 34008
rect 28356 34060 28408 34066
rect 28356 34002 28408 34008
rect 28172 33992 28224 33998
rect 28172 33934 28224 33940
rect 28276 33590 28304 34002
rect 28828 33998 28856 34070
rect 29092 34060 29144 34066
rect 29092 34002 29144 34008
rect 28816 33992 28868 33998
rect 28816 33934 28868 33940
rect 28264 33584 28316 33590
rect 28264 33526 28316 33532
rect 28276 33046 28304 33526
rect 29104 33522 29132 34002
rect 28724 33516 28776 33522
rect 28724 33458 28776 33464
rect 29092 33516 29144 33522
rect 29092 33458 29144 33464
rect 28736 33289 28764 33458
rect 29000 33380 29052 33386
rect 29000 33322 29052 33328
rect 28722 33280 28778 33289
rect 28722 33215 28778 33224
rect 28264 33040 28316 33046
rect 28264 32982 28316 32988
rect 28736 32910 28764 33215
rect 28724 32904 28776 32910
rect 28724 32846 28776 32852
rect 28736 32570 28764 32846
rect 28448 32564 28500 32570
rect 28448 32506 28500 32512
rect 28724 32564 28776 32570
rect 28724 32506 28776 32512
rect 28460 32298 28488 32506
rect 28908 32360 28960 32366
rect 28908 32302 28960 32308
rect 28448 32292 28500 32298
rect 28448 32234 28500 32240
rect 28920 31754 28948 32302
rect 29012 31958 29040 33322
rect 29104 33046 29132 33458
rect 29196 33386 29224 35090
rect 29276 34128 29328 34134
rect 29276 34070 29328 34076
rect 29288 33658 29316 34070
rect 29276 33652 29328 33658
rect 29276 33594 29328 33600
rect 29368 33448 29420 33454
rect 29366 33416 29368 33425
rect 29420 33416 29422 33425
rect 29184 33380 29236 33386
rect 29366 33351 29422 33360
rect 29184 33322 29236 33328
rect 29092 33040 29144 33046
rect 29092 32982 29144 32988
rect 29000 31952 29052 31958
rect 29000 31894 29052 31900
rect 28908 31748 28960 31754
rect 28908 31690 28960 31696
rect 28920 31346 28948 31690
rect 28908 31340 28960 31346
rect 28908 31282 28960 31288
rect 27988 31204 28040 31210
rect 27988 31146 28040 31152
rect 27712 30592 27764 30598
rect 27712 30534 27764 30540
rect 27620 29504 27672 29510
rect 27620 29446 27672 29452
rect 27632 27538 27660 29446
rect 27724 29034 27752 30534
rect 27804 29708 27856 29714
rect 27804 29650 27856 29656
rect 27816 29170 27844 29650
rect 27804 29164 27856 29170
rect 27804 29106 27856 29112
rect 27712 29028 27764 29034
rect 27712 28970 27764 28976
rect 27816 28626 27844 29106
rect 27804 28620 27856 28626
rect 27804 28562 27856 28568
rect 27804 28484 27856 28490
rect 27804 28426 27856 28432
rect 27816 28218 27844 28426
rect 27804 28212 27856 28218
rect 27804 28154 27856 28160
rect 27896 28008 27948 28014
rect 28000 27996 28028 31146
rect 28356 31136 28408 31142
rect 28356 31078 28408 31084
rect 28368 30734 28396 31078
rect 28356 30728 28408 30734
rect 28356 30670 28408 30676
rect 28080 28416 28132 28422
rect 28080 28358 28132 28364
rect 28092 28082 28120 28358
rect 28080 28076 28132 28082
rect 28080 28018 28132 28024
rect 27948 27968 28028 27996
rect 27896 27950 27948 27956
rect 27908 27674 27936 27950
rect 27896 27668 27948 27674
rect 27896 27610 27948 27616
rect 27620 27532 27672 27538
rect 27620 27474 27672 27480
rect 27620 27396 27672 27402
rect 27620 27338 27672 27344
rect 27632 27062 27660 27338
rect 27804 27328 27856 27334
rect 27804 27270 27856 27276
rect 27620 27056 27672 27062
rect 27620 26998 27672 27004
rect 27632 26586 27660 26998
rect 27620 26580 27672 26586
rect 27620 26522 27672 26528
rect 27816 26450 27844 27270
rect 27896 26988 27948 26994
rect 27896 26930 27948 26936
rect 27988 26988 28040 26994
rect 27988 26930 28040 26936
rect 27804 26444 27856 26450
rect 27804 26386 27856 26392
rect 27620 26308 27672 26314
rect 27620 26250 27672 26256
rect 27632 25838 27660 26250
rect 27908 26042 27936 26930
rect 28000 26042 28028 26930
rect 28092 26586 28120 28018
rect 28172 27464 28224 27470
rect 28172 27406 28224 27412
rect 28184 26858 28212 27406
rect 28264 26988 28316 26994
rect 28264 26930 28316 26936
rect 28172 26852 28224 26858
rect 28172 26794 28224 26800
rect 28080 26580 28132 26586
rect 28080 26522 28132 26528
rect 28276 26518 28304 26930
rect 28264 26512 28316 26518
rect 28264 26454 28316 26460
rect 27896 26036 27948 26042
rect 27896 25978 27948 25984
rect 27988 26036 28040 26042
rect 27988 25978 28040 25984
rect 27620 25832 27672 25838
rect 27620 25774 27672 25780
rect 27620 25220 27672 25226
rect 27620 25162 27672 25168
rect 27632 24614 27660 25162
rect 28276 25158 28304 26454
rect 28264 25152 28316 25158
rect 28264 25094 28316 25100
rect 28276 24818 28304 25094
rect 28264 24812 28316 24818
rect 28264 24754 28316 24760
rect 27620 24608 27672 24614
rect 27620 24550 27672 24556
rect 28080 24608 28132 24614
rect 28080 24550 28132 24556
rect 27632 24274 27660 24550
rect 27620 24268 27672 24274
rect 27620 24210 27672 24216
rect 27448 22066 27568 22094
rect 27448 11626 27476 22066
rect 28092 16574 28120 24550
rect 28092 16546 28212 16574
rect 27436 11620 27488 11626
rect 27436 11562 27488 11568
rect 28184 2650 28212 16546
rect 28172 2644 28224 2650
rect 28172 2586 28224 2592
rect 27712 2372 27764 2378
rect 27712 2314 27764 2320
rect 26792 1964 26844 1970
rect 26792 1906 26844 1912
rect 27724 800 27752 2314
rect 28368 2038 28396 30670
rect 28816 29640 28868 29646
rect 28816 29582 28868 29588
rect 28540 29164 28592 29170
rect 28540 29106 28592 29112
rect 28552 28762 28580 29106
rect 28724 28960 28776 28966
rect 28724 28902 28776 28908
rect 28540 28756 28592 28762
rect 28540 28698 28592 28704
rect 28448 28552 28500 28558
rect 28448 28494 28500 28500
rect 28460 27946 28488 28494
rect 28736 28150 28764 28902
rect 28828 28150 28856 29582
rect 29092 29504 29144 29510
rect 29092 29446 29144 29452
rect 29000 28552 29052 28558
rect 29000 28494 29052 28500
rect 28724 28144 28776 28150
rect 28724 28086 28776 28092
rect 28816 28144 28868 28150
rect 28816 28086 28868 28092
rect 28448 27940 28500 27946
rect 28448 27882 28500 27888
rect 28724 27872 28776 27878
rect 28724 27814 28776 27820
rect 28736 27470 28764 27814
rect 28828 27606 28856 28086
rect 29012 27606 29040 28494
rect 29104 28014 29132 29446
rect 29092 28008 29144 28014
rect 29092 27950 29144 27956
rect 28816 27600 28868 27606
rect 28816 27542 28868 27548
rect 29000 27600 29052 27606
rect 29000 27542 29052 27548
rect 29104 27470 29132 27950
rect 28724 27464 28776 27470
rect 28724 27406 28776 27412
rect 29092 27464 29144 27470
rect 29092 27406 29144 27412
rect 28632 27396 28684 27402
rect 28632 27338 28684 27344
rect 28644 27130 28672 27338
rect 28632 27124 28684 27130
rect 28632 27066 28684 27072
rect 29184 26920 29236 26926
rect 29184 26862 29236 26868
rect 29276 26920 29328 26926
rect 29276 26862 29328 26868
rect 29196 25838 29224 26862
rect 29288 26382 29316 26862
rect 29276 26376 29328 26382
rect 29276 26318 29328 26324
rect 29184 25832 29236 25838
rect 29184 25774 29236 25780
rect 29288 25498 29316 26318
rect 29368 25968 29420 25974
rect 29368 25910 29420 25916
rect 29276 25492 29328 25498
rect 29276 25434 29328 25440
rect 29380 25294 29408 25910
rect 29368 25288 29420 25294
rect 29368 25230 29420 25236
rect 29380 24954 29408 25230
rect 29368 24948 29420 24954
rect 29368 24890 29420 24896
rect 29380 23866 29408 24890
rect 29368 23860 29420 23866
rect 29368 23802 29420 23808
rect 29472 8906 29500 45834
rect 30024 44946 30052 49710
rect 30196 48748 30248 48754
rect 30196 48690 30248 48696
rect 30104 48340 30156 48346
rect 30104 48282 30156 48288
rect 30116 46578 30144 48282
rect 30208 48278 30236 48690
rect 30196 48272 30248 48278
rect 30196 48214 30248 48220
rect 30288 48136 30340 48142
rect 30288 48078 30340 48084
rect 30300 47258 30328 48078
rect 30288 47252 30340 47258
rect 30288 47194 30340 47200
rect 30196 47116 30248 47122
rect 30196 47058 30248 47064
rect 30208 46714 30236 47058
rect 30196 46708 30248 46714
rect 30196 46650 30248 46656
rect 30104 46572 30156 46578
rect 30104 46514 30156 46520
rect 30196 45960 30248 45966
rect 30196 45902 30248 45908
rect 30012 44940 30064 44946
rect 30012 44882 30064 44888
rect 30024 43874 30052 44882
rect 30024 43846 30144 43874
rect 30116 43790 30144 43846
rect 30104 43784 30156 43790
rect 30104 43726 30156 43732
rect 30116 43450 30144 43726
rect 30104 43444 30156 43450
rect 30104 43386 30156 43392
rect 30012 43376 30064 43382
rect 30012 43318 30064 43324
rect 29828 43104 29880 43110
rect 29828 43046 29880 43052
rect 29552 42764 29604 42770
rect 29552 42706 29604 42712
rect 29564 42514 29592 42706
rect 29644 42560 29696 42566
rect 29564 42508 29644 42514
rect 29564 42502 29696 42508
rect 29564 42486 29684 42502
rect 29564 42362 29592 42486
rect 29552 42356 29604 42362
rect 29552 42298 29604 42304
rect 29840 41449 29868 43046
rect 30024 42702 30052 43318
rect 30012 42696 30064 42702
rect 30012 42638 30064 42644
rect 29826 41440 29882 41449
rect 29826 41375 29882 41384
rect 29550 41304 29606 41313
rect 29550 41239 29606 41248
rect 29564 41138 29592 41239
rect 29552 41132 29604 41138
rect 29552 41074 29604 41080
rect 29840 41070 29868 41375
rect 29920 41200 29972 41206
rect 29920 41142 29972 41148
rect 29932 41070 29960 41142
rect 29828 41064 29880 41070
rect 29828 41006 29880 41012
rect 29920 41064 29972 41070
rect 29920 41006 29972 41012
rect 29736 40996 29788 41002
rect 29736 40938 29788 40944
rect 29644 40928 29696 40934
rect 29644 40870 29696 40876
rect 29550 39128 29606 39137
rect 29550 39063 29552 39072
rect 29604 39063 29606 39072
rect 29552 39034 29604 39040
rect 29656 37194 29684 40870
rect 29748 40118 29776 40938
rect 29828 40588 29880 40594
rect 29828 40530 29880 40536
rect 29736 40112 29788 40118
rect 29736 40054 29788 40060
rect 29748 37262 29776 40054
rect 29840 37398 29868 40530
rect 30012 39976 30064 39982
rect 30012 39918 30064 39924
rect 29920 39364 29972 39370
rect 29920 39306 29972 39312
rect 29932 39098 29960 39306
rect 29920 39092 29972 39098
rect 29920 39034 29972 39040
rect 30024 38554 30052 39918
rect 30012 38548 30064 38554
rect 30012 38490 30064 38496
rect 29920 38412 29972 38418
rect 29920 38354 29972 38360
rect 29932 37466 29960 38354
rect 30208 38298 30236 45902
rect 30380 45824 30432 45830
rect 30380 45766 30432 45772
rect 30392 45286 30420 45766
rect 30380 45280 30432 45286
rect 30380 45222 30432 45228
rect 30380 44396 30432 44402
rect 30380 44338 30432 44344
rect 30392 43314 30420 44338
rect 30380 43308 30432 43314
rect 30380 43250 30432 43256
rect 30392 41818 30420 43250
rect 30484 42838 30512 54606
rect 30748 54528 30800 54534
rect 30748 54470 30800 54476
rect 30564 54256 30616 54262
rect 30564 54198 30616 54204
rect 30576 53582 30604 54198
rect 30760 53990 30788 54470
rect 31392 54324 31444 54330
rect 31392 54266 31444 54272
rect 31208 54256 31260 54262
rect 31208 54198 31260 54204
rect 30748 53984 30800 53990
rect 30748 53926 30800 53932
rect 30760 53582 30788 53926
rect 30564 53576 30616 53582
rect 30564 53518 30616 53524
rect 30748 53576 30800 53582
rect 30748 53518 30800 53524
rect 30576 52494 30604 53518
rect 30564 52488 30616 52494
rect 30564 52430 30616 52436
rect 30760 52426 30788 53518
rect 30840 52964 30892 52970
rect 30840 52906 30892 52912
rect 30748 52420 30800 52426
rect 30748 52362 30800 52368
rect 30760 52306 30788 52362
rect 30668 52278 30788 52306
rect 30564 47660 30616 47666
rect 30564 47602 30616 47608
rect 30576 45014 30604 47602
rect 30668 46986 30696 52278
rect 30748 51808 30800 51814
rect 30748 51750 30800 51756
rect 30760 51474 30788 51750
rect 30748 51468 30800 51474
rect 30748 51410 30800 51416
rect 30760 50862 30788 51410
rect 30852 51406 30880 52906
rect 30840 51400 30892 51406
rect 30840 51342 30892 51348
rect 30852 50930 30880 51342
rect 30840 50924 30892 50930
rect 30840 50866 30892 50872
rect 30748 50856 30800 50862
rect 30748 50798 30800 50804
rect 30760 49638 30788 50798
rect 31024 50380 31076 50386
rect 31024 50322 31076 50328
rect 31036 50182 31064 50322
rect 31024 50176 31076 50182
rect 31024 50118 31076 50124
rect 31036 49910 31064 50118
rect 31024 49904 31076 49910
rect 31024 49846 31076 49852
rect 30748 49632 30800 49638
rect 30748 49574 30800 49580
rect 31116 49088 31168 49094
rect 31116 49030 31168 49036
rect 30840 48748 30892 48754
rect 30840 48690 30892 48696
rect 31024 48748 31076 48754
rect 31024 48690 31076 48696
rect 30852 47802 30880 48690
rect 30932 48544 30984 48550
rect 30932 48486 30984 48492
rect 30944 48142 30972 48486
rect 30932 48136 30984 48142
rect 30932 48078 30984 48084
rect 30840 47796 30892 47802
rect 30840 47738 30892 47744
rect 30852 47258 30880 47738
rect 31036 47666 31064 48690
rect 31128 48142 31156 49030
rect 31116 48136 31168 48142
rect 31116 48078 31168 48084
rect 31024 47660 31076 47666
rect 31024 47602 31076 47608
rect 31128 47598 31156 48078
rect 31116 47592 31168 47598
rect 31116 47534 31168 47540
rect 30840 47252 30892 47258
rect 30840 47194 30892 47200
rect 30748 47048 30800 47054
rect 30748 46990 30800 46996
rect 30930 47016 30986 47025
rect 30656 46980 30708 46986
rect 30656 46922 30708 46928
rect 30760 46714 30788 46990
rect 30930 46951 30932 46960
rect 30984 46951 30986 46960
rect 30932 46922 30984 46928
rect 30840 46912 30892 46918
rect 30840 46854 30892 46860
rect 30748 46708 30800 46714
rect 30748 46650 30800 46656
rect 30852 46578 30880 46854
rect 31220 46714 31248 54198
rect 31300 53780 31352 53786
rect 31300 53722 31352 53728
rect 31312 52154 31340 53722
rect 31404 53718 31432 54266
rect 31392 53712 31444 53718
rect 31392 53654 31444 53660
rect 31404 53242 31432 53654
rect 31392 53236 31444 53242
rect 31392 53178 31444 53184
rect 31484 53032 31536 53038
rect 31484 52974 31536 52980
rect 31300 52148 31352 52154
rect 31300 52090 31352 52096
rect 31496 51882 31524 52974
rect 31484 51876 31536 51882
rect 31484 51818 31536 51824
rect 31300 51400 31352 51406
rect 31300 51342 31352 51348
rect 31312 51066 31340 51342
rect 31392 51264 31444 51270
rect 31392 51206 31444 51212
rect 31300 51060 31352 51066
rect 31300 51002 31352 51008
rect 31312 50386 31340 51002
rect 31300 50380 31352 50386
rect 31300 50322 31352 50328
rect 31312 49842 31340 50322
rect 31404 50318 31432 51206
rect 31392 50312 31444 50318
rect 31392 50254 31444 50260
rect 31404 50182 31432 50254
rect 31392 50176 31444 50182
rect 31392 50118 31444 50124
rect 31300 49836 31352 49842
rect 31300 49778 31352 49784
rect 31300 48612 31352 48618
rect 31300 48554 31352 48560
rect 31312 47734 31340 48554
rect 31484 48544 31536 48550
rect 31484 48486 31536 48492
rect 31496 48346 31524 48486
rect 31484 48340 31536 48346
rect 31484 48282 31536 48288
rect 31300 47728 31352 47734
rect 31300 47670 31352 47676
rect 31312 47054 31340 47670
rect 31300 47048 31352 47054
rect 31300 46990 31352 46996
rect 31208 46708 31260 46714
rect 31208 46650 31260 46656
rect 30840 46572 30892 46578
rect 30840 46514 30892 46520
rect 30852 46034 30880 46514
rect 30932 46436 30984 46442
rect 30932 46378 30984 46384
rect 30840 46028 30892 46034
rect 30840 45970 30892 45976
rect 30944 45898 30972 46378
rect 30932 45892 30984 45898
rect 30932 45834 30984 45840
rect 30944 45082 30972 45834
rect 31220 45626 31248 46650
rect 31484 45824 31536 45830
rect 31484 45766 31536 45772
rect 31208 45620 31260 45626
rect 31208 45562 31260 45568
rect 30932 45076 30984 45082
rect 30932 45018 30984 45024
rect 30564 45008 30616 45014
rect 30564 44950 30616 44956
rect 30840 44736 30892 44742
rect 30840 44678 30892 44684
rect 30852 44538 30880 44678
rect 30840 44532 30892 44538
rect 30840 44474 30892 44480
rect 30944 44470 30972 45018
rect 30932 44464 30984 44470
rect 30984 44424 31064 44452
rect 30932 44406 30984 44412
rect 30932 43784 30984 43790
rect 30932 43726 30984 43732
rect 30748 43648 30800 43654
rect 30748 43590 30800 43596
rect 30472 42832 30524 42838
rect 30472 42774 30524 42780
rect 30564 42560 30616 42566
rect 30564 42502 30616 42508
rect 30576 42362 30604 42502
rect 30564 42356 30616 42362
rect 30564 42298 30616 42304
rect 30760 42294 30788 43590
rect 30840 43376 30892 43382
rect 30840 43318 30892 43324
rect 30852 42634 30880 43318
rect 30840 42628 30892 42634
rect 30840 42570 30892 42576
rect 30840 42356 30892 42362
rect 30840 42298 30892 42304
rect 30748 42288 30800 42294
rect 30748 42230 30800 42236
rect 30656 42220 30708 42226
rect 30656 42162 30708 42168
rect 30380 41812 30432 41818
rect 30380 41754 30432 41760
rect 30288 41540 30340 41546
rect 30288 41482 30340 41488
rect 30300 41138 30328 41482
rect 30288 41132 30340 41138
rect 30288 41074 30340 41080
rect 30288 38820 30340 38826
rect 30288 38762 30340 38768
rect 30024 38270 30236 38298
rect 29920 37460 29972 37466
rect 29920 37402 29972 37408
rect 29828 37392 29880 37398
rect 29828 37334 29880 37340
rect 29736 37256 29788 37262
rect 29736 37198 29788 37204
rect 29920 37256 29972 37262
rect 29920 37198 29972 37204
rect 29644 37188 29696 37194
rect 29644 37130 29696 37136
rect 29552 36848 29604 36854
rect 29552 36790 29604 36796
rect 29564 36174 29592 36790
rect 29656 36310 29684 37130
rect 29644 36304 29696 36310
rect 29644 36246 29696 36252
rect 29552 36168 29604 36174
rect 29552 36110 29604 36116
rect 29552 35624 29604 35630
rect 29552 35566 29604 35572
rect 29564 35494 29592 35566
rect 29552 35488 29604 35494
rect 29552 35430 29604 35436
rect 29564 34950 29592 35430
rect 29644 35012 29696 35018
rect 29644 34954 29696 34960
rect 29552 34944 29604 34950
rect 29552 34886 29604 34892
rect 29564 34066 29592 34886
rect 29552 34060 29604 34066
rect 29552 34002 29604 34008
rect 29656 33658 29684 34954
rect 29748 34134 29776 37198
rect 29932 36922 29960 37198
rect 29920 36916 29972 36922
rect 29920 36858 29972 36864
rect 29920 34536 29972 34542
rect 29920 34478 29972 34484
rect 29828 34468 29880 34474
rect 29828 34410 29880 34416
rect 29736 34128 29788 34134
rect 29736 34070 29788 34076
rect 29840 34066 29868 34410
rect 29932 34202 29960 34478
rect 29920 34196 29972 34202
rect 29920 34138 29972 34144
rect 29828 34060 29880 34066
rect 29828 34002 29880 34008
rect 29736 33992 29788 33998
rect 29736 33934 29788 33940
rect 29748 33658 29776 33934
rect 29644 33652 29696 33658
rect 29644 33594 29696 33600
rect 29736 33652 29788 33658
rect 29736 33594 29788 33600
rect 29920 33516 29972 33522
rect 29840 33476 29920 33504
rect 29840 33289 29868 33476
rect 29920 33458 29972 33464
rect 29920 33380 29972 33386
rect 29920 33322 29972 33328
rect 29826 33280 29882 33289
rect 29826 33215 29882 33224
rect 29932 32978 29960 33322
rect 29552 32972 29604 32978
rect 29552 32914 29604 32920
rect 29920 32972 29972 32978
rect 29920 32914 29972 32920
rect 29564 32434 29592 32914
rect 29644 32836 29696 32842
rect 29644 32778 29696 32784
rect 29656 32570 29684 32778
rect 29644 32564 29696 32570
rect 29644 32506 29696 32512
rect 29552 32428 29604 32434
rect 29552 32370 29604 32376
rect 29736 32428 29788 32434
rect 29736 32370 29788 32376
rect 29748 32230 29776 32370
rect 29736 32224 29788 32230
rect 29736 32166 29788 32172
rect 29932 31958 29960 32914
rect 29920 31952 29972 31958
rect 29920 31894 29972 31900
rect 30024 31754 30052 38270
rect 30104 38208 30156 38214
rect 30104 38150 30156 38156
rect 30116 37262 30144 38150
rect 30300 38010 30328 38762
rect 30288 38004 30340 38010
rect 30288 37946 30340 37952
rect 30104 37256 30156 37262
rect 30104 37198 30156 37204
rect 30104 36304 30156 36310
rect 30104 36246 30156 36252
rect 30116 34474 30144 36246
rect 30196 36100 30248 36106
rect 30196 36042 30248 36048
rect 30208 34542 30236 36042
rect 30300 35562 30328 37946
rect 30392 36854 30420 41754
rect 30668 41274 30696 42162
rect 30656 41268 30708 41274
rect 30656 41210 30708 41216
rect 30746 41032 30802 41041
rect 30746 40967 30802 40976
rect 30760 40526 30788 40967
rect 30852 40526 30880 42298
rect 30944 42226 30972 43726
rect 31036 42634 31064 44424
rect 31220 43450 31248 45562
rect 31300 44396 31352 44402
rect 31300 44338 31352 44344
rect 31312 44198 31340 44338
rect 31300 44192 31352 44198
rect 31300 44134 31352 44140
rect 31116 43444 31168 43450
rect 31116 43386 31168 43392
rect 31208 43444 31260 43450
rect 31208 43386 31260 43392
rect 31128 42906 31156 43386
rect 31312 43382 31340 44134
rect 31496 43654 31524 45766
rect 31588 44198 31616 56841
rect 34164 56794 34192 56841
rect 34256 56794 34284 56902
rect 34164 56766 34284 56794
rect 34440 55214 34468 56902
rect 36082 56841 36138 57641
rect 38658 56841 38714 57641
rect 40590 56841 40646 57641
rect 42522 56841 42578 57641
rect 45098 56841 45154 57641
rect 47030 56841 47086 57641
rect 48962 56841 49018 57641
rect 51538 56841 51594 57641
rect 53470 56841 53526 57641
rect 55402 56841 55458 57641
rect 34440 55186 34560 55214
rect 33876 54732 33928 54738
rect 33876 54674 33928 54680
rect 32680 54664 32732 54670
rect 32680 54606 32732 54612
rect 32404 54596 32456 54602
rect 32404 54538 32456 54544
rect 32416 54126 32444 54538
rect 32692 54194 32720 54606
rect 33048 54528 33100 54534
rect 33048 54470 33100 54476
rect 33060 54194 33088 54470
rect 32680 54188 32732 54194
rect 32680 54130 32732 54136
rect 33048 54188 33100 54194
rect 33048 54130 33100 54136
rect 33324 54188 33376 54194
rect 33324 54130 33376 54136
rect 31944 54120 31996 54126
rect 31944 54062 31996 54068
rect 32404 54120 32456 54126
rect 33336 54074 33364 54130
rect 32404 54062 32456 54068
rect 31668 53440 31720 53446
rect 31668 53382 31720 53388
rect 31680 53106 31708 53382
rect 31668 53100 31720 53106
rect 31668 53042 31720 53048
rect 31680 52698 31708 53042
rect 31668 52692 31720 52698
rect 31668 52634 31720 52640
rect 31760 52012 31812 52018
rect 31760 51954 31812 51960
rect 31772 51066 31800 51954
rect 31956 51270 31984 54062
rect 33244 54046 33364 54074
rect 33244 53990 33272 54046
rect 32220 53984 32272 53990
rect 32220 53926 32272 53932
rect 33232 53984 33284 53990
rect 33232 53926 33284 53932
rect 33416 53984 33468 53990
rect 33416 53926 33468 53932
rect 32128 53576 32180 53582
rect 32128 53518 32180 53524
rect 32036 53508 32088 53514
rect 32036 53450 32088 53456
rect 32048 53106 32076 53450
rect 32036 53100 32088 53106
rect 32036 53042 32088 53048
rect 32048 52562 32076 53042
rect 32036 52556 32088 52562
rect 32036 52498 32088 52504
rect 31944 51264 31996 51270
rect 31944 51206 31996 51212
rect 31760 51060 31812 51066
rect 31760 51002 31812 51008
rect 31772 49230 31800 51002
rect 31956 49366 31984 51206
rect 32140 49842 32168 53518
rect 32232 52902 32260 53926
rect 33428 53786 33456 53926
rect 33416 53780 33468 53786
rect 33416 53722 33468 53728
rect 33324 53712 33376 53718
rect 33324 53654 33376 53660
rect 32956 53508 33008 53514
rect 32956 53450 33008 53456
rect 32220 52896 32272 52902
rect 32220 52838 32272 52844
rect 32232 52086 32260 52838
rect 32220 52080 32272 52086
rect 32220 52022 32272 52028
rect 32588 51604 32640 51610
rect 32588 51546 32640 51552
rect 32600 51270 32628 51546
rect 32588 51264 32640 51270
rect 32588 51206 32640 51212
rect 32404 50924 32456 50930
rect 32404 50866 32456 50872
rect 32220 50720 32272 50726
rect 32220 50662 32272 50668
rect 32312 50720 32364 50726
rect 32312 50662 32364 50668
rect 32128 49836 32180 49842
rect 32128 49778 32180 49784
rect 31944 49360 31996 49366
rect 31944 49302 31996 49308
rect 32232 49230 32260 50662
rect 32324 50318 32352 50662
rect 32416 50522 32444 50866
rect 32496 50856 32548 50862
rect 32496 50798 32548 50804
rect 32404 50516 32456 50522
rect 32404 50458 32456 50464
rect 32508 50318 32536 50798
rect 32312 50312 32364 50318
rect 32312 50254 32364 50260
rect 32496 50312 32548 50318
rect 32496 50254 32548 50260
rect 32404 50176 32456 50182
rect 32404 50118 32456 50124
rect 32416 49230 32444 50118
rect 32508 49978 32536 50254
rect 32496 49972 32548 49978
rect 32496 49914 32548 49920
rect 32600 49858 32628 51206
rect 32508 49830 32628 49858
rect 32508 49298 32536 49830
rect 32588 49768 32640 49774
rect 32588 49710 32640 49716
rect 32600 49434 32628 49710
rect 32588 49428 32640 49434
rect 32588 49370 32640 49376
rect 32496 49292 32548 49298
rect 32496 49234 32548 49240
rect 32588 49292 32640 49298
rect 32588 49234 32640 49240
rect 31760 49224 31812 49230
rect 31760 49166 31812 49172
rect 32220 49224 32272 49230
rect 32220 49166 32272 49172
rect 32404 49224 32456 49230
rect 32404 49166 32456 49172
rect 31772 48006 31800 49166
rect 32508 49162 32536 49234
rect 32496 49156 32548 49162
rect 32496 49098 32548 49104
rect 32220 48272 32272 48278
rect 32220 48214 32272 48220
rect 31760 48000 31812 48006
rect 31760 47942 31812 47948
rect 31668 46980 31720 46986
rect 31668 46922 31720 46928
rect 31680 46442 31708 46922
rect 31772 46753 31800 47942
rect 32036 47660 32088 47666
rect 32036 47602 32088 47608
rect 32048 47569 32076 47602
rect 32034 47560 32090 47569
rect 32034 47495 32090 47504
rect 32048 47025 32076 47495
rect 32232 47054 32260 48214
rect 32404 48204 32456 48210
rect 32404 48146 32456 48152
rect 32416 47666 32444 48146
rect 32600 48142 32628 49234
rect 32680 49224 32732 49230
rect 32680 49166 32732 49172
rect 32588 48136 32640 48142
rect 32588 48078 32640 48084
rect 32600 47802 32628 48078
rect 32588 47796 32640 47802
rect 32588 47738 32640 47744
rect 32404 47660 32456 47666
rect 32404 47602 32456 47608
rect 32692 47258 32720 49166
rect 32680 47252 32732 47258
rect 32680 47194 32732 47200
rect 32496 47116 32548 47122
rect 32496 47058 32548 47064
rect 32220 47048 32272 47054
rect 32034 47016 32090 47025
rect 32272 47008 32352 47036
rect 32220 46990 32272 46996
rect 32034 46951 32090 46960
rect 31758 46744 31814 46753
rect 31758 46679 31814 46688
rect 32128 46572 32180 46578
rect 32128 46514 32180 46520
rect 31668 46436 31720 46442
rect 31668 46378 31720 46384
rect 32140 46102 32168 46514
rect 32220 46504 32272 46510
rect 32220 46446 32272 46452
rect 32128 46096 32180 46102
rect 32128 46038 32180 46044
rect 32140 45898 32168 46038
rect 32232 45898 32260 46446
rect 32128 45892 32180 45898
rect 32128 45834 32180 45840
rect 32220 45892 32272 45898
rect 32220 45834 32272 45840
rect 32140 45626 32168 45834
rect 32128 45620 32180 45626
rect 32128 45562 32180 45568
rect 32232 45490 32260 45834
rect 32220 45484 32272 45490
rect 32220 45426 32272 45432
rect 32324 44826 32352 47008
rect 32404 46368 32456 46374
rect 32404 46310 32456 46316
rect 32416 46170 32444 46310
rect 32508 46170 32536 47058
rect 32968 46646 32996 53450
rect 33336 53242 33364 53654
rect 33508 53440 33560 53446
rect 33508 53382 33560 53388
rect 33784 53440 33836 53446
rect 33784 53382 33836 53388
rect 33520 53242 33548 53382
rect 33324 53236 33376 53242
rect 33324 53178 33376 53184
rect 33508 53236 33560 53242
rect 33508 53178 33560 53184
rect 33508 53032 33560 53038
rect 33428 52980 33508 52986
rect 33428 52974 33560 52980
rect 33428 52958 33548 52974
rect 33428 52578 33456 52958
rect 33508 52896 33560 52902
rect 33508 52838 33560 52844
rect 33692 52896 33744 52902
rect 33692 52838 33744 52844
rect 33048 52556 33100 52562
rect 33152 52550 33456 52578
rect 33152 52544 33180 52550
rect 33100 52516 33180 52544
rect 33048 52498 33100 52504
rect 33324 52420 33376 52426
rect 33324 52362 33376 52368
rect 33336 52018 33364 52362
rect 33428 52154 33456 52550
rect 33416 52148 33468 52154
rect 33416 52090 33468 52096
rect 33324 52012 33376 52018
rect 33324 51954 33376 51960
rect 33140 51944 33192 51950
rect 33140 51886 33192 51892
rect 33152 51338 33180 51886
rect 33520 51406 33548 52838
rect 33600 52556 33652 52562
rect 33600 52498 33652 52504
rect 33612 51882 33640 52498
rect 33704 52358 33732 52838
rect 33692 52352 33744 52358
rect 33692 52294 33744 52300
rect 33704 52018 33732 52294
rect 33692 52012 33744 52018
rect 33692 51954 33744 51960
rect 33600 51876 33652 51882
rect 33600 51818 33652 51824
rect 33796 51406 33824 53382
rect 33888 52494 33916 54674
rect 34532 54602 34560 55186
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 36096 54874 36124 56841
rect 38672 54874 38700 56841
rect 40604 54874 40632 56841
rect 42536 55214 42564 56841
rect 42536 55186 42840 55214
rect 36084 54868 36136 54874
rect 36084 54810 36136 54816
rect 38660 54868 38712 54874
rect 38660 54810 38712 54816
rect 40592 54868 40644 54874
rect 40592 54810 40644 54816
rect 38672 54670 38700 54810
rect 42812 54670 42840 55186
rect 45112 54738 45140 56841
rect 47044 54874 47072 56841
rect 48976 54874 49004 56841
rect 51552 54874 51580 56841
rect 47032 54868 47084 54874
rect 47032 54810 47084 54816
rect 48964 54868 49016 54874
rect 48964 54810 49016 54816
rect 51540 54868 51592 54874
rect 51540 54810 51592 54816
rect 45100 54732 45152 54738
rect 45100 54674 45152 54680
rect 36084 54664 36136 54670
rect 36084 54606 36136 54612
rect 38660 54664 38712 54670
rect 38660 54606 38712 54612
rect 42800 54664 42852 54670
rect 42800 54606 42852 54612
rect 34520 54596 34572 54602
rect 34520 54538 34572 54544
rect 34532 54330 34560 54538
rect 34796 54528 34848 54534
rect 34796 54470 34848 54476
rect 34520 54324 34572 54330
rect 34520 54266 34572 54272
rect 34428 53780 34480 53786
rect 34428 53722 34480 53728
rect 34440 53242 34468 53722
rect 34520 53508 34572 53514
rect 34520 53450 34572 53456
rect 34152 53236 34204 53242
rect 34152 53178 34204 53184
rect 34428 53236 34480 53242
rect 34428 53178 34480 53184
rect 34164 52494 34192 53178
rect 34244 53100 34296 53106
rect 34244 53042 34296 53048
rect 34336 53100 34388 53106
rect 34336 53042 34388 53048
rect 34256 52698 34284 53042
rect 34244 52692 34296 52698
rect 34244 52634 34296 52640
rect 33876 52488 33928 52494
rect 33876 52430 33928 52436
rect 34152 52488 34204 52494
rect 34152 52430 34204 52436
rect 34164 52086 34192 52430
rect 34152 52080 34204 52086
rect 34152 52022 34204 52028
rect 33508 51400 33560 51406
rect 33508 51342 33560 51348
rect 33784 51400 33836 51406
rect 33784 51342 33836 51348
rect 34348 51338 34376 53042
rect 34532 53038 34560 53450
rect 34520 53032 34572 53038
rect 34520 52974 34572 52980
rect 34532 52018 34560 52974
rect 34612 52352 34664 52358
rect 34612 52294 34664 52300
rect 34520 52012 34572 52018
rect 34520 51954 34572 51960
rect 33140 51332 33192 51338
rect 33140 51274 33192 51280
rect 34336 51332 34388 51338
rect 34336 51274 34388 51280
rect 34532 50862 34560 51954
rect 34520 50856 34572 50862
rect 34520 50798 34572 50804
rect 33784 50720 33836 50726
rect 33784 50662 33836 50668
rect 33324 50448 33376 50454
rect 33324 50390 33376 50396
rect 33048 49768 33100 49774
rect 33048 49710 33100 49716
rect 33060 49366 33088 49710
rect 33048 49360 33100 49366
rect 33048 49302 33100 49308
rect 33232 49224 33284 49230
rect 33232 49166 33284 49172
rect 33244 48142 33272 49166
rect 33232 48136 33284 48142
rect 33232 48078 33284 48084
rect 33048 48068 33100 48074
rect 33048 48010 33100 48016
rect 33060 47666 33088 48010
rect 33140 48000 33192 48006
rect 33140 47942 33192 47948
rect 33048 47660 33100 47666
rect 33048 47602 33100 47608
rect 33152 47054 33180 47942
rect 33244 47666 33272 48078
rect 33232 47660 33284 47666
rect 33232 47602 33284 47608
rect 33232 47524 33284 47530
rect 33232 47466 33284 47472
rect 33244 47122 33272 47466
rect 33232 47116 33284 47122
rect 33336 47104 33364 50390
rect 33796 50318 33824 50662
rect 34624 50386 34652 52294
rect 34704 51400 34756 51406
rect 34704 51342 34756 51348
rect 34716 50862 34744 51342
rect 34704 50856 34756 50862
rect 34704 50798 34756 50804
rect 34612 50380 34664 50386
rect 34612 50322 34664 50328
rect 33784 50312 33836 50318
rect 33784 50254 33836 50260
rect 34152 50312 34204 50318
rect 34152 50254 34204 50260
rect 33796 49910 33824 50254
rect 34164 49978 34192 50254
rect 34336 50244 34388 50250
rect 34336 50186 34388 50192
rect 34152 49972 34204 49978
rect 34152 49914 34204 49920
rect 33784 49904 33836 49910
rect 33784 49846 33836 49852
rect 33796 49638 33824 49846
rect 33784 49632 33836 49638
rect 33784 49574 33836 49580
rect 33508 49224 33560 49230
rect 33508 49166 33560 49172
rect 33600 49224 33652 49230
rect 33600 49166 33652 49172
rect 33416 49088 33468 49094
rect 33416 49030 33468 49036
rect 33428 47666 33456 49030
rect 33520 48618 33548 49166
rect 33612 48890 33640 49166
rect 33600 48884 33652 48890
rect 33600 48826 33652 48832
rect 33796 48822 33824 49574
rect 33784 48816 33836 48822
rect 33784 48758 33836 48764
rect 33508 48612 33560 48618
rect 33508 48554 33560 48560
rect 33416 47660 33468 47666
rect 33416 47602 33468 47608
rect 33520 47598 33548 48554
rect 33600 48544 33652 48550
rect 33600 48486 33652 48492
rect 33508 47592 33560 47598
rect 33508 47534 33560 47540
rect 33612 47161 33640 48486
rect 33784 47728 33836 47734
rect 33784 47670 33836 47676
rect 33692 47456 33744 47462
rect 33692 47398 33744 47404
rect 33598 47152 33654 47161
rect 33336 47076 33456 47104
rect 33598 47087 33654 47096
rect 33232 47058 33284 47064
rect 33140 47048 33192 47054
rect 33140 46990 33192 46996
rect 33230 47016 33286 47025
rect 33230 46951 33232 46960
rect 33284 46951 33286 46960
rect 33324 46980 33376 46986
rect 33232 46922 33284 46928
rect 33324 46922 33376 46928
rect 33140 46912 33192 46918
rect 33140 46854 33192 46860
rect 32956 46640 33008 46646
rect 32956 46582 33008 46588
rect 32588 46572 32640 46578
rect 32588 46514 32640 46520
rect 32404 46164 32456 46170
rect 32404 46106 32456 46112
rect 32496 46164 32548 46170
rect 32496 46106 32548 46112
rect 32416 45558 32444 46106
rect 32404 45552 32456 45558
rect 32404 45494 32456 45500
rect 32600 45490 32628 46514
rect 33152 46510 33180 46854
rect 33336 46714 33364 46922
rect 33324 46708 33376 46714
rect 33324 46650 33376 46656
rect 33140 46504 33192 46510
rect 33140 46446 33192 46452
rect 33140 46164 33192 46170
rect 33140 46106 33192 46112
rect 32588 45484 32640 45490
rect 32588 45426 32640 45432
rect 32496 44872 32548 44878
rect 32324 44798 32444 44826
rect 32600 44860 32628 45426
rect 33152 45354 33180 46106
rect 33232 46028 33284 46034
rect 33232 45970 33284 45976
rect 33140 45348 33192 45354
rect 33140 45290 33192 45296
rect 33244 44928 33272 45970
rect 33428 45898 33456 47076
rect 33600 46572 33652 46578
rect 33520 46532 33600 46560
rect 33416 45892 33468 45898
rect 33416 45834 33468 45840
rect 33324 45824 33376 45830
rect 33324 45766 33376 45772
rect 33060 44900 33272 44928
rect 32548 44832 32628 44860
rect 32496 44814 32548 44820
rect 32312 44736 32364 44742
rect 32312 44678 32364 44684
rect 32324 44402 32352 44678
rect 32416 44470 32444 44798
rect 32404 44464 32456 44470
rect 32404 44406 32456 44412
rect 32312 44396 32364 44402
rect 32312 44338 32364 44344
rect 31576 44192 31628 44198
rect 31576 44134 31628 44140
rect 31484 43648 31536 43654
rect 31484 43590 31536 43596
rect 31300 43376 31352 43382
rect 31300 43318 31352 43324
rect 31392 43376 31444 43382
rect 31392 43318 31444 43324
rect 31208 43308 31260 43314
rect 31208 43250 31260 43256
rect 31116 42900 31168 42906
rect 31116 42842 31168 42848
rect 31024 42628 31076 42634
rect 31024 42570 31076 42576
rect 30932 42220 30984 42226
rect 30932 42162 30984 42168
rect 30944 41682 30972 42162
rect 30932 41676 30984 41682
rect 30932 41618 30984 41624
rect 30932 41132 30984 41138
rect 30932 41074 30984 41080
rect 30944 40730 30972 41074
rect 30932 40724 30984 40730
rect 30932 40666 30984 40672
rect 30748 40520 30800 40526
rect 30748 40462 30800 40468
rect 30840 40520 30892 40526
rect 30840 40462 30892 40468
rect 31024 40520 31076 40526
rect 31128 40508 31156 42842
rect 31220 42362 31248 43250
rect 31300 43240 31352 43246
rect 31300 43182 31352 43188
rect 31208 42356 31260 42362
rect 31208 42298 31260 42304
rect 31208 40928 31260 40934
rect 31208 40870 31260 40876
rect 31076 40480 31156 40508
rect 31024 40462 31076 40468
rect 30564 40384 30616 40390
rect 30564 40326 30616 40332
rect 30576 40050 30604 40326
rect 30564 40044 30616 40050
rect 30564 39986 30616 39992
rect 30576 38962 30604 39986
rect 30748 39976 30800 39982
rect 30748 39918 30800 39924
rect 30760 39438 30788 39918
rect 30840 39568 30892 39574
rect 30840 39510 30892 39516
rect 30748 39432 30800 39438
rect 30748 39374 30800 39380
rect 30656 39364 30708 39370
rect 30656 39306 30708 39312
rect 30564 38956 30616 38962
rect 30564 38898 30616 38904
rect 30472 38888 30524 38894
rect 30472 38830 30524 38836
rect 30484 37806 30512 38830
rect 30562 38448 30618 38457
rect 30562 38383 30618 38392
rect 30576 38214 30604 38383
rect 30564 38208 30616 38214
rect 30564 38150 30616 38156
rect 30472 37800 30524 37806
rect 30472 37742 30524 37748
rect 30668 37262 30696 39306
rect 30760 38457 30788 39374
rect 30852 39302 30880 39510
rect 31036 39386 31064 40462
rect 31220 40186 31248 40870
rect 31208 40180 31260 40186
rect 31208 40122 31260 40128
rect 31116 40044 31168 40050
rect 31116 39986 31168 39992
rect 31128 39506 31156 39986
rect 31116 39500 31168 39506
rect 31116 39442 31168 39448
rect 31036 39358 31156 39386
rect 30840 39296 30892 39302
rect 30840 39238 30892 39244
rect 31024 39296 31076 39302
rect 31024 39238 31076 39244
rect 30852 38486 30880 39238
rect 31036 38962 31064 39238
rect 30932 38956 30984 38962
rect 30932 38898 30984 38904
rect 31024 38956 31076 38962
rect 31024 38898 31076 38904
rect 30944 38554 30972 38898
rect 30932 38548 30984 38554
rect 30932 38490 30984 38496
rect 30840 38480 30892 38486
rect 30746 38448 30802 38457
rect 30840 38422 30892 38428
rect 30746 38383 30802 38392
rect 30852 38010 30880 38422
rect 30932 38208 30984 38214
rect 30932 38150 30984 38156
rect 30840 38004 30892 38010
rect 30840 37946 30892 37952
rect 30944 37330 30972 38150
rect 31024 37868 31076 37874
rect 31024 37810 31076 37816
rect 30932 37324 30984 37330
rect 30932 37266 30984 37272
rect 30656 37256 30708 37262
rect 30656 37198 30708 37204
rect 30748 37120 30800 37126
rect 30748 37062 30800 37068
rect 30380 36848 30432 36854
rect 30380 36790 30432 36796
rect 30392 35766 30420 36790
rect 30656 36576 30708 36582
rect 30656 36518 30708 36524
rect 30472 36168 30524 36174
rect 30472 36110 30524 36116
rect 30380 35760 30432 35766
rect 30380 35702 30432 35708
rect 30288 35556 30340 35562
rect 30288 35498 30340 35504
rect 30484 34678 30512 36110
rect 30668 36106 30696 36518
rect 30760 36174 30788 37062
rect 31036 36786 31064 37810
rect 31128 36854 31156 39358
rect 31208 38888 31260 38894
rect 31208 38830 31260 38836
rect 31220 38758 31248 38830
rect 31208 38752 31260 38758
rect 31208 38694 31260 38700
rect 31116 36848 31168 36854
rect 31116 36790 31168 36796
rect 30840 36780 30892 36786
rect 30840 36722 30892 36728
rect 31024 36780 31076 36786
rect 31024 36722 31076 36728
rect 30748 36168 30800 36174
rect 30748 36110 30800 36116
rect 30656 36100 30708 36106
rect 30656 36042 30708 36048
rect 30562 35048 30618 35057
rect 30562 34983 30618 34992
rect 30576 34950 30604 34983
rect 30564 34944 30616 34950
rect 30564 34886 30616 34892
rect 30472 34672 30524 34678
rect 30472 34614 30524 34620
rect 30288 34604 30340 34610
rect 30288 34546 30340 34552
rect 30196 34536 30248 34542
rect 30196 34478 30248 34484
rect 30104 34468 30156 34474
rect 30104 34410 30156 34416
rect 30116 33998 30144 34410
rect 30104 33992 30156 33998
rect 30104 33934 30156 33940
rect 30104 33448 30156 33454
rect 30102 33416 30104 33425
rect 30156 33416 30158 33425
rect 30102 33351 30158 33360
rect 30300 32774 30328 34546
rect 30380 33856 30432 33862
rect 30380 33798 30432 33804
rect 30472 33856 30524 33862
rect 30472 33798 30524 33804
rect 30392 32858 30420 33798
rect 30484 33590 30512 33798
rect 30472 33584 30524 33590
rect 30472 33526 30524 33532
rect 30392 32830 30512 32858
rect 30288 32768 30340 32774
rect 30288 32710 30340 32716
rect 30380 32768 30432 32774
rect 30380 32710 30432 32716
rect 30104 32496 30156 32502
rect 30102 32464 30104 32473
rect 30156 32464 30158 32473
rect 30102 32399 30158 32408
rect 30300 32212 30328 32710
rect 30392 32366 30420 32710
rect 30380 32360 30432 32366
rect 30380 32302 30432 32308
rect 30484 32298 30512 32830
rect 30472 32292 30524 32298
rect 30472 32234 30524 32240
rect 30300 32184 30420 32212
rect 30024 31726 30328 31754
rect 29552 31680 29604 31686
rect 29552 31622 29604 31628
rect 29564 31346 29592 31622
rect 29552 31340 29604 31346
rect 29552 31282 29604 31288
rect 29828 31136 29880 31142
rect 29828 31078 29880 31084
rect 29840 30734 29868 31078
rect 29828 30728 29880 30734
rect 29828 30670 29880 30676
rect 29828 29640 29880 29646
rect 29828 29582 29880 29588
rect 29840 29034 29868 29582
rect 29644 29028 29696 29034
rect 29644 28970 29696 28976
rect 29828 29028 29880 29034
rect 29828 28970 29880 28976
rect 29656 27606 29684 28970
rect 29828 28552 29880 28558
rect 29828 28494 29880 28500
rect 29840 28082 29868 28494
rect 29828 28076 29880 28082
rect 29828 28018 29880 28024
rect 29644 27600 29696 27606
rect 29644 27542 29696 27548
rect 29552 27532 29604 27538
rect 29552 27474 29604 27480
rect 29564 27130 29592 27474
rect 29552 27124 29604 27130
rect 29552 27066 29604 27072
rect 29656 26382 29684 27542
rect 29840 26858 29868 28018
rect 30012 27464 30064 27470
rect 30012 27406 30064 27412
rect 29828 26852 29880 26858
rect 29828 26794 29880 26800
rect 29644 26376 29696 26382
rect 30024 26364 30052 27406
rect 30104 26988 30156 26994
rect 30104 26930 30156 26936
rect 30116 26432 30144 26930
rect 30196 26784 30248 26790
rect 30196 26726 30248 26732
rect 30208 26586 30236 26726
rect 30196 26580 30248 26586
rect 30196 26522 30248 26528
rect 30196 26444 30248 26450
rect 30116 26404 30196 26432
rect 30196 26386 30248 26392
rect 30024 26336 30144 26364
rect 29644 26318 29696 26324
rect 29552 26240 29604 26246
rect 29552 26182 29604 26188
rect 29564 25906 29592 26182
rect 29656 25974 29684 26318
rect 29736 26308 29788 26314
rect 29736 26250 29788 26256
rect 29644 25968 29696 25974
rect 29644 25910 29696 25916
rect 29552 25900 29604 25906
rect 29552 25842 29604 25848
rect 29644 25832 29696 25838
rect 29644 25774 29696 25780
rect 29656 25498 29684 25774
rect 29644 25492 29696 25498
rect 29644 25434 29696 25440
rect 29748 25294 29776 26250
rect 30012 25900 30064 25906
rect 30012 25842 30064 25848
rect 30024 25362 30052 25842
rect 30012 25356 30064 25362
rect 30012 25298 30064 25304
rect 29736 25288 29788 25294
rect 29736 25230 29788 25236
rect 30024 24954 30052 25298
rect 30012 24948 30064 24954
rect 30012 24890 30064 24896
rect 30116 24274 30144 26336
rect 30208 26042 30236 26386
rect 30196 26036 30248 26042
rect 30196 25978 30248 25984
rect 30104 24268 30156 24274
rect 30104 24210 30156 24216
rect 30300 16658 30328 31726
rect 30392 31210 30420 32184
rect 30380 31204 30432 31210
rect 30380 31146 30432 31152
rect 30392 29510 30420 31146
rect 30380 29504 30432 29510
rect 30380 29446 30432 29452
rect 30392 28490 30420 29446
rect 30380 28484 30432 28490
rect 30380 28426 30432 28432
rect 30392 27946 30420 28426
rect 30380 27940 30432 27946
rect 30380 27882 30432 27888
rect 30380 27328 30432 27334
rect 30380 27270 30432 27276
rect 30392 27130 30420 27270
rect 30380 27124 30432 27130
rect 30380 27066 30432 27072
rect 30380 26920 30432 26926
rect 30380 26862 30432 26868
rect 30392 26382 30420 26862
rect 30380 26376 30432 26382
rect 30380 26318 30432 26324
rect 30392 24682 30420 26318
rect 30472 25696 30524 25702
rect 30472 25638 30524 25644
rect 30484 25362 30512 25638
rect 30472 25356 30524 25362
rect 30472 25298 30524 25304
rect 30472 25220 30524 25226
rect 30472 25162 30524 25168
rect 30484 24886 30512 25162
rect 30472 24880 30524 24886
rect 30472 24822 30524 24828
rect 30472 24744 30524 24750
rect 30472 24686 30524 24692
rect 30380 24676 30432 24682
rect 30380 24618 30432 24624
rect 30484 24410 30512 24686
rect 30472 24404 30524 24410
rect 30472 24346 30524 24352
rect 30288 16652 30340 16658
rect 30288 16594 30340 16600
rect 29460 8900 29512 8906
rect 29460 8842 29512 8848
rect 30576 2922 30604 34886
rect 30668 34610 30696 36042
rect 30748 35760 30800 35766
rect 30748 35702 30800 35708
rect 30760 34746 30788 35702
rect 30748 34740 30800 34746
rect 30748 34682 30800 34688
rect 30656 34604 30708 34610
rect 30656 34546 30708 34552
rect 30852 33318 30880 36722
rect 31116 36712 31168 36718
rect 31116 36654 31168 36660
rect 31128 36174 31156 36654
rect 31116 36168 31168 36174
rect 31116 36110 31168 36116
rect 31312 36020 31340 43182
rect 31404 42770 31432 43318
rect 31496 43314 31524 43590
rect 31484 43308 31536 43314
rect 31484 43250 31536 43256
rect 31392 42764 31444 42770
rect 31392 42706 31444 42712
rect 31404 40458 31432 42706
rect 31484 42356 31536 42362
rect 31484 42298 31536 42304
rect 31496 40662 31524 42298
rect 31588 41614 31616 44134
rect 32128 43308 32180 43314
rect 32128 43250 32180 43256
rect 32140 42906 32168 43250
rect 32416 43110 32444 44406
rect 32600 44402 32628 44832
rect 32772 44872 32824 44878
rect 32772 44814 32824 44820
rect 32588 44396 32640 44402
rect 32588 44338 32640 44344
rect 32600 43382 32628 44338
rect 32784 43994 32812 44814
rect 33060 44402 33088 44900
rect 33336 44810 33364 45766
rect 33520 45354 33548 46532
rect 33600 46514 33652 46520
rect 33600 45824 33652 45830
rect 33600 45766 33652 45772
rect 33612 45626 33640 45766
rect 33600 45620 33652 45626
rect 33600 45562 33652 45568
rect 33508 45348 33560 45354
rect 33508 45290 33560 45296
rect 33508 44872 33560 44878
rect 33508 44814 33560 44820
rect 33324 44804 33376 44810
rect 33324 44746 33376 44752
rect 33232 44736 33284 44742
rect 33232 44678 33284 44684
rect 33048 44396 33100 44402
rect 33048 44338 33100 44344
rect 33140 44328 33192 44334
rect 33140 44270 33192 44276
rect 32956 44260 33008 44266
rect 32956 44202 33008 44208
rect 32772 43988 32824 43994
rect 32772 43930 32824 43936
rect 32680 43716 32732 43722
rect 32680 43658 32732 43664
rect 32692 43450 32720 43658
rect 32680 43444 32732 43450
rect 32680 43386 32732 43392
rect 32588 43376 32640 43382
rect 32588 43318 32640 43324
rect 32404 43104 32456 43110
rect 32404 43046 32456 43052
rect 32128 42900 32180 42906
rect 32128 42842 32180 42848
rect 32128 42220 32180 42226
rect 32128 42162 32180 42168
rect 31576 41608 31628 41614
rect 31576 41550 31628 41556
rect 32140 41274 32168 42162
rect 32404 42016 32456 42022
rect 32404 41958 32456 41964
rect 32416 41614 32444 41958
rect 32404 41608 32456 41614
rect 32404 41550 32456 41556
rect 32220 41540 32272 41546
rect 32220 41482 32272 41488
rect 32128 41268 32180 41274
rect 32128 41210 32180 41216
rect 31484 40656 31536 40662
rect 31484 40598 31536 40604
rect 31392 40452 31444 40458
rect 31392 40394 31444 40400
rect 31576 40384 31628 40390
rect 31576 40326 31628 40332
rect 31760 40384 31812 40390
rect 31760 40326 31812 40332
rect 31484 39636 31536 39642
rect 31484 39578 31536 39584
rect 31392 39296 31444 39302
rect 31392 39238 31444 39244
rect 31404 39030 31432 39238
rect 31392 39024 31444 39030
rect 31392 38966 31444 38972
rect 31496 37262 31524 39578
rect 31588 39137 31616 40326
rect 31772 40050 31800 40326
rect 32232 40186 32260 41482
rect 32600 41313 32628 43318
rect 32586 41304 32642 41313
rect 32586 41239 32642 41248
rect 32600 41138 32628 41239
rect 32680 41200 32732 41206
rect 32680 41142 32732 41148
rect 32404 41132 32456 41138
rect 32404 41074 32456 41080
rect 32588 41132 32640 41138
rect 32588 41074 32640 41080
rect 32416 40730 32444 41074
rect 32404 40724 32456 40730
rect 32404 40666 32456 40672
rect 32220 40180 32272 40186
rect 32220 40122 32272 40128
rect 31760 40044 31812 40050
rect 31760 39986 31812 39992
rect 31668 39908 31720 39914
rect 31668 39850 31720 39856
rect 31574 39128 31630 39137
rect 31574 39063 31630 39072
rect 31588 39030 31616 39063
rect 31576 39024 31628 39030
rect 31576 38966 31628 38972
rect 31588 37874 31616 38966
rect 31576 37868 31628 37874
rect 31576 37810 31628 37816
rect 31680 37738 31708 39850
rect 31944 38344 31996 38350
rect 31944 38286 31996 38292
rect 32036 38344 32088 38350
rect 32036 38286 32088 38292
rect 31956 37806 31984 38286
rect 32048 37874 32076 38286
rect 32036 37868 32088 37874
rect 32036 37810 32088 37816
rect 31944 37800 31996 37806
rect 31944 37742 31996 37748
rect 31668 37732 31720 37738
rect 31668 37674 31720 37680
rect 31484 37256 31536 37262
rect 31484 37198 31536 37204
rect 31760 37256 31812 37262
rect 31760 37198 31812 37204
rect 31128 35992 31340 36020
rect 30932 35488 30984 35494
rect 30932 35430 30984 35436
rect 30840 33312 30892 33318
rect 30944 33289 30972 35430
rect 30840 33254 30892 33260
rect 30930 33280 30986 33289
rect 30748 33040 30800 33046
rect 30748 32982 30800 32988
rect 30656 30388 30708 30394
rect 30656 30330 30708 30336
rect 30668 28966 30696 30330
rect 30656 28960 30708 28966
rect 30656 28902 30708 28908
rect 30668 26518 30696 28902
rect 30760 28801 30788 32982
rect 30852 32910 30880 33254
rect 30930 33215 30986 33224
rect 30840 32904 30892 32910
rect 30840 32846 30892 32852
rect 30932 32768 30984 32774
rect 30932 32710 30984 32716
rect 30840 32496 30892 32502
rect 30838 32464 30840 32473
rect 30892 32464 30894 32473
rect 30838 32399 30894 32408
rect 30944 32230 30972 32710
rect 30932 32224 30984 32230
rect 30932 32166 30984 32172
rect 30944 31822 30972 32166
rect 30840 31816 30892 31822
rect 30840 31758 30892 31764
rect 30932 31816 30984 31822
rect 30932 31758 30984 31764
rect 30852 31210 30880 31758
rect 31024 31680 31076 31686
rect 31024 31622 31076 31628
rect 30840 31204 30892 31210
rect 30840 31146 30892 31152
rect 31036 30394 31064 31622
rect 31024 30388 31076 30394
rect 31024 30330 31076 30336
rect 30746 28792 30802 28801
rect 30746 28727 30802 28736
rect 30840 28416 30892 28422
rect 30840 28358 30892 28364
rect 30852 28082 30880 28358
rect 30840 28076 30892 28082
rect 30840 28018 30892 28024
rect 30932 28076 30984 28082
rect 30932 28018 30984 28024
rect 30852 27130 30880 28018
rect 30944 27946 30972 28018
rect 30932 27940 30984 27946
rect 30932 27882 30984 27888
rect 31024 27940 31076 27946
rect 31024 27882 31076 27888
rect 30944 27606 30972 27882
rect 30932 27600 30984 27606
rect 30932 27542 30984 27548
rect 31036 27402 31064 27882
rect 31024 27396 31076 27402
rect 31024 27338 31076 27344
rect 30840 27124 30892 27130
rect 30840 27066 30892 27072
rect 30656 26512 30708 26518
rect 30656 26454 30708 26460
rect 30748 25152 30800 25158
rect 30748 25094 30800 25100
rect 30760 24818 30788 25094
rect 30748 24812 30800 24818
rect 30748 24754 30800 24760
rect 30656 24064 30708 24070
rect 30656 24006 30708 24012
rect 30564 2916 30616 2922
rect 30564 2858 30616 2864
rect 30668 2514 30696 24006
rect 31128 2922 31156 35992
rect 31300 35284 31352 35290
rect 31300 35226 31352 35232
rect 31312 34610 31340 35226
rect 31392 34944 31444 34950
rect 31392 34886 31444 34892
rect 31404 34678 31432 34886
rect 31392 34672 31444 34678
rect 31392 34614 31444 34620
rect 31300 34604 31352 34610
rect 31300 34546 31352 34552
rect 31300 34400 31352 34406
rect 31300 34342 31352 34348
rect 31312 33998 31340 34342
rect 31392 34060 31444 34066
rect 31392 34002 31444 34008
rect 31300 33992 31352 33998
rect 31300 33934 31352 33940
rect 31208 32904 31260 32910
rect 31208 32846 31260 32852
rect 31220 32434 31248 32846
rect 31208 32428 31260 32434
rect 31208 32370 31260 32376
rect 31220 30938 31248 32370
rect 31208 30932 31260 30938
rect 31208 30874 31260 30880
rect 31220 29850 31248 30874
rect 31208 29844 31260 29850
rect 31208 29786 31260 29792
rect 31312 29170 31340 33934
rect 31404 33590 31432 34002
rect 31392 33584 31444 33590
rect 31392 33526 31444 33532
rect 31404 32978 31432 33526
rect 31392 32972 31444 32978
rect 31392 32914 31444 32920
rect 31404 32230 31432 32914
rect 31496 32570 31524 37198
rect 31772 36582 31800 37198
rect 31760 36576 31812 36582
rect 31760 36518 31812 36524
rect 31576 36032 31628 36038
rect 31576 35974 31628 35980
rect 31588 33862 31616 35974
rect 31772 35834 31800 36518
rect 31956 36106 31984 37742
rect 32128 37664 32180 37670
rect 32128 37606 32180 37612
rect 32140 37194 32168 37606
rect 32232 37262 32260 40122
rect 32600 39506 32628 41074
rect 32692 39642 32720 41142
rect 32968 40458 32996 44202
rect 33048 43852 33100 43858
rect 33048 43794 33100 43800
rect 33060 42702 33088 43794
rect 33152 43246 33180 44270
rect 33244 43790 33272 44678
rect 33520 44538 33548 44814
rect 33600 44804 33652 44810
rect 33600 44746 33652 44752
rect 33508 44532 33560 44538
rect 33508 44474 33560 44480
rect 33416 44260 33468 44266
rect 33416 44202 33468 44208
rect 33428 43994 33456 44202
rect 33416 43988 33468 43994
rect 33416 43930 33468 43936
rect 33612 43790 33640 44746
rect 33232 43784 33284 43790
rect 33232 43726 33284 43732
rect 33600 43784 33652 43790
rect 33600 43726 33652 43732
rect 33140 43240 33192 43246
rect 33140 43182 33192 43188
rect 33704 43178 33732 47398
rect 33796 47258 33824 47670
rect 33784 47252 33836 47258
rect 33784 47194 33836 47200
rect 33968 47048 34020 47054
rect 33968 46990 34020 46996
rect 33876 46504 33928 46510
rect 33876 46446 33928 46452
rect 33888 46034 33916 46446
rect 33876 46028 33928 46034
rect 33876 45970 33928 45976
rect 33874 45928 33930 45937
rect 33874 45863 33876 45872
rect 33928 45863 33930 45872
rect 33876 45834 33928 45840
rect 33888 45626 33916 45834
rect 33876 45620 33928 45626
rect 33876 45562 33928 45568
rect 33980 45082 34008 46990
rect 34060 46980 34112 46986
rect 34060 46922 34112 46928
rect 34072 46753 34100 46922
rect 34058 46744 34114 46753
rect 34058 46679 34060 46688
rect 34112 46679 34114 46688
rect 34060 46650 34112 46656
rect 34164 45966 34192 49914
rect 34348 49842 34376 50186
rect 34428 50176 34480 50182
rect 34428 50118 34480 50124
rect 34440 49910 34468 50118
rect 34624 49910 34652 50322
rect 34428 49904 34480 49910
rect 34428 49846 34480 49852
rect 34612 49904 34664 49910
rect 34612 49846 34664 49852
rect 34336 49836 34388 49842
rect 34336 49778 34388 49784
rect 34336 49156 34388 49162
rect 34336 49098 34388 49104
rect 34244 48816 34296 48822
rect 34244 48758 34296 48764
rect 34256 48074 34284 48758
rect 34244 48068 34296 48074
rect 34244 48010 34296 48016
rect 34256 46102 34284 48010
rect 34348 46866 34376 49098
rect 34612 49088 34664 49094
rect 34612 49030 34664 49036
rect 34624 48822 34652 49030
rect 34612 48816 34664 48822
rect 34612 48758 34664 48764
rect 34808 48634 34836 54470
rect 36096 53990 36124 54606
rect 38844 54528 38896 54534
rect 38844 54470 38896 54476
rect 40132 54528 40184 54534
rect 40132 54470 40184 54476
rect 42616 54528 42668 54534
rect 42616 54470 42668 54476
rect 36084 53984 36136 53990
rect 36084 53926 36136 53932
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 35624 52896 35676 52902
rect 35624 52838 35676 52844
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 35348 52692 35400 52698
rect 35348 52634 35400 52640
rect 35360 52154 35388 52634
rect 35348 52148 35400 52154
rect 35348 52090 35400 52096
rect 35532 52012 35584 52018
rect 35532 51954 35584 51960
rect 35348 51944 35400 51950
rect 35348 51886 35400 51892
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 34888 51332 34940 51338
rect 34888 51274 34940 51280
rect 34900 50930 34928 51274
rect 34888 50924 34940 50930
rect 34888 50866 34940 50872
rect 35360 50862 35388 51886
rect 35440 51808 35492 51814
rect 35440 51750 35492 51756
rect 35348 50856 35400 50862
rect 35348 50798 35400 50804
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 35360 50182 35388 50798
rect 35348 50176 35400 50182
rect 35348 50118 35400 50124
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 35256 49292 35308 49298
rect 35256 49234 35308 49240
rect 35268 48754 35296 49234
rect 35256 48748 35308 48754
rect 35256 48690 35308 48696
rect 34716 48606 34836 48634
rect 34428 48136 34480 48142
rect 34428 48078 34480 48084
rect 34440 47802 34468 48078
rect 34612 48000 34664 48006
rect 34612 47942 34664 47948
rect 34428 47796 34480 47802
rect 34428 47738 34480 47744
rect 34624 47598 34652 47942
rect 34612 47592 34664 47598
rect 34612 47534 34664 47540
rect 34612 46912 34664 46918
rect 34348 46860 34612 46866
rect 34348 46854 34664 46860
rect 34348 46838 34652 46854
rect 34244 46096 34296 46102
rect 34244 46038 34296 46044
rect 34152 45960 34204 45966
rect 34152 45902 34204 45908
rect 34348 45558 34376 46838
rect 34520 46096 34572 46102
rect 34520 46038 34572 46044
rect 34428 45824 34480 45830
rect 34428 45766 34480 45772
rect 34060 45552 34112 45558
rect 34060 45494 34112 45500
rect 34336 45552 34388 45558
rect 34336 45494 34388 45500
rect 33968 45076 34020 45082
rect 33968 45018 34020 45024
rect 34072 44146 34100 45494
rect 34336 45416 34388 45422
rect 34336 45358 34388 45364
rect 34348 44878 34376 45358
rect 34440 45014 34468 45766
rect 34532 45286 34560 46038
rect 34612 45960 34664 45966
rect 34610 45928 34612 45937
rect 34664 45928 34666 45937
rect 34610 45863 34666 45872
rect 34612 45824 34664 45830
rect 34612 45766 34664 45772
rect 34624 45490 34652 45766
rect 34612 45484 34664 45490
rect 34612 45426 34664 45432
rect 34716 45370 34744 48606
rect 34796 48544 34848 48550
rect 34796 48486 34848 48492
rect 34808 47666 34836 48486
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 35348 48204 35400 48210
rect 35348 48146 35400 48152
rect 35360 47666 35388 48146
rect 34796 47660 34848 47666
rect 34796 47602 34848 47608
rect 35348 47660 35400 47666
rect 35348 47602 35400 47608
rect 35346 47560 35402 47569
rect 35346 47495 35348 47504
rect 35400 47495 35402 47504
rect 35348 47466 35400 47472
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 35360 47190 35388 47466
rect 35348 47184 35400 47190
rect 35348 47126 35400 47132
rect 35452 46646 35480 51750
rect 35544 51610 35572 51954
rect 35636 51882 35664 52838
rect 35716 52420 35768 52426
rect 35716 52362 35768 52368
rect 35728 52154 35756 52362
rect 35900 52352 35952 52358
rect 35900 52294 35952 52300
rect 35716 52148 35768 52154
rect 35716 52090 35768 52096
rect 35624 51876 35676 51882
rect 35624 51818 35676 51824
rect 35532 51604 35584 51610
rect 35532 51546 35584 51552
rect 35636 51542 35664 51818
rect 35624 51536 35676 51542
rect 35624 51478 35676 51484
rect 35532 51264 35584 51270
rect 35636 51252 35664 51478
rect 35728 51406 35756 52090
rect 35912 51950 35940 52294
rect 35900 51944 35952 51950
rect 35900 51886 35952 51892
rect 35716 51400 35768 51406
rect 35716 51342 35768 51348
rect 35584 51224 35664 51252
rect 35532 51206 35584 51212
rect 35544 49638 35572 51206
rect 35728 51066 35756 51342
rect 35716 51060 35768 51066
rect 35716 51002 35768 51008
rect 35912 50930 35940 51886
rect 35900 50924 35952 50930
rect 35900 50866 35952 50872
rect 35912 50794 35940 50866
rect 35900 50788 35952 50794
rect 35900 50730 35952 50736
rect 35532 49632 35584 49638
rect 35532 49574 35584 49580
rect 35900 49632 35952 49638
rect 35900 49574 35952 49580
rect 35544 48686 35572 49574
rect 35912 49230 35940 49574
rect 35900 49224 35952 49230
rect 35900 49166 35952 49172
rect 35912 49094 35940 49166
rect 35900 49088 35952 49094
rect 35900 49030 35952 49036
rect 35532 48680 35584 48686
rect 35532 48622 35584 48628
rect 35544 48550 35572 48622
rect 35532 48544 35584 48550
rect 35532 48486 35584 48492
rect 35808 48544 35860 48550
rect 35808 48486 35860 48492
rect 35544 48074 35572 48486
rect 35820 48210 35848 48486
rect 35808 48204 35860 48210
rect 35808 48146 35860 48152
rect 35532 48068 35584 48074
rect 35532 48010 35584 48016
rect 35440 46640 35492 46646
rect 35440 46582 35492 46588
rect 34796 46572 34848 46578
rect 34796 46514 34848 46520
rect 34808 46374 34836 46514
rect 34796 46368 34848 46374
rect 34796 46310 34848 46316
rect 35348 46368 35400 46374
rect 35348 46310 35400 46316
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 34980 45960 35032 45966
rect 34980 45902 35032 45908
rect 34992 45626 35020 45902
rect 34980 45620 35032 45626
rect 34980 45562 35032 45568
rect 35360 45490 35388 46310
rect 35452 45966 35480 46582
rect 35440 45960 35492 45966
rect 35440 45902 35492 45908
rect 35348 45484 35400 45490
rect 35348 45426 35400 45432
rect 34624 45342 34744 45370
rect 34796 45416 34848 45422
rect 34796 45358 34848 45364
rect 34520 45280 34572 45286
rect 34520 45222 34572 45228
rect 34428 45008 34480 45014
rect 34428 44950 34480 44956
rect 34152 44872 34204 44878
rect 34152 44814 34204 44820
rect 34336 44872 34388 44878
rect 34336 44814 34388 44820
rect 34164 44266 34192 44814
rect 34440 44402 34468 44950
rect 34428 44396 34480 44402
rect 34428 44338 34480 44344
rect 34152 44260 34204 44266
rect 34152 44202 34204 44208
rect 34072 44118 34192 44146
rect 33784 43308 33836 43314
rect 33784 43250 33836 43256
rect 33692 43172 33744 43178
rect 33692 43114 33744 43120
rect 33232 43104 33284 43110
rect 33232 43046 33284 43052
rect 33048 42696 33100 42702
rect 33048 42638 33100 42644
rect 33244 42158 33272 43046
rect 33600 42764 33652 42770
rect 33600 42706 33652 42712
rect 33612 42566 33640 42706
rect 33692 42696 33744 42702
rect 33692 42638 33744 42644
rect 33600 42560 33652 42566
rect 33600 42502 33652 42508
rect 33232 42152 33284 42158
rect 33232 42094 33284 42100
rect 33600 42084 33652 42090
rect 33600 42026 33652 42032
rect 33612 41206 33640 42026
rect 33704 41818 33732 42638
rect 33796 42294 33824 43250
rect 33968 43240 34020 43246
rect 33968 43182 34020 43188
rect 33876 43172 33928 43178
rect 33876 43114 33928 43120
rect 33784 42288 33836 42294
rect 33784 42230 33836 42236
rect 33888 42090 33916 43114
rect 33980 42566 34008 43182
rect 34060 42832 34112 42838
rect 34060 42774 34112 42780
rect 33968 42560 34020 42566
rect 33968 42502 34020 42508
rect 34072 42226 34100 42774
rect 34060 42220 34112 42226
rect 34060 42162 34112 42168
rect 34164 42106 34192 44118
rect 34624 43466 34652 45342
rect 34704 45280 34756 45286
rect 34704 45222 34756 45228
rect 34532 43438 34652 43466
rect 34244 43308 34296 43314
rect 34244 43250 34296 43256
rect 34336 43308 34388 43314
rect 34336 43250 34388 43256
rect 34256 42702 34284 43250
rect 34348 42770 34376 43250
rect 34336 42764 34388 42770
rect 34336 42706 34388 42712
rect 34244 42696 34296 42702
rect 34244 42638 34296 42644
rect 34348 42548 34376 42706
rect 34348 42520 34468 42548
rect 33876 42084 33928 42090
rect 33876 42026 33928 42032
rect 33980 42078 34192 42106
rect 33692 41812 33744 41818
rect 33692 41754 33744 41760
rect 33980 41478 34008 42078
rect 34336 42016 34388 42022
rect 34336 41958 34388 41964
rect 34152 41812 34204 41818
rect 34152 41754 34204 41760
rect 34164 41614 34192 41754
rect 34152 41608 34204 41614
rect 34152 41550 34204 41556
rect 33876 41472 33928 41478
rect 33876 41414 33928 41420
rect 33968 41472 34020 41478
rect 33968 41414 34020 41420
rect 33600 41200 33652 41206
rect 33600 41142 33652 41148
rect 33784 41200 33836 41206
rect 33784 41142 33836 41148
rect 33416 41132 33468 41138
rect 33416 41074 33468 41080
rect 33232 40928 33284 40934
rect 33232 40870 33284 40876
rect 33244 40594 33272 40870
rect 33428 40662 33456 41074
rect 33796 40769 33824 41142
rect 33782 40760 33838 40769
rect 33782 40695 33838 40704
rect 33416 40656 33468 40662
rect 33416 40598 33468 40604
rect 33796 40594 33824 40695
rect 33232 40588 33284 40594
rect 33232 40530 33284 40536
rect 33784 40588 33836 40594
rect 33784 40530 33836 40536
rect 33416 40520 33468 40526
rect 33416 40462 33468 40468
rect 33508 40520 33560 40526
rect 33508 40462 33560 40468
rect 32956 40452 33008 40458
rect 32956 40394 33008 40400
rect 32968 40050 32996 40394
rect 32956 40044 33008 40050
rect 32956 39986 33008 39992
rect 33324 40044 33376 40050
rect 33324 39986 33376 39992
rect 32680 39636 32732 39642
rect 32680 39578 32732 39584
rect 32588 39500 32640 39506
rect 32588 39442 32640 39448
rect 32968 39370 32996 39986
rect 33232 39840 33284 39846
rect 33232 39782 33284 39788
rect 33140 39636 33192 39642
rect 33140 39578 33192 39584
rect 32956 39364 33008 39370
rect 32956 39306 33008 39312
rect 33048 39296 33100 39302
rect 33048 39238 33100 39244
rect 32956 38956 33008 38962
rect 32956 38898 33008 38904
rect 32496 38752 32548 38758
rect 32496 38694 32548 38700
rect 32508 37670 32536 38694
rect 32968 38554 32996 38898
rect 32956 38548 33008 38554
rect 32956 38490 33008 38496
rect 32588 38276 32640 38282
rect 32588 38218 32640 38224
rect 32600 37874 32628 38218
rect 33060 37874 33088 39238
rect 32588 37868 32640 37874
rect 32588 37810 32640 37816
rect 33048 37868 33100 37874
rect 33048 37810 33100 37816
rect 32496 37664 32548 37670
rect 32496 37606 32548 37612
rect 32404 37392 32456 37398
rect 32404 37334 32456 37340
rect 32220 37256 32272 37262
rect 32220 37198 32272 37204
rect 32128 37188 32180 37194
rect 32128 37130 32180 37136
rect 32036 36576 32088 36582
rect 32036 36518 32088 36524
rect 31944 36100 31996 36106
rect 31944 36042 31996 36048
rect 31852 36032 31904 36038
rect 31852 35974 31904 35980
rect 31760 35828 31812 35834
rect 31760 35770 31812 35776
rect 31864 35086 31892 35974
rect 32048 35698 32076 36518
rect 32140 35714 32168 37130
rect 32416 37126 32444 37334
rect 32600 37330 32628 37810
rect 32588 37324 32640 37330
rect 32588 37266 32640 37272
rect 32956 37188 33008 37194
rect 32956 37130 33008 37136
rect 32404 37120 32456 37126
rect 32404 37062 32456 37068
rect 32864 36168 32916 36174
rect 32864 36110 32916 36116
rect 32036 35692 32088 35698
rect 32140 35686 32260 35714
rect 32036 35634 32088 35640
rect 32128 35556 32180 35562
rect 32128 35498 32180 35504
rect 32140 35086 32168 35498
rect 31852 35080 31904 35086
rect 31852 35022 31904 35028
rect 32128 35080 32180 35086
rect 32128 35022 32180 35028
rect 31668 34944 31720 34950
rect 31668 34886 31720 34892
rect 31576 33856 31628 33862
rect 31576 33798 31628 33804
rect 31588 32910 31616 33798
rect 31680 32978 31708 34886
rect 31668 32972 31720 32978
rect 31668 32914 31720 32920
rect 31576 32904 31628 32910
rect 31576 32846 31628 32852
rect 31484 32564 31536 32570
rect 31484 32506 31536 32512
rect 31680 32434 31708 32914
rect 31944 32836 31996 32842
rect 31944 32778 31996 32784
rect 31668 32428 31720 32434
rect 31588 32388 31668 32416
rect 31392 32224 31444 32230
rect 31392 32166 31444 32172
rect 31484 32224 31536 32230
rect 31484 32166 31536 32172
rect 31392 32020 31444 32026
rect 31392 31962 31444 31968
rect 31404 31686 31432 31962
rect 31496 31822 31524 32166
rect 31484 31816 31536 31822
rect 31484 31758 31536 31764
rect 31392 31680 31444 31686
rect 31392 31622 31444 31628
rect 31484 29708 31536 29714
rect 31484 29650 31536 29656
rect 31392 29504 31444 29510
rect 31392 29446 31444 29452
rect 31300 29164 31352 29170
rect 31300 29106 31352 29112
rect 31300 29028 31352 29034
rect 31300 28970 31352 28976
rect 31312 28150 31340 28970
rect 31404 28422 31432 29446
rect 31392 28416 31444 28422
rect 31392 28358 31444 28364
rect 31300 28144 31352 28150
rect 31300 28086 31352 28092
rect 31300 27668 31352 27674
rect 31300 27610 31352 27616
rect 31312 26586 31340 27610
rect 31496 27606 31524 29650
rect 31588 29238 31616 32388
rect 31668 32370 31720 32376
rect 31956 32366 31984 32778
rect 31944 32360 31996 32366
rect 31996 32308 32076 32314
rect 31944 32302 32076 32308
rect 31956 32286 32076 32302
rect 31668 32224 31720 32230
rect 31668 32166 31720 32172
rect 31680 32026 31708 32166
rect 31668 32020 31720 32026
rect 31668 31962 31720 31968
rect 31760 31816 31812 31822
rect 31760 31758 31812 31764
rect 31772 31210 31800 31758
rect 31852 31272 31904 31278
rect 31852 31214 31904 31220
rect 31760 31204 31812 31210
rect 31760 31146 31812 31152
rect 31864 30734 31892 31214
rect 31944 31204 31996 31210
rect 31944 31146 31996 31152
rect 31956 30938 31984 31146
rect 31944 30932 31996 30938
rect 31944 30874 31996 30880
rect 31852 30728 31904 30734
rect 31852 30670 31904 30676
rect 31668 29776 31720 29782
rect 31668 29718 31720 29724
rect 31680 29646 31708 29718
rect 31668 29640 31720 29646
rect 31668 29582 31720 29588
rect 31852 29640 31904 29646
rect 31852 29582 31904 29588
rect 31576 29232 31628 29238
rect 31576 29174 31628 29180
rect 31588 28506 31616 29174
rect 31588 28478 31708 28506
rect 31576 28416 31628 28422
rect 31576 28358 31628 28364
rect 31588 28082 31616 28358
rect 31576 28076 31628 28082
rect 31576 28018 31628 28024
rect 31484 27600 31536 27606
rect 31484 27542 31536 27548
rect 31588 27538 31616 28018
rect 31680 27946 31708 28478
rect 31864 28218 31892 29582
rect 32048 29170 32076 32286
rect 32140 30802 32168 35022
rect 32232 32434 32260 35686
rect 32404 35556 32456 35562
rect 32404 35498 32456 35504
rect 32416 34746 32444 35498
rect 32680 35488 32732 35494
rect 32680 35430 32732 35436
rect 32692 35086 32720 35430
rect 32680 35080 32732 35086
rect 32680 35022 32732 35028
rect 32404 34740 32456 34746
rect 32404 34682 32456 34688
rect 32876 34610 32904 36110
rect 32404 34604 32456 34610
rect 32404 34546 32456 34552
rect 32588 34604 32640 34610
rect 32588 34546 32640 34552
rect 32864 34604 32916 34610
rect 32864 34546 32916 34552
rect 32416 34406 32444 34546
rect 32404 34400 32456 34406
rect 32404 34342 32456 34348
rect 32416 33318 32444 34342
rect 32600 34202 32628 34546
rect 32588 34196 32640 34202
rect 32588 34138 32640 34144
rect 32680 34196 32732 34202
rect 32680 34138 32732 34144
rect 32588 33856 32640 33862
rect 32588 33798 32640 33804
rect 32600 33454 32628 33798
rect 32692 33658 32720 34138
rect 32772 33992 32824 33998
rect 32772 33934 32824 33940
rect 32680 33652 32732 33658
rect 32680 33594 32732 33600
rect 32784 33538 32812 33934
rect 32876 33862 32904 34546
rect 32864 33856 32916 33862
rect 32864 33798 32916 33804
rect 32784 33510 32904 33538
rect 32876 33454 32904 33510
rect 32496 33448 32548 33454
rect 32496 33390 32548 33396
rect 32588 33448 32640 33454
rect 32588 33390 32640 33396
rect 32864 33448 32916 33454
rect 32864 33390 32916 33396
rect 32404 33312 32456 33318
rect 32508 33289 32536 33390
rect 32404 33254 32456 33260
rect 32494 33280 32550 33289
rect 32494 33215 32550 33224
rect 32508 32978 32536 33215
rect 32496 32972 32548 32978
rect 32496 32914 32548 32920
rect 32876 32842 32904 33390
rect 32864 32836 32916 32842
rect 32864 32778 32916 32784
rect 32968 32552 32996 37130
rect 33060 36310 33088 37810
rect 33152 37738 33180 39578
rect 33244 37874 33272 39782
rect 33336 39642 33364 39986
rect 33324 39636 33376 39642
rect 33324 39578 33376 39584
rect 33324 39500 33376 39506
rect 33324 39442 33376 39448
rect 33336 38654 33364 39442
rect 33428 39438 33456 40462
rect 33520 40186 33548 40462
rect 33888 40458 33916 41414
rect 34164 41138 34192 41550
rect 34244 41540 34296 41546
rect 34244 41482 34296 41488
rect 34152 41132 34204 41138
rect 34152 41074 34204 41080
rect 34164 40594 34192 41074
rect 34256 41070 34284 41482
rect 34244 41064 34296 41070
rect 34244 41006 34296 41012
rect 34152 40588 34204 40594
rect 34152 40530 34204 40536
rect 33876 40452 33928 40458
rect 33876 40394 33928 40400
rect 33508 40180 33560 40186
rect 33508 40122 33560 40128
rect 34164 40118 34192 40530
rect 34152 40112 34204 40118
rect 34152 40054 34204 40060
rect 34164 39982 34192 40054
rect 33508 39976 33560 39982
rect 33508 39918 33560 39924
rect 34152 39976 34204 39982
rect 34152 39918 34204 39924
rect 33416 39432 33468 39438
rect 33416 39374 33468 39380
rect 33520 39370 33548 39918
rect 33784 39636 33836 39642
rect 33784 39578 33836 39584
rect 34152 39636 34204 39642
rect 34152 39578 34204 39584
rect 33508 39364 33560 39370
rect 33508 39306 33560 39312
rect 33796 39302 33824 39578
rect 33784 39296 33836 39302
rect 33784 39238 33836 39244
rect 33416 38888 33468 38894
rect 33416 38830 33468 38836
rect 33428 38758 33456 38830
rect 33796 38758 33824 39238
rect 34164 38962 34192 39578
rect 34152 38956 34204 38962
rect 34152 38898 34204 38904
rect 33416 38752 33468 38758
rect 33416 38694 33468 38700
rect 33784 38752 33836 38758
rect 33784 38694 33836 38700
rect 34060 38752 34112 38758
rect 34060 38694 34112 38700
rect 33336 38626 33456 38654
rect 33428 38350 33456 38626
rect 33416 38344 33468 38350
rect 33414 38312 33416 38321
rect 33600 38344 33652 38350
rect 33468 38312 33470 38321
rect 33470 38270 33548 38298
rect 33600 38286 33652 38292
rect 33692 38344 33744 38350
rect 33692 38286 33744 38292
rect 33414 38247 33470 38256
rect 33416 38208 33468 38214
rect 33416 38150 33468 38156
rect 33428 38010 33456 38150
rect 33416 38004 33468 38010
rect 33416 37946 33468 37952
rect 33232 37868 33284 37874
rect 33232 37810 33284 37816
rect 33140 37732 33192 37738
rect 33140 37674 33192 37680
rect 33520 37466 33548 38270
rect 33612 38010 33640 38286
rect 33600 38004 33652 38010
rect 33600 37946 33652 37952
rect 33600 37664 33652 37670
rect 33600 37606 33652 37612
rect 33508 37460 33560 37466
rect 33508 37402 33560 37408
rect 33416 37188 33468 37194
rect 33416 37130 33468 37136
rect 33428 36786 33456 37130
rect 33416 36780 33468 36786
rect 33416 36722 33468 36728
rect 33520 36650 33548 37402
rect 33140 36644 33192 36650
rect 33140 36586 33192 36592
rect 33508 36644 33560 36650
rect 33508 36586 33560 36592
rect 33048 36304 33100 36310
rect 33048 36246 33100 36252
rect 33060 34678 33088 36246
rect 33048 34672 33100 34678
rect 33048 34614 33100 34620
rect 33060 33590 33088 34614
rect 33048 33584 33100 33590
rect 33048 33526 33100 33532
rect 33152 32570 33180 36586
rect 33324 36576 33376 36582
rect 33612 36530 33640 37606
rect 33704 36718 33732 38286
rect 33796 36854 33824 38694
rect 34072 38282 34100 38694
rect 34060 38276 34112 38282
rect 34060 38218 34112 38224
rect 33968 37868 34020 37874
rect 33968 37810 34020 37816
rect 33876 37120 33928 37126
rect 33876 37062 33928 37068
rect 33784 36848 33836 36854
rect 33784 36790 33836 36796
rect 33692 36712 33744 36718
rect 33692 36654 33744 36660
rect 33784 36644 33836 36650
rect 33784 36586 33836 36592
rect 33324 36518 33376 36524
rect 33232 35488 33284 35494
rect 33232 35430 33284 35436
rect 33244 34950 33272 35430
rect 33232 34944 33284 34950
rect 33232 34886 33284 34892
rect 33232 34400 33284 34406
rect 33232 34342 33284 34348
rect 33244 33998 33272 34342
rect 33232 33992 33284 33998
rect 33232 33934 33284 33940
rect 33336 33844 33364 36518
rect 33520 36502 33640 36530
rect 33520 36174 33548 36502
rect 33692 36372 33744 36378
rect 33692 36314 33744 36320
rect 33508 36168 33560 36174
rect 33508 36110 33560 36116
rect 33416 35216 33468 35222
rect 33416 35158 33468 35164
rect 33428 34406 33456 35158
rect 33416 34400 33468 34406
rect 33416 34342 33468 34348
rect 33244 33816 33364 33844
rect 33140 32564 33192 32570
rect 32968 32524 33088 32552
rect 32220 32428 32272 32434
rect 32220 32370 32272 32376
rect 32680 32428 32732 32434
rect 32680 32370 32732 32376
rect 32864 32428 32916 32434
rect 32864 32370 32916 32376
rect 32956 32428 33008 32434
rect 33060 32416 33088 32524
rect 33140 32506 33192 32512
rect 33060 32388 33180 32416
rect 32956 32370 33008 32376
rect 32232 31804 32260 32370
rect 32496 32292 32548 32298
rect 32496 32234 32548 32240
rect 32312 31816 32364 31822
rect 32232 31776 32312 31804
rect 32312 31758 32364 31764
rect 32508 31346 32536 32234
rect 32692 31890 32720 32370
rect 32680 31884 32732 31890
rect 32680 31826 32732 31832
rect 32680 31680 32732 31686
rect 32680 31622 32732 31628
rect 32220 31340 32272 31346
rect 32220 31282 32272 31288
rect 32496 31340 32548 31346
rect 32496 31282 32548 31288
rect 32232 30938 32260 31282
rect 32496 31136 32548 31142
rect 32496 31078 32548 31084
rect 32220 30932 32272 30938
rect 32220 30874 32272 30880
rect 32128 30796 32180 30802
rect 32128 30738 32180 30744
rect 32140 30190 32168 30738
rect 32508 30326 32536 31078
rect 32496 30320 32548 30326
rect 32496 30262 32548 30268
rect 32128 30184 32180 30190
rect 32128 30126 32180 30132
rect 32496 30048 32548 30054
rect 32496 29990 32548 29996
rect 32404 29504 32456 29510
rect 32404 29446 32456 29452
rect 32036 29164 32088 29170
rect 32036 29106 32088 29112
rect 31944 28960 31996 28966
rect 31944 28902 31996 28908
rect 31852 28212 31904 28218
rect 31852 28154 31904 28160
rect 31668 27940 31720 27946
rect 31668 27882 31720 27888
rect 31576 27532 31628 27538
rect 31576 27474 31628 27480
rect 31484 27396 31536 27402
rect 31484 27338 31536 27344
rect 31496 26994 31524 27338
rect 31484 26988 31536 26994
rect 31484 26930 31536 26936
rect 31680 26586 31708 27882
rect 31956 27538 31984 28902
rect 32048 28014 32076 29106
rect 32312 28756 32364 28762
rect 32312 28698 32364 28704
rect 32128 28144 32180 28150
rect 32128 28086 32180 28092
rect 32036 28008 32088 28014
rect 32036 27950 32088 27956
rect 31944 27532 31996 27538
rect 31944 27474 31996 27480
rect 32140 27470 32168 28086
rect 32324 28082 32352 28698
rect 32416 28558 32444 29446
rect 32508 28626 32536 29990
rect 32588 29640 32640 29646
rect 32588 29582 32640 29588
rect 32600 29170 32628 29582
rect 32588 29164 32640 29170
rect 32588 29106 32640 29112
rect 32600 28762 32628 29106
rect 32588 28756 32640 28762
rect 32588 28698 32640 28704
rect 32496 28620 32548 28626
rect 32496 28562 32548 28568
rect 32404 28552 32456 28558
rect 32404 28494 32456 28500
rect 32692 28082 32720 31622
rect 32772 31272 32824 31278
rect 32772 31214 32824 31220
rect 32784 30938 32812 31214
rect 32772 30932 32824 30938
rect 32772 30874 32824 30880
rect 32876 30666 32904 32370
rect 32968 31754 32996 32370
rect 33048 32292 33100 32298
rect 33048 32234 33100 32240
rect 33060 31822 33088 32234
rect 33152 31958 33180 32388
rect 33140 31952 33192 31958
rect 33140 31894 33192 31900
rect 33048 31816 33100 31822
rect 33048 31758 33100 31764
rect 32956 31748 33008 31754
rect 32956 31690 33008 31696
rect 32968 31482 32996 31690
rect 32956 31476 33008 31482
rect 32956 31418 33008 31424
rect 32968 31142 32996 31418
rect 32956 31136 33008 31142
rect 32956 31078 33008 31084
rect 32968 30734 32996 31078
rect 32956 30728 33008 30734
rect 32956 30670 33008 30676
rect 32864 30660 32916 30666
rect 32864 30602 32916 30608
rect 33060 29850 33088 31758
rect 33140 31340 33192 31346
rect 33140 31282 33192 31288
rect 33048 29844 33100 29850
rect 33048 29786 33100 29792
rect 32772 29776 32824 29782
rect 32772 29718 32824 29724
rect 32312 28076 32364 28082
rect 32312 28018 32364 28024
rect 32680 28076 32732 28082
rect 32680 28018 32732 28024
rect 32128 27464 32180 27470
rect 32128 27406 32180 27412
rect 32404 27464 32456 27470
rect 32404 27406 32456 27412
rect 32140 27062 32168 27406
rect 32416 27062 32444 27406
rect 32128 27056 32180 27062
rect 32128 26998 32180 27004
rect 32404 27056 32456 27062
rect 32404 26998 32456 27004
rect 32784 26586 32812 29718
rect 33152 29646 33180 31282
rect 33140 29640 33192 29646
rect 33140 29582 33192 29588
rect 32956 28552 33008 28558
rect 32956 28494 33008 28500
rect 32968 27130 32996 28494
rect 32956 27124 33008 27130
rect 32956 27066 33008 27072
rect 31300 26580 31352 26586
rect 31300 26522 31352 26528
rect 31668 26580 31720 26586
rect 31668 26522 31720 26528
rect 32772 26580 32824 26586
rect 32772 26522 32824 26528
rect 31392 26376 31444 26382
rect 31392 26318 31444 26324
rect 31300 26240 31352 26246
rect 31300 26182 31352 26188
rect 31312 25294 31340 26182
rect 31404 25906 31432 26318
rect 31760 26308 31812 26314
rect 31760 26250 31812 26256
rect 31772 25906 31800 26250
rect 32784 26042 32812 26522
rect 32772 26036 32824 26042
rect 32772 25978 32824 25984
rect 32784 25906 32812 25978
rect 31392 25900 31444 25906
rect 31392 25842 31444 25848
rect 31760 25900 31812 25906
rect 31760 25842 31812 25848
rect 32772 25900 32824 25906
rect 32772 25842 32824 25848
rect 32220 25696 32272 25702
rect 32220 25638 32272 25644
rect 32232 25498 32260 25638
rect 32220 25492 32272 25498
rect 32220 25434 32272 25440
rect 32784 25430 32812 25842
rect 32772 25424 32824 25430
rect 32772 25366 32824 25372
rect 31300 25288 31352 25294
rect 31300 25230 31352 25236
rect 31300 25152 31352 25158
rect 31300 25094 31352 25100
rect 31312 24886 31340 25094
rect 32784 24954 32812 25366
rect 32772 24948 32824 24954
rect 32772 24890 32824 24896
rect 31300 24880 31352 24886
rect 31300 24822 31352 24828
rect 33244 22094 33272 33816
rect 33324 33652 33376 33658
rect 33324 33594 33376 33600
rect 33336 33386 33364 33594
rect 33428 33522 33456 34342
rect 33416 33516 33468 33522
rect 33416 33458 33468 33464
rect 33520 33402 33548 36110
rect 33324 33380 33376 33386
rect 33324 33322 33376 33328
rect 33428 33374 33548 33402
rect 33324 32564 33376 32570
rect 33324 32506 33376 32512
rect 33336 29850 33364 32506
rect 33428 31686 33456 33374
rect 33704 33114 33732 36314
rect 33796 36310 33824 36586
rect 33784 36304 33836 36310
rect 33784 36246 33836 36252
rect 33888 36242 33916 37062
rect 33980 36922 34008 37810
rect 34164 37670 34192 38898
rect 34152 37664 34204 37670
rect 34152 37606 34204 37612
rect 34256 37346 34284 41006
rect 34072 37318 34284 37346
rect 33968 36916 34020 36922
rect 33968 36858 34020 36864
rect 33968 36712 34020 36718
rect 33968 36654 34020 36660
rect 33980 36582 34008 36654
rect 33968 36576 34020 36582
rect 33968 36518 34020 36524
rect 33876 36236 33928 36242
rect 33876 36178 33928 36184
rect 33888 35544 33916 36178
rect 33968 35692 34020 35698
rect 34072 35680 34100 37318
rect 34244 37256 34296 37262
rect 34348 37244 34376 41958
rect 34440 41682 34468 42520
rect 34428 41676 34480 41682
rect 34428 41618 34480 41624
rect 34428 41472 34480 41478
rect 34428 41414 34480 41420
rect 34440 41274 34468 41414
rect 34428 41268 34480 41274
rect 34428 41210 34480 41216
rect 34428 39568 34480 39574
rect 34428 39510 34480 39516
rect 34440 38962 34468 39510
rect 34428 38956 34480 38962
rect 34428 38898 34480 38904
rect 34296 37216 34376 37244
rect 34244 37198 34296 37204
rect 34256 36786 34284 37198
rect 34244 36780 34296 36786
rect 34244 36722 34296 36728
rect 34152 36576 34204 36582
rect 34152 36518 34204 36524
rect 34164 35698 34192 36518
rect 34256 36281 34284 36722
rect 34242 36272 34298 36281
rect 34242 36207 34298 36216
rect 34336 36168 34388 36174
rect 34336 36110 34388 36116
rect 34348 35834 34376 36110
rect 34428 36032 34480 36038
rect 34428 35974 34480 35980
rect 34336 35828 34388 35834
rect 34336 35770 34388 35776
rect 34020 35652 34100 35680
rect 33968 35634 34020 35640
rect 33888 35516 34008 35544
rect 33692 33108 33744 33114
rect 33692 33050 33744 33056
rect 33508 32904 33560 32910
rect 33508 32846 33560 32852
rect 33416 31680 33468 31686
rect 33416 31622 33468 31628
rect 33520 31362 33548 32846
rect 33600 32496 33652 32502
rect 33600 32438 33652 32444
rect 33428 31334 33548 31362
rect 33428 31278 33456 31334
rect 33416 31272 33468 31278
rect 33416 31214 33468 31220
rect 33324 29844 33376 29850
rect 33324 29786 33376 29792
rect 33336 29714 33364 29786
rect 33324 29708 33376 29714
rect 33324 29650 33376 29656
rect 33428 29578 33456 31214
rect 33612 29594 33640 32438
rect 33784 31884 33836 31890
rect 33784 31826 33836 31832
rect 33796 31278 33824 31826
rect 33876 31816 33928 31822
rect 33876 31758 33928 31764
rect 33888 31482 33916 31758
rect 33876 31476 33928 31482
rect 33876 31418 33928 31424
rect 33784 31272 33836 31278
rect 33784 31214 33836 31220
rect 33796 30802 33824 31214
rect 33784 30796 33836 30802
rect 33784 30738 33836 30744
rect 33796 29714 33824 30738
rect 33784 29708 33836 29714
rect 33784 29650 33836 29656
rect 33416 29572 33468 29578
rect 33416 29514 33468 29520
rect 33520 29566 33640 29594
rect 33324 29504 33376 29510
rect 33324 29446 33376 29452
rect 33336 28506 33364 29446
rect 33520 28994 33548 29566
rect 33612 29306 33916 29322
rect 33600 29300 33928 29306
rect 33652 29294 33876 29300
rect 33600 29242 33652 29248
rect 33876 29242 33928 29248
rect 33428 28966 33548 28994
rect 33980 28966 34008 35516
rect 34072 35494 34100 35652
rect 34152 35692 34204 35698
rect 34152 35634 34204 35640
rect 34060 35488 34112 35494
rect 34112 35448 34192 35476
rect 34060 35430 34112 35436
rect 34060 33380 34112 33386
rect 34060 33322 34112 33328
rect 34072 32026 34100 33322
rect 34164 32570 34192 35448
rect 34336 34944 34388 34950
rect 34336 34886 34388 34892
rect 34348 34678 34376 34886
rect 34336 34672 34388 34678
rect 34336 34614 34388 34620
rect 34336 33856 34388 33862
rect 34336 33798 34388 33804
rect 34348 33454 34376 33798
rect 34336 33448 34388 33454
rect 34336 33390 34388 33396
rect 34244 32972 34296 32978
rect 34244 32914 34296 32920
rect 34152 32564 34204 32570
rect 34152 32506 34204 32512
rect 34060 32020 34112 32026
rect 34060 31962 34112 31968
rect 34060 31748 34112 31754
rect 34060 31690 34112 31696
rect 34072 31346 34100 31690
rect 34060 31340 34112 31346
rect 34060 31282 34112 31288
rect 34072 30734 34100 31282
rect 34060 30728 34112 30734
rect 34060 30670 34112 30676
rect 34072 30394 34100 30670
rect 34060 30388 34112 30394
rect 34060 30330 34112 30336
rect 34152 29844 34204 29850
rect 34152 29786 34204 29792
rect 33428 28626 33456 28966
rect 33968 28960 34020 28966
rect 33968 28902 34020 28908
rect 33966 28792 34022 28801
rect 33966 28727 34022 28736
rect 33416 28620 33468 28626
rect 33416 28562 33468 28568
rect 33980 28558 34008 28727
rect 33968 28552 34020 28558
rect 33336 28478 33456 28506
rect 33968 28494 34020 28500
rect 33324 26308 33376 26314
rect 33324 26250 33376 26256
rect 33336 26042 33364 26250
rect 33324 26036 33376 26042
rect 33324 25978 33376 25984
rect 33152 22066 33272 22094
rect 33428 22094 33456 28478
rect 33980 28150 34008 28494
rect 33968 28144 34020 28150
rect 33968 28086 34020 28092
rect 33784 27464 33836 27470
rect 33784 27406 33836 27412
rect 33796 27062 33824 27406
rect 33784 27056 33836 27062
rect 33784 26998 33836 27004
rect 33796 26586 33824 26998
rect 33784 26580 33836 26586
rect 33784 26522 33836 26528
rect 33796 26042 33824 26522
rect 33784 26036 33836 26042
rect 33784 25978 33836 25984
rect 33428 22066 33548 22094
rect 33152 18086 33180 22066
rect 33140 18080 33192 18086
rect 33140 18022 33192 18028
rect 33520 3466 33548 22066
rect 33980 11082 34008 28086
rect 34164 27962 34192 29786
rect 34256 28014 34284 32914
rect 34336 32224 34388 32230
rect 34336 32166 34388 32172
rect 34348 31958 34376 32166
rect 34336 31952 34388 31958
rect 34336 31894 34388 31900
rect 34440 29102 34468 35974
rect 34532 33810 34560 43438
rect 34612 42152 34664 42158
rect 34612 42094 34664 42100
rect 34624 40730 34652 42094
rect 34716 41664 34744 45222
rect 34808 45082 34836 45358
rect 35348 45348 35400 45354
rect 35348 45290 35400 45296
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34796 45076 34848 45082
rect 34796 45018 34848 45024
rect 35360 44946 35388 45290
rect 35348 44940 35400 44946
rect 35348 44882 35400 44888
rect 34888 44872 34940 44878
rect 35544 44826 35572 48010
rect 35808 47456 35860 47462
rect 35808 47398 35860 47404
rect 35820 47258 35848 47398
rect 35808 47252 35860 47258
rect 35808 47194 35860 47200
rect 35808 46572 35860 46578
rect 35912 46560 35940 49030
rect 35860 46532 35940 46560
rect 35808 46514 35860 46520
rect 35820 45966 35848 46514
rect 35808 45960 35860 45966
rect 35808 45902 35860 45908
rect 35808 45824 35860 45830
rect 35808 45766 35860 45772
rect 35820 45422 35848 45766
rect 35808 45416 35860 45422
rect 35808 45358 35860 45364
rect 35624 44940 35676 44946
rect 35624 44882 35676 44888
rect 34888 44814 34940 44820
rect 34796 44804 34848 44810
rect 34796 44746 34848 44752
rect 34808 44538 34836 44746
rect 34900 44538 34928 44814
rect 35360 44798 35572 44826
rect 34796 44532 34848 44538
rect 34796 44474 34848 44480
rect 34888 44532 34940 44538
rect 34888 44474 34940 44480
rect 34796 44192 34848 44198
rect 34796 44134 34848 44140
rect 34808 43994 34836 44134
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 34796 43988 34848 43994
rect 34796 43930 34848 43936
rect 34796 43852 34848 43858
rect 34796 43794 34848 43800
rect 34808 42702 34836 43794
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 35360 42922 35388 44798
rect 35532 43308 35584 43314
rect 35532 43250 35584 43256
rect 35268 42894 35388 42922
rect 35544 42906 35572 43250
rect 35532 42900 35584 42906
rect 34796 42696 34848 42702
rect 34796 42638 34848 42644
rect 34808 42022 34836 42638
rect 34980 42628 35032 42634
rect 34980 42570 35032 42576
rect 34992 42362 35020 42570
rect 34980 42356 35032 42362
rect 34980 42298 35032 42304
rect 35268 42106 35296 42894
rect 35532 42842 35584 42848
rect 35348 42696 35400 42702
rect 35348 42638 35400 42644
rect 35532 42696 35584 42702
rect 35532 42638 35584 42644
rect 35360 42294 35388 42638
rect 35348 42288 35400 42294
rect 35348 42230 35400 42236
rect 35268 42078 35388 42106
rect 35544 42090 35572 42638
rect 34796 42016 34848 42022
rect 34796 41958 34848 41964
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 35360 41834 35388 42078
rect 35532 42084 35584 42090
rect 35532 42026 35584 42032
rect 35360 41806 35480 41834
rect 34716 41636 34836 41664
rect 34704 41132 34756 41138
rect 34704 41074 34756 41080
rect 34612 40724 34664 40730
rect 34612 40666 34664 40672
rect 34716 40526 34744 41074
rect 34704 40520 34756 40526
rect 34704 40462 34756 40468
rect 34808 40050 34836 41636
rect 35348 41472 35400 41478
rect 35348 41414 35400 41420
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 35360 40526 35388 41414
rect 35348 40520 35400 40526
rect 35348 40462 35400 40468
rect 35348 40384 35400 40390
rect 35348 40326 35400 40332
rect 34796 40044 34848 40050
rect 34796 39986 34848 39992
rect 34808 39438 34836 39986
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 35360 39642 35388 40326
rect 35348 39636 35400 39642
rect 35348 39578 35400 39584
rect 35348 39500 35400 39506
rect 35348 39442 35400 39448
rect 34796 39432 34848 39438
rect 34796 39374 34848 39380
rect 35256 39432 35308 39438
rect 35256 39374 35308 39380
rect 34980 39364 35032 39370
rect 34980 39306 35032 39312
rect 34704 39296 34756 39302
rect 34704 39238 34756 39244
rect 34716 38282 34744 39238
rect 34992 39030 35020 39306
rect 34980 39024 35032 39030
rect 34980 38966 35032 38972
rect 35268 38962 35296 39374
rect 35256 38956 35308 38962
rect 35256 38898 35308 38904
rect 34796 38752 34848 38758
rect 34796 38694 34848 38700
rect 34808 38554 34836 38694
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 35360 38554 35388 39442
rect 34796 38548 34848 38554
rect 34796 38490 34848 38496
rect 35348 38548 35400 38554
rect 35348 38490 35400 38496
rect 35360 38350 35388 38490
rect 35348 38344 35400 38350
rect 35348 38286 35400 38292
rect 34704 38276 34756 38282
rect 34704 38218 34756 38224
rect 35164 38276 35216 38282
rect 35164 38218 35216 38224
rect 35176 38010 35204 38218
rect 35164 38004 35216 38010
rect 35164 37946 35216 37952
rect 34612 37868 34664 37874
rect 34612 37810 34664 37816
rect 34624 37398 34652 37810
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34704 37460 34756 37466
rect 34704 37402 34756 37408
rect 34612 37392 34664 37398
rect 34612 37334 34664 37340
rect 34624 36378 34652 37334
rect 34716 37262 34744 37402
rect 34888 37392 34940 37398
rect 34888 37334 34940 37340
rect 34704 37256 34756 37262
rect 34704 37198 34756 37204
rect 34716 36718 34744 37198
rect 34796 37120 34848 37126
rect 34796 37062 34848 37068
rect 34808 36854 34836 37062
rect 34796 36848 34848 36854
rect 34796 36790 34848 36796
rect 34704 36712 34756 36718
rect 34900 36666 34928 37334
rect 35072 37256 35124 37262
rect 35072 37198 35124 37204
rect 35084 36922 35112 37198
rect 35348 37188 35400 37194
rect 35348 37130 35400 37136
rect 35072 36916 35124 36922
rect 35072 36858 35124 36864
rect 35164 36780 35216 36786
rect 35164 36722 35216 36728
rect 34704 36654 34756 36660
rect 34808 36638 34928 36666
rect 34612 36372 34664 36378
rect 34612 36314 34664 36320
rect 34624 35630 34652 36314
rect 34704 35828 34756 35834
rect 34704 35770 34756 35776
rect 34612 35624 34664 35630
rect 34612 35566 34664 35572
rect 34612 35080 34664 35086
rect 34610 35048 34612 35057
rect 34664 35048 34666 35057
rect 34610 34983 34666 34992
rect 34612 34672 34664 34678
rect 34612 34614 34664 34620
rect 34624 33998 34652 34614
rect 34716 34542 34744 35770
rect 34808 35086 34836 36638
rect 35176 36582 35204 36722
rect 35360 36582 35388 37130
rect 35164 36576 35216 36582
rect 35164 36518 35216 36524
rect 35348 36576 35400 36582
rect 35348 36518 35400 36524
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34888 36304 34940 36310
rect 34888 36246 34940 36252
rect 35070 36272 35126 36281
rect 34900 36106 34928 36246
rect 35070 36207 35126 36216
rect 35164 36236 35216 36242
rect 34888 36100 34940 36106
rect 34888 36042 34940 36048
rect 35084 35698 35112 36207
rect 35164 36178 35216 36184
rect 35072 35692 35124 35698
rect 35072 35634 35124 35640
rect 35176 35630 35204 36178
rect 35360 35766 35388 36518
rect 35348 35760 35400 35766
rect 35348 35702 35400 35708
rect 35164 35624 35216 35630
rect 35164 35566 35216 35572
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35346 35184 35402 35193
rect 35346 35119 35402 35128
rect 35360 35086 35388 35119
rect 34796 35080 34848 35086
rect 34796 35022 34848 35028
rect 35348 35080 35400 35086
rect 35348 35022 35400 35028
rect 35348 34944 35400 34950
rect 35348 34886 35400 34892
rect 35360 34610 35388 34886
rect 34796 34604 34848 34610
rect 34796 34546 34848 34552
rect 35348 34604 35400 34610
rect 35348 34546 35400 34552
rect 34704 34536 34756 34542
rect 34704 34478 34756 34484
rect 34716 34134 34744 34478
rect 34704 34128 34756 34134
rect 34704 34070 34756 34076
rect 34612 33992 34664 33998
rect 34612 33934 34664 33940
rect 34532 33782 34652 33810
rect 34520 33584 34572 33590
rect 34520 33526 34572 33532
rect 34428 29096 34480 29102
rect 34428 29038 34480 29044
rect 34428 28076 34480 28082
rect 34428 28018 34480 28024
rect 34072 27946 34192 27962
rect 34244 28008 34296 28014
rect 34244 27950 34296 27956
rect 34060 27940 34192 27946
rect 34112 27934 34192 27940
rect 34060 27882 34112 27888
rect 34164 27538 34192 27934
rect 34152 27532 34204 27538
rect 34152 27474 34204 27480
rect 34336 26988 34388 26994
rect 34336 26930 34388 26936
rect 34060 26920 34112 26926
rect 34060 26862 34112 26868
rect 34072 26450 34100 26862
rect 34060 26444 34112 26450
rect 34060 26386 34112 26392
rect 34348 26042 34376 26930
rect 34336 26036 34388 26042
rect 34336 25978 34388 25984
rect 33968 11076 34020 11082
rect 33968 11018 34020 11024
rect 33508 3460 33560 3466
rect 33508 3402 33560 3408
rect 34440 2990 34468 28018
rect 34532 15910 34560 33526
rect 34624 26994 34652 33782
rect 34808 33658 34836 34546
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35360 34202 35388 34546
rect 35348 34196 35400 34202
rect 35348 34138 35400 34144
rect 35348 33992 35400 33998
rect 35348 33934 35400 33940
rect 34704 33652 34756 33658
rect 34704 33594 34756 33600
rect 34796 33652 34848 33658
rect 34796 33594 34848 33600
rect 35256 33652 35308 33658
rect 35256 33594 35308 33600
rect 34716 32230 34744 33594
rect 35268 33522 35296 33594
rect 35256 33516 35308 33522
rect 35256 33458 35308 33464
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35360 33114 35388 33934
rect 35348 33108 35400 33114
rect 35348 33050 35400 33056
rect 35072 32904 35124 32910
rect 35072 32846 35124 32852
rect 35084 32502 35112 32846
rect 35072 32496 35124 32502
rect 35072 32438 35124 32444
rect 34704 32224 34756 32230
rect 34704 32166 34756 32172
rect 34716 31822 34744 32166
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34704 31816 34756 31822
rect 34704 31758 34756 31764
rect 35452 31754 35480 41806
rect 35544 40202 35572 42026
rect 35636 40390 35664 44882
rect 35716 44872 35768 44878
rect 35716 44814 35768 44820
rect 35728 44334 35756 44814
rect 35820 44810 35848 45358
rect 35808 44804 35860 44810
rect 35808 44746 35860 44752
rect 35716 44328 35768 44334
rect 35716 44270 35768 44276
rect 35716 44192 35768 44198
rect 35716 44134 35768 44140
rect 35728 41818 35756 44134
rect 35900 43852 35952 43858
rect 35900 43794 35952 43800
rect 35912 43246 35940 43794
rect 35992 43376 36044 43382
rect 35992 43318 36044 43324
rect 35900 43240 35952 43246
rect 35900 43182 35952 43188
rect 36004 42906 36032 43318
rect 35992 42900 36044 42906
rect 35992 42842 36044 42848
rect 35898 42800 35954 42809
rect 35898 42735 35954 42744
rect 35808 42356 35860 42362
rect 35808 42298 35860 42304
rect 35716 41812 35768 41818
rect 35716 41754 35768 41760
rect 35728 40474 35756 41754
rect 35820 41478 35848 42298
rect 35912 42226 35940 42735
rect 35900 42220 35952 42226
rect 35900 42162 35952 42168
rect 35992 42220 36044 42226
rect 35992 42162 36044 42168
rect 36004 41614 36032 42162
rect 35992 41608 36044 41614
rect 35992 41550 36044 41556
rect 35808 41472 35860 41478
rect 35808 41414 35860 41420
rect 35900 41132 35952 41138
rect 35900 41074 35952 41080
rect 35808 40928 35860 40934
rect 35808 40870 35860 40876
rect 35820 40594 35848 40870
rect 35912 40662 35940 41074
rect 35900 40656 35952 40662
rect 35900 40598 35952 40604
rect 35808 40588 35860 40594
rect 35808 40530 35860 40536
rect 35728 40446 35940 40474
rect 35624 40384 35676 40390
rect 35624 40326 35676 40332
rect 35544 40174 35756 40202
rect 35624 39840 35676 39846
rect 35624 39782 35676 39788
rect 35636 39438 35664 39782
rect 35624 39432 35676 39438
rect 35624 39374 35676 39380
rect 35532 39024 35584 39030
rect 35532 38966 35584 38972
rect 35544 38214 35572 38966
rect 35636 38962 35664 39374
rect 35624 38956 35676 38962
rect 35624 38898 35676 38904
rect 35532 38208 35584 38214
rect 35532 38150 35584 38156
rect 35544 38010 35572 38150
rect 35532 38004 35584 38010
rect 35532 37946 35584 37952
rect 35532 36780 35584 36786
rect 35532 36722 35584 36728
rect 35544 36174 35572 36722
rect 35728 36394 35756 40174
rect 35808 39908 35860 39914
rect 35808 39850 35860 39856
rect 35820 39302 35848 39850
rect 35808 39296 35860 39302
rect 35808 39238 35860 39244
rect 35820 38486 35848 39238
rect 35808 38480 35860 38486
rect 35808 38422 35860 38428
rect 35820 37874 35848 38422
rect 35912 38282 35940 40446
rect 35992 38752 36044 38758
rect 35992 38694 36044 38700
rect 35900 38276 35952 38282
rect 35900 38218 35952 38224
rect 35808 37868 35860 37874
rect 35808 37810 35860 37816
rect 36004 37466 36032 38694
rect 35992 37460 36044 37466
rect 35992 37402 36044 37408
rect 35636 36366 35756 36394
rect 35532 36168 35584 36174
rect 35532 36110 35584 36116
rect 35532 35080 35584 35086
rect 35532 35022 35584 35028
rect 35544 33998 35572 35022
rect 35532 33992 35584 33998
rect 35532 33934 35584 33940
rect 35544 33658 35572 33934
rect 35532 33652 35584 33658
rect 35532 33594 35584 33600
rect 35544 32842 35572 33594
rect 35636 33590 35664 36366
rect 35808 36236 35860 36242
rect 35808 36178 35860 36184
rect 35820 35290 35848 36178
rect 36004 36106 36032 37402
rect 35992 36100 36044 36106
rect 35992 36042 36044 36048
rect 35808 35284 35860 35290
rect 35808 35226 35860 35232
rect 36096 35154 36124 53926
rect 36176 53780 36228 53786
rect 36176 53722 36228 53728
rect 36188 49638 36216 53722
rect 37280 51808 37332 51814
rect 37280 51750 37332 51756
rect 36452 51468 36504 51474
rect 36452 51410 36504 51416
rect 36176 49632 36228 49638
rect 36176 49574 36228 49580
rect 36176 44872 36228 44878
rect 36176 44814 36228 44820
rect 36188 44538 36216 44814
rect 36268 44804 36320 44810
rect 36268 44746 36320 44752
rect 36176 44532 36228 44538
rect 36176 44474 36228 44480
rect 36280 44402 36308 44746
rect 36268 44396 36320 44402
rect 36268 44338 36320 44344
rect 36280 43926 36308 44338
rect 36268 43920 36320 43926
rect 36268 43862 36320 43868
rect 36464 43790 36492 51410
rect 37188 51264 37240 51270
rect 37188 51206 37240 51212
rect 37200 50794 37228 51206
rect 37188 50788 37240 50794
rect 37188 50730 37240 50736
rect 37200 50522 37228 50730
rect 37292 50726 37320 51750
rect 37280 50720 37332 50726
rect 37280 50662 37332 50668
rect 37188 50516 37240 50522
rect 37188 50458 37240 50464
rect 36912 49768 36964 49774
rect 36912 49710 36964 49716
rect 36544 48544 36596 48550
rect 36544 48486 36596 48492
rect 36556 48142 36584 48486
rect 36544 48136 36596 48142
rect 36544 48078 36596 48084
rect 36556 48006 36584 48078
rect 36544 48000 36596 48006
rect 36544 47942 36596 47948
rect 36556 46918 36584 47942
rect 36544 46912 36596 46918
rect 36544 46854 36596 46860
rect 36556 45830 36584 46854
rect 36636 46504 36688 46510
rect 36636 46446 36688 46452
rect 36648 46374 36676 46446
rect 36636 46368 36688 46374
rect 36636 46310 36688 46316
rect 36544 45824 36596 45830
rect 36544 45766 36596 45772
rect 36544 44872 36596 44878
rect 36544 44814 36596 44820
rect 36556 44402 36584 44814
rect 36648 44538 36676 46310
rect 36636 44532 36688 44538
rect 36636 44474 36688 44480
rect 36544 44396 36596 44402
rect 36544 44338 36596 44344
rect 36556 43994 36584 44338
rect 36728 44260 36780 44266
rect 36728 44202 36780 44208
rect 36544 43988 36596 43994
rect 36544 43930 36596 43936
rect 36268 43784 36320 43790
rect 36268 43726 36320 43732
rect 36452 43784 36504 43790
rect 36452 43726 36504 43732
rect 36280 43314 36308 43726
rect 36740 43654 36768 44202
rect 36728 43648 36780 43654
rect 36728 43590 36780 43596
rect 36268 43308 36320 43314
rect 36268 43250 36320 43256
rect 36176 43104 36228 43110
rect 36176 43046 36228 43052
rect 36360 43104 36412 43110
rect 36360 43046 36412 43052
rect 36188 40730 36216 43046
rect 36268 42832 36320 42838
rect 36268 42774 36320 42780
rect 36280 41546 36308 42774
rect 36372 41682 36400 43046
rect 36452 42900 36504 42906
rect 36452 42842 36504 42848
rect 36464 42702 36492 42842
rect 36740 42770 36768 43590
rect 36728 42764 36780 42770
rect 36728 42706 36780 42712
rect 36820 42764 36872 42770
rect 36820 42706 36872 42712
rect 36452 42696 36504 42702
rect 36452 42638 36504 42644
rect 36832 42294 36860 42706
rect 36820 42288 36872 42294
rect 36820 42230 36872 42236
rect 36360 41676 36412 41682
rect 36360 41618 36412 41624
rect 36268 41540 36320 41546
rect 36268 41482 36320 41488
rect 36360 41472 36412 41478
rect 36360 41414 36412 41420
rect 36728 41472 36780 41478
rect 36728 41414 36780 41420
rect 36176 40724 36228 40730
rect 36176 40666 36228 40672
rect 36372 40050 36400 41414
rect 36636 41268 36688 41274
rect 36636 41210 36688 41216
rect 36648 40526 36676 41210
rect 36740 41138 36768 41414
rect 36728 41132 36780 41138
rect 36728 41074 36780 41080
rect 36740 40526 36768 41074
rect 36636 40520 36688 40526
rect 36636 40462 36688 40468
rect 36728 40520 36780 40526
rect 36728 40462 36780 40468
rect 36176 40044 36228 40050
rect 36176 39986 36228 39992
rect 36360 40044 36412 40050
rect 36360 39986 36412 39992
rect 36188 39506 36216 39986
rect 36176 39500 36228 39506
rect 36176 39442 36228 39448
rect 36372 39438 36400 39986
rect 36360 39432 36412 39438
rect 36360 39374 36412 39380
rect 36360 39092 36412 39098
rect 36360 39034 36412 39040
rect 36372 37466 36400 39034
rect 36452 38752 36504 38758
rect 36452 38694 36504 38700
rect 36464 38554 36492 38694
rect 36452 38548 36504 38554
rect 36452 38490 36504 38496
rect 36464 37874 36492 38490
rect 36636 38208 36688 38214
rect 36636 38150 36688 38156
rect 36452 37868 36504 37874
rect 36452 37810 36504 37816
rect 36648 37466 36676 38150
rect 36360 37460 36412 37466
rect 36360 37402 36412 37408
rect 36636 37460 36688 37466
rect 36636 37402 36688 37408
rect 36648 36718 36676 37402
rect 36636 36712 36688 36718
rect 36636 36654 36688 36660
rect 36176 36168 36228 36174
rect 36176 36110 36228 36116
rect 36188 35630 36216 36110
rect 36636 35828 36688 35834
rect 36636 35770 36688 35776
rect 36452 35692 36504 35698
rect 36452 35634 36504 35640
rect 36176 35624 36228 35630
rect 36176 35566 36228 35572
rect 36084 35148 36136 35154
rect 36084 35090 36136 35096
rect 36464 35018 36492 35634
rect 36544 35216 36596 35222
rect 36544 35158 36596 35164
rect 36452 35012 36504 35018
rect 36452 34954 36504 34960
rect 36464 34610 36492 34954
rect 36556 34746 36584 35158
rect 36648 34950 36676 35770
rect 36636 34944 36688 34950
rect 36636 34886 36688 34892
rect 36544 34740 36596 34746
rect 36544 34682 36596 34688
rect 35808 34604 35860 34610
rect 35808 34546 35860 34552
rect 35992 34604 36044 34610
rect 35992 34546 36044 34552
rect 36452 34604 36504 34610
rect 36452 34546 36504 34552
rect 35716 33856 35768 33862
rect 35716 33798 35768 33804
rect 35624 33584 35676 33590
rect 35624 33526 35676 33532
rect 35728 32910 35756 33798
rect 35716 32904 35768 32910
rect 35716 32846 35768 32852
rect 35532 32836 35584 32842
rect 35532 32778 35584 32784
rect 35716 32768 35768 32774
rect 35716 32710 35768 32716
rect 35728 32434 35756 32710
rect 35820 32570 35848 34546
rect 35900 34400 35952 34406
rect 35900 34342 35952 34348
rect 35912 34066 35940 34342
rect 35900 34060 35952 34066
rect 35900 34002 35952 34008
rect 35912 33454 35940 34002
rect 36004 33930 36032 34546
rect 36556 34202 36584 34682
rect 36544 34196 36596 34202
rect 36544 34138 36596 34144
rect 35992 33924 36044 33930
rect 35992 33866 36044 33872
rect 36004 33658 36032 33866
rect 35992 33652 36044 33658
rect 35992 33594 36044 33600
rect 36556 33590 36584 34138
rect 36544 33584 36596 33590
rect 36544 33526 36596 33532
rect 36084 33516 36136 33522
rect 36084 33458 36136 33464
rect 36176 33516 36228 33522
rect 36176 33458 36228 33464
rect 35900 33448 35952 33454
rect 35900 33390 35952 33396
rect 36096 33114 36124 33458
rect 36084 33108 36136 33114
rect 36084 33050 36136 33056
rect 35808 32564 35860 32570
rect 35808 32506 35860 32512
rect 36096 32434 36124 33050
rect 36188 32502 36216 33458
rect 36636 32768 36688 32774
rect 36636 32710 36688 32716
rect 36728 32768 36780 32774
rect 36728 32710 36780 32716
rect 36176 32496 36228 32502
rect 36176 32438 36228 32444
rect 36648 32434 36676 32710
rect 35716 32428 35768 32434
rect 35716 32370 35768 32376
rect 36084 32428 36136 32434
rect 36084 32370 36136 32376
rect 36268 32428 36320 32434
rect 36268 32370 36320 32376
rect 36636 32428 36688 32434
rect 36636 32370 36688 32376
rect 34808 31726 35480 31754
rect 34704 31272 34756 31278
rect 34704 31214 34756 31220
rect 34716 30938 34744 31214
rect 34704 30932 34756 30938
rect 34704 30874 34756 30880
rect 34612 26988 34664 26994
rect 34612 26930 34664 26936
rect 34808 22574 34836 31726
rect 35728 31414 35756 32370
rect 36280 31958 36308 32370
rect 36360 32224 36412 32230
rect 36360 32166 36412 32172
rect 36268 31952 36320 31958
rect 36268 31894 36320 31900
rect 35992 31748 36044 31754
rect 35992 31690 36044 31696
rect 35716 31408 35768 31414
rect 35716 31350 35768 31356
rect 35440 31340 35492 31346
rect 35440 31282 35492 31288
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35452 30734 35480 31282
rect 35728 30734 35756 31350
rect 35440 30728 35492 30734
rect 35440 30670 35492 30676
rect 35716 30728 35768 30734
rect 35716 30670 35768 30676
rect 35164 30252 35216 30258
rect 35164 30194 35216 30200
rect 35176 30036 35204 30194
rect 35176 30008 35388 30036
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35360 29102 35388 30008
rect 35348 29096 35400 29102
rect 35348 29038 35400 29044
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35360 28558 35388 29038
rect 34980 28552 35032 28558
rect 34978 28520 34980 28529
rect 35348 28552 35400 28558
rect 35032 28520 35034 28529
rect 35348 28494 35400 28500
rect 34978 28455 35034 28464
rect 35360 28218 35388 28494
rect 35348 28212 35400 28218
rect 35348 28154 35400 28160
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35348 27464 35400 27470
rect 35348 27406 35400 27412
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35360 26382 35388 27406
rect 35348 26376 35400 26382
rect 35348 26318 35400 26324
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34796 22568 34848 22574
rect 34796 22510 34848 22516
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35452 22094 35480 30670
rect 35716 30252 35768 30258
rect 35716 30194 35768 30200
rect 35728 29646 35756 30194
rect 35808 30184 35860 30190
rect 35808 30126 35860 30132
rect 35716 29640 35768 29646
rect 35716 29582 35768 29588
rect 35728 29186 35756 29582
rect 35636 29158 35756 29186
rect 35636 29102 35664 29158
rect 35624 29096 35676 29102
rect 35624 29038 35676 29044
rect 35532 28688 35584 28694
rect 35532 28630 35584 28636
rect 35544 28490 35572 28630
rect 35532 28484 35584 28490
rect 35532 28426 35584 28432
rect 35544 28082 35572 28426
rect 35636 28150 35664 29038
rect 35820 29034 35848 30126
rect 36004 30054 36032 31690
rect 36280 31346 36308 31894
rect 36268 31340 36320 31346
rect 36268 31282 36320 31288
rect 36084 30932 36136 30938
rect 36084 30874 36136 30880
rect 36096 30258 36124 30874
rect 36176 30592 36228 30598
rect 36176 30534 36228 30540
rect 36084 30252 36136 30258
rect 36084 30194 36136 30200
rect 35992 30048 36044 30054
rect 35992 29990 36044 29996
rect 36188 29714 36216 30534
rect 36280 30394 36308 31282
rect 36372 30802 36400 32166
rect 36648 31890 36676 32370
rect 36740 32366 36768 32710
rect 36728 32360 36780 32366
rect 36728 32302 36780 32308
rect 36636 31884 36688 31890
rect 36636 31826 36688 31832
rect 36740 31822 36768 32302
rect 36728 31816 36780 31822
rect 36728 31758 36780 31764
rect 36544 31340 36596 31346
rect 36544 31282 36596 31288
rect 36452 31204 36504 31210
rect 36452 31146 36504 31152
rect 36360 30796 36412 30802
rect 36360 30738 36412 30744
rect 36268 30388 36320 30394
rect 36268 30330 36320 30336
rect 36464 30258 36492 31146
rect 36556 30938 36584 31282
rect 36636 31136 36688 31142
rect 36636 31078 36688 31084
rect 36544 30932 36596 30938
rect 36544 30874 36596 30880
rect 36648 30802 36676 31078
rect 36636 30796 36688 30802
rect 36636 30738 36688 30744
rect 36452 30252 36504 30258
rect 36452 30194 36504 30200
rect 36452 30048 36504 30054
rect 36452 29990 36504 29996
rect 36464 29850 36492 29990
rect 36452 29844 36504 29850
rect 36452 29786 36504 29792
rect 36176 29708 36228 29714
rect 36176 29650 36228 29656
rect 36188 29170 36216 29650
rect 36648 29646 36676 30738
rect 36636 29640 36688 29646
rect 36636 29582 36688 29588
rect 36268 29504 36320 29510
rect 36268 29446 36320 29452
rect 36176 29164 36228 29170
rect 36176 29106 36228 29112
rect 35808 29028 35860 29034
rect 35808 28970 35860 28976
rect 35820 28762 35848 28970
rect 35808 28756 35860 28762
rect 35808 28698 35860 28704
rect 36280 28626 36308 29446
rect 36452 29096 36504 29102
rect 36452 29038 36504 29044
rect 36268 28620 36320 28626
rect 36268 28562 36320 28568
rect 35900 28552 35952 28558
rect 36464 28529 36492 29038
rect 35900 28494 35952 28500
rect 36450 28520 36506 28529
rect 35912 28422 35940 28494
rect 36450 28455 36506 28464
rect 35900 28416 35952 28422
rect 35900 28358 35952 28364
rect 35624 28144 35676 28150
rect 35624 28086 35676 28092
rect 35912 28082 35940 28358
rect 36464 28218 36492 28455
rect 36452 28212 36504 28218
rect 36452 28154 36504 28160
rect 35532 28076 35584 28082
rect 35532 28018 35584 28024
rect 35900 28076 35952 28082
rect 35900 28018 35952 28024
rect 36452 28076 36504 28082
rect 36452 28018 36504 28024
rect 35912 27334 35940 28018
rect 36464 27674 36492 28018
rect 36452 27668 36504 27674
rect 36452 27610 36504 27616
rect 35900 27328 35952 27334
rect 35900 27270 35952 27276
rect 35912 26790 35940 27270
rect 36084 26988 36136 26994
rect 36084 26930 36136 26936
rect 35900 26784 35952 26790
rect 35900 26726 35952 26732
rect 35360 22066 35480 22094
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34520 15904 34572 15910
rect 34520 15846 34572 15852
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34428 2984 34480 2990
rect 34428 2926 34480 2932
rect 31116 2916 31168 2922
rect 31116 2858 31168 2864
rect 32220 2848 32272 2854
rect 32220 2790 32272 2796
rect 34520 2848 34572 2854
rect 34520 2790 34572 2796
rect 30656 2508 30708 2514
rect 30656 2450 30708 2456
rect 32232 2446 32260 2790
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 32220 2440 32272 2446
rect 32220 2382 32272 2388
rect 28356 2032 28408 2038
rect 28356 1974 28408 1980
rect 30300 800 30328 2382
rect 32232 800 32260 2382
rect 34532 2378 34560 2790
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35360 2446 35388 22066
rect 35912 2582 35940 26726
rect 36096 26314 36124 26930
rect 36084 26308 36136 26314
rect 36084 26250 36136 26256
rect 36096 18698 36124 26250
rect 36084 18692 36136 18698
rect 36084 18634 36136 18640
rect 36924 2582 36952 49710
rect 37200 49434 37228 50458
rect 37292 50182 37320 50662
rect 37280 50176 37332 50182
rect 37280 50118 37332 50124
rect 37292 49774 37320 50118
rect 37280 49768 37332 49774
rect 37280 49710 37332 49716
rect 37188 49428 37240 49434
rect 37188 49370 37240 49376
rect 37464 47456 37516 47462
rect 37464 47398 37516 47404
rect 37188 47116 37240 47122
rect 37188 47058 37240 47064
rect 37200 43382 37228 47058
rect 37476 47025 37504 47398
rect 37462 47016 37518 47025
rect 37462 46951 37518 46960
rect 37280 46368 37332 46374
rect 37280 46310 37332 46316
rect 37292 45558 37320 46310
rect 37280 45552 37332 45558
rect 37280 45494 37332 45500
rect 37292 45082 37320 45494
rect 37280 45076 37332 45082
rect 37280 45018 37332 45024
rect 37188 43376 37240 43382
rect 37188 43318 37240 43324
rect 37372 43308 37424 43314
rect 37372 43250 37424 43256
rect 37188 43240 37240 43246
rect 37188 43182 37240 43188
rect 37002 42800 37058 42809
rect 37002 42735 37058 42744
rect 37016 42702 37044 42735
rect 37004 42696 37056 42702
rect 37004 42638 37056 42644
rect 37016 41682 37044 42638
rect 37200 42226 37228 43182
rect 37384 42294 37412 43250
rect 37476 42838 37504 46951
rect 37832 46368 37884 46374
rect 37832 46310 37884 46316
rect 37844 45966 37872 46310
rect 37832 45960 37884 45966
rect 37832 45902 37884 45908
rect 37740 45824 37792 45830
rect 37740 45766 37792 45772
rect 37752 45286 37780 45766
rect 37740 45280 37792 45286
rect 37740 45222 37792 45228
rect 37752 43058 37780 45222
rect 38108 45076 38160 45082
rect 38108 45018 38160 45024
rect 37832 43920 37884 43926
rect 37832 43862 37884 43868
rect 37844 43382 37872 43862
rect 37832 43376 37884 43382
rect 37832 43318 37884 43324
rect 37752 43030 37964 43058
rect 37464 42832 37516 42838
rect 37464 42774 37516 42780
rect 37464 42560 37516 42566
rect 37464 42502 37516 42508
rect 37372 42288 37424 42294
rect 37292 42236 37372 42242
rect 37292 42230 37424 42236
rect 37188 42220 37240 42226
rect 37188 42162 37240 42168
rect 37292 42214 37412 42230
rect 37200 41750 37228 42162
rect 37188 41744 37240 41750
rect 37188 41686 37240 41692
rect 37004 41676 37056 41682
rect 37004 41618 37056 41624
rect 37292 41414 37320 42214
rect 37372 42084 37424 42090
rect 37372 42026 37424 42032
rect 37384 41478 37412 42026
rect 37476 41546 37504 42502
rect 37832 42220 37884 42226
rect 37832 42162 37884 42168
rect 37556 42016 37608 42022
rect 37556 41958 37608 41964
rect 37464 41540 37516 41546
rect 37464 41482 37516 41488
rect 37372 41472 37424 41478
rect 37372 41414 37424 41420
rect 37200 41386 37320 41414
rect 37200 41274 37228 41386
rect 37188 41268 37240 41274
rect 37188 41210 37240 41216
rect 37096 40520 37148 40526
rect 37096 40462 37148 40468
rect 37108 31958 37136 40462
rect 37384 39438 37412 41414
rect 37568 40050 37596 41958
rect 37844 41138 37872 42162
rect 37832 41132 37884 41138
rect 37832 41074 37884 41080
rect 37648 40928 37700 40934
rect 37648 40870 37700 40876
rect 37556 40044 37608 40050
rect 37556 39986 37608 39992
rect 37464 39840 37516 39846
rect 37464 39782 37516 39788
rect 37372 39432 37424 39438
rect 37372 39374 37424 39380
rect 37280 39296 37332 39302
rect 37280 39238 37332 39244
rect 37292 39098 37320 39238
rect 37280 39092 37332 39098
rect 37280 39034 37332 39040
rect 37292 38962 37320 39034
rect 37280 38956 37332 38962
rect 37280 38898 37332 38904
rect 37476 38894 37504 39782
rect 37568 39438 37596 39986
rect 37556 39432 37608 39438
rect 37556 39374 37608 39380
rect 37464 38888 37516 38894
rect 37464 38830 37516 38836
rect 37476 38758 37504 38830
rect 37280 38752 37332 38758
rect 37280 38694 37332 38700
rect 37464 38752 37516 38758
rect 37464 38694 37516 38700
rect 37292 38350 37320 38694
rect 37188 38344 37240 38350
rect 37188 38286 37240 38292
rect 37280 38344 37332 38350
rect 37280 38286 37332 38292
rect 37200 38214 37228 38286
rect 37188 38208 37240 38214
rect 37188 38150 37240 38156
rect 37200 37398 37228 38150
rect 37292 37942 37320 38286
rect 37280 37936 37332 37942
rect 37660 37890 37688 40870
rect 37844 40662 37872 41074
rect 37832 40656 37884 40662
rect 37832 40598 37884 40604
rect 37280 37878 37332 37884
rect 37476 37862 37688 37890
rect 37740 37868 37792 37874
rect 37188 37392 37240 37398
rect 37188 37334 37240 37340
rect 37280 37256 37332 37262
rect 37280 37198 37332 37204
rect 37292 36922 37320 37198
rect 37372 37188 37424 37194
rect 37372 37130 37424 37136
rect 37280 36916 37332 36922
rect 37280 36858 37332 36864
rect 37384 36174 37412 37130
rect 37372 36168 37424 36174
rect 37372 36110 37424 36116
rect 37476 35850 37504 37862
rect 37740 37810 37792 37816
rect 37556 37732 37608 37738
rect 37556 37674 37608 37680
rect 37568 37398 37596 37674
rect 37556 37392 37608 37398
rect 37556 37334 37608 37340
rect 37648 37256 37700 37262
rect 37752 37244 37780 37810
rect 37700 37216 37780 37244
rect 37648 37198 37700 37204
rect 37648 36100 37700 36106
rect 37648 36042 37700 36048
rect 37384 35822 37504 35850
rect 37384 33454 37412 35822
rect 37660 35766 37688 36042
rect 37752 35834 37780 37216
rect 37832 36780 37884 36786
rect 37832 36722 37884 36728
rect 37844 36106 37872 36722
rect 37832 36100 37884 36106
rect 37832 36042 37884 36048
rect 37740 35828 37792 35834
rect 37740 35770 37792 35776
rect 37464 35760 37516 35766
rect 37464 35702 37516 35708
rect 37648 35760 37700 35766
rect 37648 35702 37700 35708
rect 37476 35290 37504 35702
rect 37740 35488 37792 35494
rect 37740 35430 37792 35436
rect 37464 35284 37516 35290
rect 37464 35226 37516 35232
rect 37648 35012 37700 35018
rect 37648 34954 37700 34960
rect 37660 34610 37688 34954
rect 37648 34604 37700 34610
rect 37648 34546 37700 34552
rect 37648 33856 37700 33862
rect 37648 33798 37700 33804
rect 37464 33516 37516 33522
rect 37464 33458 37516 33464
rect 37372 33448 37424 33454
rect 37372 33390 37424 33396
rect 37096 31952 37148 31958
rect 37096 31894 37148 31900
rect 37384 31822 37412 33390
rect 37476 32570 37504 33458
rect 37660 32978 37688 33798
rect 37648 32972 37700 32978
rect 37648 32914 37700 32920
rect 37464 32564 37516 32570
rect 37464 32506 37516 32512
rect 37476 31958 37504 32506
rect 37648 32360 37700 32366
rect 37648 32302 37700 32308
rect 37464 31952 37516 31958
rect 37464 31894 37516 31900
rect 37372 31816 37424 31822
rect 37372 31758 37424 31764
rect 37280 31680 37332 31686
rect 37280 31622 37332 31628
rect 37292 31414 37320 31622
rect 37280 31408 37332 31414
rect 37280 31350 37332 31356
rect 37384 30870 37412 31758
rect 37372 30864 37424 30870
rect 37372 30806 37424 30812
rect 37476 30734 37504 31894
rect 37660 31890 37688 32302
rect 37648 31884 37700 31890
rect 37648 31826 37700 31832
rect 37660 31482 37688 31826
rect 37648 31476 37700 31482
rect 37648 31418 37700 31424
rect 37464 30728 37516 30734
rect 37464 30670 37516 30676
rect 37556 27940 37608 27946
rect 37556 27882 37608 27888
rect 37568 27674 37596 27882
rect 37556 27668 37608 27674
rect 37556 27610 37608 27616
rect 37568 27334 37596 27610
rect 37556 27328 37608 27334
rect 37556 27270 37608 27276
rect 35900 2576 35952 2582
rect 35900 2518 35952 2524
rect 36912 2576 36964 2582
rect 36912 2518 36964 2524
rect 37752 2446 37780 35430
rect 37844 35086 37872 36042
rect 37832 35080 37884 35086
rect 37832 35022 37884 35028
rect 37936 31754 37964 43030
rect 38016 42288 38068 42294
rect 38016 42230 38068 42236
rect 38028 41274 38056 42230
rect 38120 42158 38148 45018
rect 38384 44260 38436 44266
rect 38384 44202 38436 44208
rect 38396 43110 38424 44202
rect 38660 43648 38712 43654
rect 38660 43590 38712 43596
rect 38384 43104 38436 43110
rect 38384 43046 38436 43052
rect 38396 42566 38424 43046
rect 38672 42770 38700 43590
rect 38660 42764 38712 42770
rect 38660 42706 38712 42712
rect 38384 42560 38436 42566
rect 38384 42502 38436 42508
rect 38396 42362 38424 42502
rect 38384 42356 38436 42362
rect 38384 42298 38436 42304
rect 38108 42152 38160 42158
rect 38108 42094 38160 42100
rect 38108 41608 38160 41614
rect 38108 41550 38160 41556
rect 38016 41268 38068 41274
rect 38016 41210 38068 41216
rect 38120 41138 38148 41550
rect 38200 41472 38252 41478
rect 38200 41414 38252 41420
rect 38108 41132 38160 41138
rect 38108 41074 38160 41080
rect 38120 40526 38148 41074
rect 38212 41070 38240 41414
rect 38660 41268 38712 41274
rect 38660 41210 38712 41216
rect 38672 41177 38700 41210
rect 38658 41168 38714 41177
rect 38658 41103 38660 41112
rect 38712 41103 38714 41112
rect 38660 41074 38712 41080
rect 38200 41064 38252 41070
rect 38200 41006 38252 41012
rect 38108 40520 38160 40526
rect 38108 40462 38160 40468
rect 38108 40384 38160 40390
rect 38108 40326 38160 40332
rect 38120 40050 38148 40326
rect 38108 40044 38160 40050
rect 38108 39986 38160 39992
rect 38212 39370 38240 41006
rect 38384 40656 38436 40662
rect 38384 40598 38436 40604
rect 38292 39908 38344 39914
rect 38292 39850 38344 39856
rect 38304 39506 38332 39850
rect 38292 39500 38344 39506
rect 38292 39442 38344 39448
rect 38200 39364 38252 39370
rect 38200 39306 38252 39312
rect 38396 39098 38424 40598
rect 38672 40526 38700 41074
rect 38660 40520 38712 40526
rect 38660 40462 38712 40468
rect 38476 40452 38528 40458
rect 38476 40394 38528 40400
rect 38488 39438 38516 40394
rect 38672 40118 38700 40462
rect 38660 40112 38712 40118
rect 38660 40054 38712 40060
rect 38660 39976 38712 39982
rect 38660 39918 38712 39924
rect 38568 39636 38620 39642
rect 38568 39578 38620 39584
rect 38476 39432 38528 39438
rect 38476 39374 38528 39380
rect 38580 39098 38608 39578
rect 38384 39092 38436 39098
rect 38384 39034 38436 39040
rect 38568 39092 38620 39098
rect 38568 39034 38620 39040
rect 38672 38962 38700 39918
rect 38384 38956 38436 38962
rect 38384 38898 38436 38904
rect 38660 38956 38712 38962
rect 38660 38898 38712 38904
rect 38396 38282 38424 38898
rect 38476 38344 38528 38350
rect 38474 38312 38476 38321
rect 38528 38312 38530 38321
rect 38384 38276 38436 38282
rect 38474 38247 38530 38256
rect 38384 38218 38436 38224
rect 38396 37670 38424 38218
rect 38672 38214 38700 38898
rect 38856 38826 38884 54470
rect 40144 54330 40172 54470
rect 40132 54324 40184 54330
rect 40132 54266 40184 54272
rect 42628 54058 42656 54470
rect 45112 54330 45140 54674
rect 48976 54670 49004 54810
rect 53484 54670 53512 56841
rect 53562 55176 53618 55185
rect 53562 55111 53618 55120
rect 45468 54664 45520 54670
rect 45468 54606 45520 54612
rect 47584 54664 47636 54670
rect 47584 54606 47636 54612
rect 48964 54664 49016 54670
rect 48964 54606 49016 54612
rect 51632 54664 51684 54670
rect 51632 54606 51684 54612
rect 53472 54664 53524 54670
rect 53472 54606 53524 54612
rect 45100 54324 45152 54330
rect 45100 54266 45152 54272
rect 42616 54052 42668 54058
rect 42616 53994 42668 54000
rect 45480 53174 45508 54606
rect 45468 53168 45520 53174
rect 45468 53110 45520 53116
rect 39120 44192 39172 44198
rect 39120 44134 39172 44140
rect 39132 43654 39160 44134
rect 39120 43648 39172 43654
rect 39120 43590 39172 43596
rect 38936 42696 38988 42702
rect 38936 42638 38988 42644
rect 38948 41818 38976 42638
rect 39132 42634 39160 43590
rect 39948 43172 40000 43178
rect 39948 43114 40000 43120
rect 39488 43104 39540 43110
rect 39488 43046 39540 43052
rect 39500 42838 39528 43046
rect 39488 42832 39540 42838
rect 39488 42774 39540 42780
rect 39120 42628 39172 42634
rect 39120 42570 39172 42576
rect 39028 42016 39080 42022
rect 39028 41958 39080 41964
rect 38936 41812 38988 41818
rect 38936 41754 38988 41760
rect 39040 41614 39068 41958
rect 39132 41614 39160 42570
rect 39960 42566 39988 43114
rect 40500 43104 40552 43110
rect 40500 43046 40552 43052
rect 40040 42764 40092 42770
rect 40040 42706 40092 42712
rect 39948 42560 40000 42566
rect 39948 42502 40000 42508
rect 39028 41608 39080 41614
rect 39028 41550 39080 41556
rect 39120 41608 39172 41614
rect 39120 41550 39172 41556
rect 39212 41132 39264 41138
rect 39212 41074 39264 41080
rect 39396 41132 39448 41138
rect 39396 41074 39448 41080
rect 39224 40526 39252 41074
rect 39212 40520 39264 40526
rect 39212 40462 39264 40468
rect 39408 40186 39436 41074
rect 39672 40452 39724 40458
rect 39672 40394 39724 40400
rect 39396 40180 39448 40186
rect 39396 40122 39448 40128
rect 39684 40050 39712 40394
rect 38936 40044 38988 40050
rect 38936 39986 38988 39992
rect 39672 40044 39724 40050
rect 39672 39986 39724 39992
rect 39856 40044 39908 40050
rect 39856 39986 39908 39992
rect 38948 38894 38976 39986
rect 39028 39296 39080 39302
rect 39028 39238 39080 39244
rect 38936 38888 38988 38894
rect 38936 38830 38988 38836
rect 38844 38820 38896 38826
rect 38844 38762 38896 38768
rect 38660 38208 38712 38214
rect 38660 38150 38712 38156
rect 38384 37664 38436 37670
rect 38384 37606 38436 37612
rect 38200 37460 38252 37466
rect 38200 37402 38252 37408
rect 38016 37188 38068 37194
rect 38016 37130 38068 37136
rect 38028 36718 38056 37130
rect 38212 36922 38240 37402
rect 38396 37194 38424 37606
rect 38672 37466 38700 38150
rect 38752 37868 38804 37874
rect 38752 37810 38804 37816
rect 38660 37460 38712 37466
rect 38660 37402 38712 37408
rect 38672 37244 38700 37402
rect 38580 37216 38700 37244
rect 38384 37188 38436 37194
rect 38384 37130 38436 37136
rect 38292 37120 38344 37126
rect 38292 37062 38344 37068
rect 38200 36916 38252 36922
rect 38200 36858 38252 36864
rect 38016 36712 38068 36718
rect 38016 36654 38068 36660
rect 38304 36242 38332 37062
rect 38292 36236 38344 36242
rect 38292 36178 38344 36184
rect 38292 35692 38344 35698
rect 38292 35634 38344 35640
rect 38304 34746 38332 35634
rect 38396 35494 38424 37130
rect 38580 35766 38608 37216
rect 38764 36786 38792 37810
rect 38752 36780 38804 36786
rect 38752 36722 38804 36728
rect 38764 36378 38792 36722
rect 39040 36718 39068 39238
rect 39028 36712 39080 36718
rect 39028 36654 39080 36660
rect 38752 36372 38804 36378
rect 38752 36314 38804 36320
rect 39040 36310 39068 36654
rect 39028 36304 39080 36310
rect 39028 36246 39080 36252
rect 38752 36168 38804 36174
rect 38752 36110 38804 36116
rect 38568 35760 38620 35766
rect 38568 35702 38620 35708
rect 38764 35698 38792 36110
rect 39684 35834 39712 39986
rect 39868 39914 39896 39986
rect 39856 39908 39908 39914
rect 39856 39850 39908 39856
rect 39868 39370 39896 39850
rect 39856 39364 39908 39370
rect 39856 39306 39908 39312
rect 39868 38214 39896 39306
rect 39856 38208 39908 38214
rect 39856 38150 39908 38156
rect 39764 36100 39816 36106
rect 39764 36042 39816 36048
rect 39672 35828 39724 35834
rect 39672 35770 39724 35776
rect 38752 35692 38804 35698
rect 38752 35634 38804 35640
rect 38384 35488 38436 35494
rect 38384 35430 38436 35436
rect 38292 34740 38344 34746
rect 38292 34682 38344 34688
rect 38016 34400 38068 34406
rect 38016 34342 38068 34348
rect 38028 33930 38056 34342
rect 38016 33924 38068 33930
rect 38016 33866 38068 33872
rect 38028 33046 38056 33866
rect 38200 33856 38252 33862
rect 38200 33798 38252 33804
rect 38212 33590 38240 33798
rect 38200 33584 38252 33590
rect 38200 33526 38252 33532
rect 38016 33040 38068 33046
rect 38016 32982 38068 32988
rect 38028 32842 38056 32982
rect 38016 32836 38068 32842
rect 38016 32778 38068 32784
rect 38212 32774 38240 33526
rect 38764 33454 38792 35634
rect 38844 34944 38896 34950
rect 38844 34886 38896 34892
rect 38856 34542 38884 34886
rect 39684 34746 39712 35770
rect 39776 35698 39804 36042
rect 39764 35692 39816 35698
rect 39764 35634 39816 35640
rect 39776 35290 39804 35634
rect 39764 35284 39816 35290
rect 39764 35226 39816 35232
rect 39672 34740 39724 34746
rect 39672 34682 39724 34688
rect 39684 34542 39712 34682
rect 38844 34536 38896 34542
rect 38844 34478 38896 34484
rect 39672 34536 39724 34542
rect 39672 34478 39724 34484
rect 38936 33992 38988 33998
rect 38936 33934 38988 33940
rect 38752 33448 38804 33454
rect 38752 33390 38804 33396
rect 38948 33114 38976 33934
rect 38292 33108 38344 33114
rect 38292 33050 38344 33056
rect 38936 33108 38988 33114
rect 38936 33050 38988 33056
rect 38200 32768 38252 32774
rect 38200 32710 38252 32716
rect 38212 32570 38240 32710
rect 38200 32564 38252 32570
rect 38200 32506 38252 32512
rect 38304 31754 38332 33050
rect 38660 32836 38712 32842
rect 38660 32778 38712 32784
rect 38672 32570 38700 32778
rect 38660 32564 38712 32570
rect 38660 32506 38712 32512
rect 37936 31726 38148 31754
rect 37832 28688 37884 28694
rect 37832 28630 37884 28636
rect 37844 28218 37872 28630
rect 37832 28212 37884 28218
rect 37832 28154 37884 28160
rect 38120 5098 38148 31726
rect 38212 31726 38332 31754
rect 38212 31142 38240 31726
rect 38200 31136 38252 31142
rect 38200 31078 38252 31084
rect 38212 30394 38240 31078
rect 38200 30388 38252 30394
rect 38200 30330 38252 30336
rect 39960 21418 39988 42502
rect 40052 41818 40080 42706
rect 40512 42362 40540 43046
rect 40960 42560 41012 42566
rect 40960 42502 41012 42508
rect 40500 42356 40552 42362
rect 40500 42298 40552 42304
rect 40972 42022 41000 42502
rect 40960 42016 41012 42022
rect 40960 41958 41012 41964
rect 40972 41818 41000 41958
rect 40040 41812 40092 41818
rect 40040 41754 40092 41760
rect 40408 41812 40460 41818
rect 40408 41754 40460 41760
rect 40960 41812 41012 41818
rect 40960 41754 41012 41760
rect 40040 41676 40092 41682
rect 40040 41618 40092 41624
rect 40052 40526 40080 41618
rect 40420 40934 40448 41754
rect 42064 41472 42116 41478
rect 42064 41414 42116 41420
rect 41052 41268 41104 41274
rect 41052 41210 41104 41216
rect 40408 40928 40460 40934
rect 40408 40870 40460 40876
rect 40040 40520 40092 40526
rect 40040 40462 40092 40468
rect 40420 40390 40448 40870
rect 41064 40730 41092 41210
rect 41512 40928 41564 40934
rect 41512 40870 41564 40876
rect 41052 40724 41104 40730
rect 41052 40666 41104 40672
rect 41524 40458 41552 40870
rect 41512 40452 41564 40458
rect 41512 40394 41564 40400
rect 40408 40384 40460 40390
rect 40408 40326 40460 40332
rect 40420 40186 40448 40326
rect 40040 40180 40092 40186
rect 40040 40122 40092 40128
rect 40408 40180 40460 40186
rect 40408 40122 40460 40128
rect 41052 40180 41104 40186
rect 41052 40122 41104 40128
rect 40052 39574 40080 40122
rect 41064 39982 41092 40122
rect 41052 39976 41104 39982
rect 41052 39918 41104 39924
rect 41524 39642 41552 40394
rect 41512 39636 41564 39642
rect 41512 39578 41564 39584
rect 40040 39568 40092 39574
rect 40040 39510 40092 39516
rect 40052 39098 40080 39510
rect 40408 39296 40460 39302
rect 40408 39238 40460 39244
rect 40040 39092 40092 39098
rect 40040 39034 40092 39040
rect 40420 38758 40448 39238
rect 40040 38752 40092 38758
rect 40040 38694 40092 38700
rect 40408 38752 40460 38758
rect 40408 38694 40460 38700
rect 40052 38282 40080 38694
rect 40040 38276 40092 38282
rect 40040 38218 40092 38224
rect 40408 33856 40460 33862
rect 40408 33798 40460 33804
rect 40420 33386 40448 33798
rect 40408 33380 40460 33386
rect 40408 33322 40460 33328
rect 40420 32774 40448 33322
rect 40408 32768 40460 32774
rect 40408 32710 40460 32716
rect 39948 21412 40000 21418
rect 39948 21354 40000 21360
rect 40420 9926 40448 32710
rect 41512 27328 41564 27334
rect 41512 27270 41564 27276
rect 40408 9920 40460 9926
rect 40408 9862 40460 9868
rect 38108 5092 38160 5098
rect 38108 5034 38160 5040
rect 41524 2582 41552 27270
rect 42076 13870 42104 41414
rect 47596 30326 47624 54606
rect 49148 54528 49200 54534
rect 49148 54470 49200 54476
rect 49160 40633 49188 54470
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 51644 43450 51672 54606
rect 53576 54262 53604 55111
rect 53656 54528 53708 54534
rect 53656 54470 53708 54476
rect 53564 54256 53616 54262
rect 53564 54198 53616 54204
rect 53380 54052 53432 54058
rect 53380 53994 53432 54000
rect 52460 53440 52512 53446
rect 52460 53382 52512 53388
rect 52472 49978 52500 53382
rect 53288 52896 53340 52902
rect 53288 52838 53340 52844
rect 52460 49972 52512 49978
rect 52460 49914 52512 49920
rect 53104 48612 53156 48618
rect 53104 48554 53156 48560
rect 52368 43648 52420 43654
rect 52368 43590 52420 43596
rect 51632 43444 51684 43450
rect 51632 43386 51684 43392
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 49146 40624 49202 40633
rect 49146 40559 49202 40568
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 52380 36038 52408 43590
rect 52828 39908 52880 39914
rect 52828 39850 52880 39856
rect 52840 37466 52868 39850
rect 52828 37460 52880 37466
rect 52828 37402 52880 37408
rect 52840 37262 52868 37402
rect 52828 37256 52880 37262
rect 52828 37198 52880 37204
rect 52368 36032 52420 36038
rect 52368 35974 52420 35980
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 52460 34944 52512 34950
rect 52460 34886 52512 34892
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 50712 34536 50764 34542
rect 50712 34478 50764 34484
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 47584 30320 47636 30326
rect 47584 30262 47636 30268
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 42064 13864 42116 13870
rect 42064 13806 42116 13812
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 45100 2848 45152 2854
rect 45100 2790 45152 2796
rect 47676 2848 47728 2854
rect 47676 2790 47728 2796
rect 50344 2848 50396 2854
rect 50344 2790 50396 2796
rect 41512 2576 41564 2582
rect 41512 2518 41564 2524
rect 45112 2446 45140 2790
rect 35348 2440 35400 2446
rect 35348 2382 35400 2388
rect 37740 2440 37792 2446
rect 37740 2382 37792 2388
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 45100 2440 45152 2446
rect 45100 2382 45152 2388
rect 45374 2408 45430 2417
rect 34520 2372 34572 2378
rect 34440 2332 34520 2360
rect 34164 870 34284 898
rect 34164 800 34192 870
rect 18 0 74 800
rect 1950 0 2006 800
rect 3882 0 3938 800
rect 6458 0 6514 800
rect 8390 0 8446 800
rect 10322 0 10378 800
rect 12898 0 12954 800
rect 14830 0 14886 800
rect 16762 0 16818 800
rect 19338 0 19394 800
rect 21270 0 21326 800
rect 23846 0 23902 800
rect 25778 0 25834 800
rect 27710 0 27766 800
rect 30286 0 30342 800
rect 32218 0 32274 800
rect 34150 0 34206 800
rect 34256 762 34284 870
rect 34440 762 34468 2332
rect 34520 2314 34572 2320
rect 36728 2304 36780 2310
rect 36728 2246 36780 2252
rect 36740 800 36768 2246
rect 38672 800 38700 2382
rect 41236 2372 41288 2378
rect 41236 2314 41288 2320
rect 41248 800 41276 2314
rect 42800 2304 42852 2310
rect 42800 2246 42852 2252
rect 43168 2304 43220 2310
rect 43168 2246 43220 2252
rect 42812 2038 42840 2246
rect 42800 2032 42852 2038
rect 42800 1974 42852 1980
rect 43180 800 43208 2246
rect 45112 800 45140 2382
rect 47688 2378 47716 2790
rect 50356 2446 50384 2790
rect 50724 2650 50752 34478
rect 51724 31816 51776 31822
rect 51724 31758 51776 31764
rect 51448 25492 51500 25498
rect 51448 25434 51500 25440
rect 51460 3194 51488 25434
rect 51736 23866 51764 31758
rect 52472 26314 52500 34886
rect 53116 33318 53144 48554
rect 53300 34649 53328 52838
rect 53392 50250 53420 53994
rect 53564 53508 53616 53514
rect 53564 53450 53616 53456
rect 53576 53145 53604 53450
rect 53562 53136 53618 53145
rect 53562 53071 53618 53080
rect 53564 50924 53616 50930
rect 53564 50866 53616 50872
rect 53472 50720 53524 50726
rect 53472 50662 53524 50668
rect 53484 50522 53512 50662
rect 53472 50516 53524 50522
rect 53472 50458 53524 50464
rect 53576 50425 53604 50866
rect 53562 50416 53618 50425
rect 53562 50351 53618 50360
rect 53380 50244 53432 50250
rect 53380 50186 53432 50192
rect 53564 48748 53616 48754
rect 53564 48690 53616 48696
rect 53576 48385 53604 48690
rect 53562 48376 53618 48385
rect 53562 48311 53618 48320
rect 53564 46368 53616 46374
rect 53562 46336 53564 46345
rect 53616 46336 53618 46345
rect 53562 46271 53618 46280
rect 53564 43648 53616 43654
rect 53562 43616 53564 43625
rect 53616 43616 53618 43625
rect 53562 43551 53618 43560
rect 53378 41576 53434 41585
rect 53378 41511 53380 41520
rect 53432 41511 53434 41520
rect 53562 41576 53618 41585
rect 53562 41511 53564 41520
rect 53380 41482 53432 41488
rect 53616 41511 53618 41520
rect 53564 41482 53616 41488
rect 53564 40044 53616 40050
rect 53564 39986 53616 39992
rect 53576 39545 53604 39986
rect 53562 39536 53618 39545
rect 53562 39471 53618 39480
rect 53564 37120 53616 37126
rect 53564 37062 53616 37068
rect 53576 36825 53604 37062
rect 53562 36816 53618 36825
rect 53562 36751 53618 36760
rect 53564 35012 53616 35018
rect 53564 34954 53616 34960
rect 53576 34785 53604 34954
rect 53562 34776 53618 34785
rect 53562 34711 53618 34720
rect 53286 34640 53342 34649
rect 53286 34575 53342 34584
rect 53668 33998 53696 54470
rect 55416 53106 55444 56841
rect 55404 53100 55456 53106
rect 55404 53042 55456 53048
rect 53656 33992 53708 33998
rect 53656 33934 53708 33940
rect 53104 33312 53156 33318
rect 53104 33254 53156 33260
rect 53564 32428 53616 32434
rect 53564 32370 53616 32376
rect 53380 32292 53432 32298
rect 53380 32234 53432 32240
rect 53392 29306 53420 32234
rect 53576 32065 53604 32370
rect 53562 32056 53618 32065
rect 53562 31991 53618 32000
rect 53564 30252 53616 30258
rect 53564 30194 53616 30200
rect 53472 30048 53524 30054
rect 53576 30025 53604 30194
rect 53472 29990 53524 29996
rect 53562 30016 53618 30025
rect 53484 29782 53512 29990
rect 53562 29951 53618 29960
rect 53472 29776 53524 29782
rect 53472 29718 53524 29724
rect 53380 29300 53432 29306
rect 53380 29242 53432 29248
rect 53380 28008 53432 28014
rect 53656 28008 53708 28014
rect 53380 27950 53432 27956
rect 53654 27976 53656 27985
rect 53708 27976 53710 27985
rect 52828 26444 52880 26450
rect 52828 26386 52880 26392
rect 52460 26308 52512 26314
rect 52460 26250 52512 26256
rect 52840 25498 52868 26386
rect 53392 26382 53420 27950
rect 53654 27911 53710 27920
rect 53668 27674 53696 27911
rect 53656 27668 53708 27674
rect 53656 27610 53708 27616
rect 53380 26376 53432 26382
rect 53380 26318 53432 26324
rect 52828 25492 52880 25498
rect 52828 25434 52880 25440
rect 52840 25294 52868 25434
rect 52828 25288 52880 25294
rect 52828 25230 52880 25236
rect 53562 25256 53618 25265
rect 53562 25191 53618 25200
rect 53576 25158 53604 25191
rect 53564 25152 53616 25158
rect 53564 25094 53616 25100
rect 51724 23860 51776 23866
rect 51724 23802 51776 23808
rect 53564 23520 53616 23526
rect 53564 23462 53616 23468
rect 53576 23225 53604 23462
rect 53562 23216 53618 23225
rect 53562 23151 53618 23160
rect 53564 21344 53616 21350
rect 53564 21286 53616 21292
rect 53576 21185 53604 21286
rect 53562 21176 53618 21185
rect 53562 21111 53618 21120
rect 53564 18692 53616 18698
rect 53564 18634 53616 18640
rect 53576 18465 53604 18634
rect 53562 18456 53618 18465
rect 53562 18391 53618 18400
rect 53564 16448 53616 16454
rect 53562 16416 53564 16425
rect 53616 16416 53618 16425
rect 53562 16351 53618 16360
rect 53656 13932 53708 13938
rect 53656 13874 53708 13880
rect 53668 13705 53696 13874
rect 53654 13696 53710 13705
rect 53654 13631 53710 13640
rect 53562 11656 53618 11665
rect 53562 11591 53564 11600
rect 53616 11591 53618 11600
rect 53564 11562 53616 11568
rect 53564 9988 53616 9994
rect 53564 9930 53616 9936
rect 53576 9625 53604 9930
rect 53562 9616 53618 9625
rect 53562 9551 53618 9560
rect 53656 7404 53708 7410
rect 53656 7346 53708 7352
rect 53668 6905 53696 7346
rect 53654 6896 53710 6905
rect 53654 6831 53710 6840
rect 53564 5024 53616 5030
rect 53564 4966 53616 4972
rect 53576 4865 53604 4966
rect 53562 4856 53618 4865
rect 53562 4791 53618 4800
rect 54116 3392 54168 3398
rect 54116 3334 54168 3340
rect 51448 3188 51500 3194
rect 51448 3130 51500 3136
rect 50712 2644 50764 2650
rect 50712 2586 50764 2592
rect 51460 2446 51488 3130
rect 52460 2848 52512 2854
rect 53564 2848 53616 2854
rect 52460 2790 52512 2796
rect 53562 2816 53564 2825
rect 53616 2816 53618 2825
rect 49700 2440 49752 2446
rect 49620 2400 49700 2428
rect 45374 2343 45430 2352
rect 47676 2372 47728 2378
rect 45388 2310 45416 2343
rect 47676 2314 47728 2320
rect 45376 2304 45428 2310
rect 45376 2246 45428 2252
rect 47688 800 47716 2314
rect 48136 2304 48188 2310
rect 48136 2246 48188 2252
rect 48148 1902 48176 2246
rect 48136 1896 48188 1902
rect 48136 1838 48188 1844
rect 49620 800 49648 2400
rect 49700 2382 49752 2388
rect 50344 2440 50396 2446
rect 50344 2382 50396 2388
rect 51448 2440 51500 2446
rect 51448 2382 51500 2388
rect 52472 2378 52500 2790
rect 53562 2751 53618 2760
rect 52460 2372 52512 2378
rect 52460 2314 52512 2320
rect 53564 2372 53616 2378
rect 53564 2314 53616 2320
rect 51540 2304 51592 2310
rect 51540 2246 51592 2252
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 51552 800 51580 2246
rect 34256 734 34468 762
rect 36726 0 36782 800
rect 38658 0 38714 800
rect 41234 0 41290 800
rect 43166 0 43222 800
rect 45098 0 45154 800
rect 47674 0 47730 800
rect 49606 0 49662 800
rect 51538 0 51594 800
rect 53576 105 53604 2314
rect 54128 800 54156 3334
rect 53562 96 53618 105
rect 53562 31 53618 40
rect 54114 0 54170 800
<< via2 >>
rect 1582 57160 1638 57216
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 1398 52436 1400 52456
rect 1400 52436 1452 52456
rect 1452 52436 1454 52456
rect 1398 52400 1454 52436
rect 1398 50396 1400 50416
rect 1400 50396 1452 50416
rect 1452 50396 1454 50416
rect 1398 50360 1454 50396
rect 1490 47640 1546 47696
rect 1582 45620 1638 45656
rect 1582 45600 1584 45620
rect 1584 45600 1636 45620
rect 1636 45600 1638 45620
rect 2778 54440 2834 54496
rect 1582 43560 1638 43616
rect 1766 42744 1822 42800
rect 1490 40876 1492 40896
rect 1492 40876 1544 40896
rect 1544 40876 1546 40896
rect 1490 40840 1546 40876
rect 1582 38800 1638 38856
rect 1858 36100 1914 36136
rect 1858 36080 1860 36100
rect 1860 36080 1912 36100
rect 1912 36080 1914 36100
rect 2226 48068 2282 48104
rect 2226 48048 2228 48068
rect 2228 48048 2280 48068
rect 2280 48048 2282 48068
rect 1950 35128 2006 35184
rect 1582 34076 1584 34096
rect 1584 34076 1636 34096
rect 1636 34076 1638 34096
rect 1582 34040 1638 34076
rect 1490 32000 1546 32056
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 8022 41112 8078 41168
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 1398 29300 1454 29336
rect 1398 29280 1400 29300
rect 1400 29280 1452 29300
rect 1452 29280 1454 29300
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 1490 27276 1492 27296
rect 1492 27276 1544 27296
rect 1544 27276 1546 27296
rect 1490 27240 1546 27276
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 1858 25220 1914 25256
rect 1858 25200 1860 25220
rect 1860 25200 1912 25220
rect 1912 25200 1914 25220
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 1398 22480 1454 22536
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 1582 20848 1638 20904
rect 1398 20476 1400 20496
rect 1400 20476 1452 20496
rect 1452 20476 1454 20496
rect 1398 20440 1454 20476
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 1582 17756 1584 17776
rect 1584 17756 1636 17776
rect 1636 17756 1638 17776
rect 1582 17720 1638 17756
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 1398 15700 1454 15736
rect 1398 15680 1400 15700
rect 1400 15680 1452 15700
rect 1452 15680 1454 15700
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 1490 13676 1492 13696
rect 1492 13676 1544 13696
rect 1544 13676 1546 13696
rect 1490 13640 1546 13676
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 1582 10920 1638 10976
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 1490 8880 1546 8936
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 1582 6840 1638 6896
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 1490 4120 1546 4176
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 1858 2080 1914 2136
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 9126 2352 9182 2408
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 21638 49680 21694 49736
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 20718 47404 20720 47424
rect 20720 47404 20772 47424
rect 20772 47404 20774 47424
rect 20718 47368 20774 47404
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 18786 40996 18842 41032
rect 18786 40976 18788 40996
rect 18788 40976 18840 40996
rect 18840 40976 18842 40996
rect 18234 34604 18290 34640
rect 18234 34584 18236 34604
rect 18236 34584 18288 34604
rect 18288 34584 18290 34604
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19982 40568 20038 40624
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 21638 41692 21640 41712
rect 21640 41692 21692 41712
rect 21692 41692 21694 41712
rect 21638 41656 21694 41692
rect 23570 48456 23626 48512
rect 23846 41540 23902 41576
rect 23846 41520 23848 41540
rect 23848 41520 23900 41540
rect 23900 41520 23902 41540
rect 21914 38664 21970 38720
rect 22558 38664 22614 38720
rect 24398 41520 24454 41576
rect 29458 48048 29514 48104
rect 27066 41656 27122 41712
rect 27342 41384 27398 41440
rect 24582 2524 24584 2544
rect 24584 2524 24636 2544
rect 24636 2524 24638 2544
rect 24582 2488 24638 2524
rect 28906 40704 28962 40760
rect 28722 33224 28778 33280
rect 29366 33396 29368 33416
rect 29368 33396 29420 33416
rect 29420 33396 29422 33416
rect 29366 33360 29422 33396
rect 29826 41384 29882 41440
rect 29550 41248 29606 41304
rect 29550 39092 29606 39128
rect 29550 39072 29552 39092
rect 29552 39072 29604 39092
rect 29604 39072 29606 39092
rect 30930 46980 30986 47016
rect 30930 46960 30932 46980
rect 30932 46960 30984 46980
rect 30984 46960 30986 46980
rect 29826 33224 29882 33280
rect 30746 40976 30802 41032
rect 32034 47504 32090 47560
rect 32034 46960 32090 47016
rect 31758 46688 31814 46744
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 33598 47096 33654 47152
rect 33230 46980 33286 47016
rect 33230 46960 33232 46980
rect 33232 46960 33284 46980
rect 33284 46960 33286 46980
rect 30562 38392 30618 38448
rect 30746 38392 30802 38448
rect 30562 34992 30618 35048
rect 30102 33396 30104 33416
rect 30104 33396 30156 33416
rect 30156 33396 30158 33416
rect 30102 33360 30158 33396
rect 30102 32444 30104 32464
rect 30104 32444 30156 32464
rect 30156 32444 30158 32464
rect 30102 32408 30158 32444
rect 32586 41248 32642 41304
rect 31574 39072 31630 39128
rect 30930 33224 30986 33280
rect 30838 32444 30840 32464
rect 30840 32444 30892 32464
rect 30892 32444 30894 32464
rect 30838 32408 30894 32444
rect 30746 28736 30802 28792
rect 33874 45892 33930 45928
rect 33874 45872 33876 45892
rect 33876 45872 33928 45892
rect 33928 45872 33930 45892
rect 34058 46708 34114 46744
rect 34058 46688 34060 46708
rect 34060 46688 34112 46708
rect 34112 46688 34114 46708
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34610 45908 34612 45928
rect 34612 45908 34664 45928
rect 34664 45908 34666 45928
rect 34610 45872 34666 45908
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 35346 47524 35402 47560
rect 35346 47504 35348 47524
rect 35348 47504 35400 47524
rect 35400 47504 35402 47524
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 33782 40704 33838 40760
rect 32494 33224 32550 33280
rect 33414 38292 33416 38312
rect 33416 38292 33468 38312
rect 33468 38292 33470 38312
rect 33414 38256 33470 38292
rect 34242 36216 34298 36272
rect 33966 28736 34022 28792
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34610 35028 34612 35048
rect 34612 35028 34664 35048
rect 34664 35028 34666 35048
rect 34610 34992 34666 35028
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 35070 36216 35126 36272
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 35346 35128 35402 35184
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35898 42744 35954 42800
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34978 28500 34980 28520
rect 34980 28500 35032 28520
rect 35032 28500 35034 28520
rect 34978 28464 35034 28500
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 36450 28464 36506 28520
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 37462 46960 37518 47016
rect 37002 42744 37058 42800
rect 38658 41132 38714 41168
rect 38658 41112 38660 41132
rect 38660 41112 38712 41132
rect 38712 41112 38714 41132
rect 38474 38292 38476 38312
rect 38476 38292 38528 38312
rect 38528 38292 38530 38312
rect 38474 38256 38530 38292
rect 53562 55120 53618 55176
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 49146 40568 49202 40624
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 45374 2352 45430 2408
rect 53562 53080 53618 53136
rect 53562 50360 53618 50416
rect 53562 48320 53618 48376
rect 53562 46316 53564 46336
rect 53564 46316 53616 46336
rect 53616 46316 53618 46336
rect 53562 46280 53618 46316
rect 53562 43596 53564 43616
rect 53564 43596 53616 43616
rect 53616 43596 53618 43616
rect 53562 43560 53618 43596
rect 53378 41540 53434 41576
rect 53378 41520 53380 41540
rect 53380 41520 53432 41540
rect 53432 41520 53434 41540
rect 53562 41540 53618 41576
rect 53562 41520 53564 41540
rect 53564 41520 53616 41540
rect 53616 41520 53618 41540
rect 53562 39480 53618 39536
rect 53562 36760 53618 36816
rect 53562 34720 53618 34776
rect 53286 34584 53342 34640
rect 53562 32000 53618 32056
rect 53562 29960 53618 30016
rect 53654 27956 53656 27976
rect 53656 27956 53708 27976
rect 53708 27956 53710 27976
rect 53654 27920 53710 27956
rect 53562 25200 53618 25256
rect 53562 23160 53618 23216
rect 53562 21120 53618 21176
rect 53562 18400 53618 18456
rect 53562 16396 53564 16416
rect 53564 16396 53616 16416
rect 53616 16396 53618 16416
rect 53562 16360 53618 16396
rect 53654 13640 53710 13696
rect 53562 11620 53618 11656
rect 53562 11600 53564 11620
rect 53564 11600 53616 11620
rect 53616 11600 53618 11620
rect 53562 9560 53618 9616
rect 53654 6840 53710 6896
rect 53562 4800 53618 4856
rect 53562 2796 53564 2816
rect 53564 2796 53616 2816
rect 53616 2796 53618 2816
rect 53562 2760 53618 2796
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 53562 40 53618 96
<< metal3 >>
rect 0 57218 800 57248
rect 1577 57218 1643 57221
rect 0 57216 1643 57218
rect 0 57160 1582 57216
rect 1638 57160 1643 57216
rect 0 57158 1643 57160
rect 0 57128 800 57158
rect 1577 57155 1643 57158
rect 53557 55178 53623 55181
rect 54697 55178 55497 55208
rect 53557 55176 55497 55178
rect 53557 55120 53562 55176
rect 53618 55120 55497 55176
rect 53557 55118 55497 55120
rect 53557 55115 53623 55118
rect 54697 55088 55497 55118
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 0 54498 800 54528
rect 2773 54498 2839 54501
rect 0 54496 2839 54498
rect 0 54440 2778 54496
rect 2834 54440 2839 54496
rect 0 54438 2839 54440
rect 0 54408 800 54438
rect 2773 54435 2839 54438
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 53557 53138 53623 53141
rect 54697 53138 55497 53168
rect 53557 53136 55497 53138
rect 53557 53080 53562 53136
rect 53618 53080 55497 53136
rect 53557 53078 55497 53080
rect 53557 53075 53623 53078
rect 54697 53048 55497 53078
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 0 52458 800 52488
rect 1393 52458 1459 52461
rect 0 52456 1459 52458
rect 0 52400 1398 52456
rect 1454 52400 1459 52456
rect 0 52398 1459 52400
rect 0 52368 800 52398
rect 1393 52395 1459 52398
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 0 50418 800 50448
rect 1393 50418 1459 50421
rect 0 50416 1459 50418
rect 0 50360 1398 50416
rect 1454 50360 1459 50416
rect 0 50358 1459 50360
rect 0 50328 800 50358
rect 1393 50355 1459 50358
rect 53557 50418 53623 50421
rect 54697 50418 55497 50448
rect 53557 50416 55497 50418
rect 53557 50360 53562 50416
rect 53618 50360 55497 50416
rect 53557 50358 55497 50360
rect 53557 50355 53623 50358
rect 54697 50328 55497 50358
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 21398 49676 21404 49740
rect 21468 49738 21474 49740
rect 21633 49738 21699 49741
rect 21468 49736 21699 49738
rect 21468 49680 21638 49736
rect 21694 49680 21699 49736
rect 21468 49678 21699 49680
rect 21468 49676 21474 49678
rect 21633 49675 21699 49678
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 23565 48514 23631 48517
rect 23790 48514 23796 48516
rect 23565 48512 23796 48514
rect 23565 48456 23570 48512
rect 23626 48456 23796 48512
rect 23565 48454 23796 48456
rect 23565 48451 23631 48454
rect 23790 48452 23796 48454
rect 23860 48452 23866 48516
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 53557 48378 53623 48381
rect 54697 48378 55497 48408
rect 53557 48376 55497 48378
rect 53557 48320 53562 48376
rect 53618 48320 55497 48376
rect 53557 48318 55497 48320
rect 53557 48315 53623 48318
rect 54697 48288 55497 48318
rect 2221 48106 2287 48109
rect 29453 48106 29519 48109
rect 2221 48104 29519 48106
rect 2221 48048 2226 48104
rect 2282 48048 29458 48104
rect 29514 48048 29519 48104
rect 2221 48046 29519 48048
rect 2221 48043 2287 48046
rect 29453 48043 29519 48046
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 0 47698 800 47728
rect 1485 47698 1551 47701
rect 0 47696 1551 47698
rect 0 47640 1490 47696
rect 1546 47640 1551 47696
rect 0 47638 1551 47640
rect 0 47608 800 47638
rect 1485 47635 1551 47638
rect 32029 47562 32095 47565
rect 35341 47562 35407 47565
rect 32029 47560 35407 47562
rect 32029 47504 32034 47560
rect 32090 47504 35346 47560
rect 35402 47504 35407 47560
rect 32029 47502 35407 47504
rect 32029 47499 32095 47502
rect 35341 47499 35407 47502
rect 20713 47428 20779 47429
rect 20662 47364 20668 47428
rect 20732 47426 20779 47428
rect 20732 47424 20824 47426
rect 20774 47368 20824 47424
rect 20732 47366 20824 47368
rect 20732 47364 20779 47366
rect 20713 47363 20779 47364
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 33593 47154 33659 47157
rect 33550 47152 33659 47154
rect 33550 47096 33598 47152
rect 33654 47096 33659 47152
rect 33550 47091 33659 47096
rect 30925 47020 30991 47021
rect 30925 47018 30972 47020
rect 30844 47016 30972 47018
rect 31036 47018 31042 47020
rect 32029 47018 32095 47021
rect 31036 47016 32095 47018
rect 30844 46960 30930 47016
rect 31036 46960 32034 47016
rect 32090 46960 32095 47016
rect 30844 46958 30972 46960
rect 30925 46956 30972 46958
rect 31036 46958 32095 46960
rect 31036 46956 31042 46958
rect 30925 46955 30991 46956
rect 32029 46955 32095 46958
rect 33225 47018 33291 47021
rect 33550 47018 33610 47091
rect 37457 47018 37523 47021
rect 33225 47016 37523 47018
rect 33225 46960 33230 47016
rect 33286 46960 37462 47016
rect 37518 46960 37523 47016
rect 33225 46958 37523 46960
rect 33225 46955 33291 46958
rect 37457 46955 37523 46958
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 31753 46746 31819 46749
rect 34053 46746 34119 46749
rect 31753 46744 34119 46746
rect 31753 46688 31758 46744
rect 31814 46688 34058 46744
rect 34114 46688 34119 46744
rect 31753 46686 34119 46688
rect 31753 46683 31819 46686
rect 34053 46683 34119 46686
rect 53557 46338 53623 46341
rect 54697 46338 55497 46368
rect 53557 46336 55497 46338
rect 53557 46280 53562 46336
rect 53618 46280 55497 46336
rect 53557 46278 55497 46280
rect 53557 46275 53623 46278
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 54697 46248 55497 46278
rect 34930 46207 35246 46208
rect 33869 45930 33935 45933
rect 34605 45930 34671 45933
rect 33869 45928 34671 45930
rect 33869 45872 33874 45928
rect 33930 45872 34610 45928
rect 34666 45872 34671 45928
rect 33869 45870 34671 45872
rect 33869 45867 33935 45870
rect 34605 45867 34671 45870
rect 19570 45728 19886 45729
rect 0 45658 800 45688
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 1577 45658 1643 45661
rect 0 45656 1643 45658
rect 0 45600 1582 45656
rect 1638 45600 1643 45656
rect 0 45598 1643 45600
rect 0 45568 800 45598
rect 1577 45595 1643 45598
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 0 43618 800 43648
rect 1577 43618 1643 43621
rect 0 43616 1643 43618
rect 0 43560 1582 43616
rect 1638 43560 1643 43616
rect 0 43558 1643 43560
rect 0 43528 800 43558
rect 1577 43555 1643 43558
rect 53557 43618 53623 43621
rect 54697 43618 55497 43648
rect 53557 43616 55497 43618
rect 53557 43560 53562 43616
rect 53618 43560 55497 43616
rect 53557 43558 55497 43560
rect 53557 43555 53623 43558
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 54697 43528 55497 43558
rect 50290 43487 50606 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 1761 42802 1827 42805
rect 35893 42802 35959 42805
rect 36997 42802 37063 42805
rect 1761 42800 37063 42802
rect 1761 42744 1766 42800
rect 1822 42744 35898 42800
rect 35954 42744 37002 42800
rect 37058 42744 37063 42800
rect 1761 42742 37063 42744
rect 1761 42739 1827 42742
rect 35893 42739 35959 42742
rect 36997 42739 37063 42742
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 21633 41714 21699 41717
rect 27061 41714 27127 41717
rect 21633 41712 27127 41714
rect 21633 41656 21638 41712
rect 21694 41656 27066 41712
rect 27122 41656 27127 41712
rect 21633 41654 27127 41656
rect 21633 41651 21699 41654
rect 27061 41651 27127 41654
rect 23841 41578 23907 41581
rect 24393 41578 24459 41581
rect 53373 41578 53439 41581
rect 23841 41576 53439 41578
rect 23841 41520 23846 41576
rect 23902 41520 24398 41576
rect 24454 41520 53378 41576
rect 53434 41520 53439 41576
rect 23841 41518 53439 41520
rect 23841 41515 23907 41518
rect 24393 41515 24459 41518
rect 53373 41515 53439 41518
rect 53557 41578 53623 41581
rect 54697 41578 55497 41608
rect 53557 41576 55497 41578
rect 53557 41520 53562 41576
rect 53618 41520 55497 41576
rect 53557 41518 55497 41520
rect 53557 41515 53623 41518
rect 54697 41488 55497 41518
rect 27337 41442 27403 41445
rect 29821 41442 29887 41445
rect 27337 41440 29887 41442
rect 27337 41384 27342 41440
rect 27398 41384 29826 41440
rect 29882 41384 29887 41440
rect 27337 41382 29887 41384
rect 27337 41379 27403 41382
rect 29821 41379 29887 41382
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 29545 41306 29611 41309
rect 32581 41306 32647 41309
rect 29545 41304 32647 41306
rect 29545 41248 29550 41304
rect 29606 41248 32586 41304
rect 32642 41248 32647 41304
rect 29545 41246 32647 41248
rect 29545 41243 29611 41246
rect 32581 41243 32647 41246
rect 8017 41170 8083 41173
rect 38653 41170 38719 41173
rect 8017 41168 38719 41170
rect 8017 41112 8022 41168
rect 8078 41112 38658 41168
rect 38714 41112 38719 41168
rect 8017 41110 38719 41112
rect 8017 41107 8083 41110
rect 38653 41107 38719 41110
rect 18781 41034 18847 41037
rect 30741 41034 30807 41037
rect 18781 41032 30807 41034
rect 18781 40976 18786 41032
rect 18842 40976 30746 41032
rect 30802 40976 30807 41032
rect 18781 40974 30807 40976
rect 18781 40971 18847 40974
rect 30741 40971 30807 40974
rect 0 40898 800 40928
rect 1485 40898 1551 40901
rect 0 40896 1551 40898
rect 0 40840 1490 40896
rect 1546 40840 1551 40896
rect 0 40838 1551 40840
rect 0 40808 800 40838
rect 1485 40835 1551 40838
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 28901 40762 28967 40765
rect 33777 40762 33843 40765
rect 28901 40760 33843 40762
rect 28901 40704 28906 40760
rect 28962 40704 33782 40760
rect 33838 40704 33843 40760
rect 28901 40702 33843 40704
rect 28901 40699 28967 40702
rect 33777 40699 33843 40702
rect 19977 40626 20043 40629
rect 49141 40626 49207 40629
rect 19977 40624 49207 40626
rect 19977 40568 19982 40624
rect 20038 40568 49146 40624
rect 49202 40568 49207 40624
rect 19977 40566 49207 40568
rect 19977 40563 20043 40566
rect 49141 40563 49207 40566
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 53557 39538 53623 39541
rect 54697 39538 55497 39568
rect 53557 39536 55497 39538
rect 53557 39480 53562 39536
rect 53618 39480 55497 39536
rect 53557 39478 55497 39480
rect 53557 39475 53623 39478
rect 54697 39448 55497 39478
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 29545 39130 29611 39133
rect 31569 39130 31635 39133
rect 29545 39128 31635 39130
rect 29545 39072 29550 39128
rect 29606 39072 31574 39128
rect 31630 39072 31635 39128
rect 29545 39070 31635 39072
rect 29545 39067 29611 39070
rect 31569 39067 31635 39070
rect 0 38858 800 38888
rect 1577 38858 1643 38861
rect 0 38856 1643 38858
rect 0 38800 1582 38856
rect 1638 38800 1643 38856
rect 0 38798 1643 38800
rect 0 38768 800 38798
rect 1577 38795 1643 38798
rect 21909 38722 21975 38725
rect 22553 38722 22619 38725
rect 21909 38720 22619 38722
rect 21909 38664 21914 38720
rect 21970 38664 22558 38720
rect 22614 38664 22619 38720
rect 21909 38662 22619 38664
rect 21909 38659 21975 38662
rect 22553 38659 22619 38662
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 30557 38450 30623 38453
rect 30741 38450 30807 38453
rect 30557 38448 30807 38450
rect 30557 38392 30562 38448
rect 30618 38392 30746 38448
rect 30802 38392 30807 38448
rect 30557 38390 30807 38392
rect 30557 38387 30623 38390
rect 30741 38387 30807 38390
rect 33409 38314 33475 38317
rect 38469 38314 38535 38317
rect 33409 38312 38535 38314
rect 33409 38256 33414 38312
rect 33470 38256 38474 38312
rect 38530 38256 38535 38312
rect 33409 38254 38535 38256
rect 33409 38251 33475 38254
rect 38469 38251 38535 38254
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 53557 36818 53623 36821
rect 54697 36818 55497 36848
rect 53557 36816 55497 36818
rect 53557 36760 53562 36816
rect 53618 36760 55497 36816
rect 53557 36758 55497 36760
rect 53557 36755 53623 36758
rect 54697 36728 55497 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 34237 36274 34303 36277
rect 35065 36274 35131 36277
rect 34237 36272 35131 36274
rect 34237 36216 34242 36272
rect 34298 36216 35070 36272
rect 35126 36216 35131 36272
rect 34237 36214 35131 36216
rect 34237 36211 34303 36214
rect 35065 36211 35131 36214
rect 0 36138 800 36168
rect 1853 36138 1919 36141
rect 0 36136 1919 36138
rect 0 36080 1858 36136
rect 1914 36080 1919 36136
rect 0 36078 1919 36080
rect 0 36048 800 36078
rect 1853 36075 1919 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 1945 35186 2011 35189
rect 35341 35186 35407 35189
rect 1945 35184 35407 35186
rect 1945 35128 1950 35184
rect 2006 35128 35346 35184
rect 35402 35128 35407 35184
rect 1945 35126 35407 35128
rect 1945 35123 2011 35126
rect 35341 35123 35407 35126
rect 30557 35050 30623 35053
rect 34605 35050 34671 35053
rect 30557 35048 34671 35050
rect 30557 34992 30562 35048
rect 30618 34992 34610 35048
rect 34666 34992 34671 35048
rect 30557 34990 34671 34992
rect 30557 34987 30623 34990
rect 34605 34987 34671 34990
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 53557 34778 53623 34781
rect 54697 34778 55497 34808
rect 53557 34776 55497 34778
rect 53557 34720 53562 34776
rect 53618 34720 55497 34776
rect 53557 34718 55497 34720
rect 53557 34715 53623 34718
rect 54697 34688 55497 34718
rect 18229 34642 18295 34645
rect 53281 34642 53347 34645
rect 18229 34640 53347 34642
rect 18229 34584 18234 34640
rect 18290 34584 53286 34640
rect 53342 34584 53347 34640
rect 18229 34582 53347 34584
rect 18229 34579 18295 34582
rect 53281 34579 53347 34582
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 0 34098 800 34128
rect 1577 34098 1643 34101
rect 0 34096 1643 34098
rect 0 34040 1582 34096
rect 1638 34040 1643 34096
rect 0 34038 1643 34040
rect 0 34008 800 34038
rect 1577 34035 1643 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 29361 33418 29427 33421
rect 30097 33418 30163 33421
rect 29361 33416 30163 33418
rect 29361 33360 29366 33416
rect 29422 33360 30102 33416
rect 30158 33360 30163 33416
rect 29361 33358 30163 33360
rect 29361 33355 29427 33358
rect 30097 33355 30163 33358
rect 28717 33282 28783 33285
rect 29821 33282 29887 33285
rect 30925 33282 30991 33285
rect 32489 33282 32555 33285
rect 28717 33280 32555 33282
rect 28717 33224 28722 33280
rect 28778 33224 29826 33280
rect 29882 33224 30930 33280
rect 30986 33224 32494 33280
rect 32550 33224 32555 33280
rect 28717 33222 32555 33224
rect 28717 33219 28783 33222
rect 29821 33219 29887 33222
rect 30925 33219 30991 33222
rect 32489 33219 32555 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 30097 32466 30163 32469
rect 30833 32466 30899 32469
rect 30097 32464 30899 32466
rect 30097 32408 30102 32464
rect 30158 32408 30838 32464
rect 30894 32408 30899 32464
rect 30097 32406 30899 32408
rect 30097 32403 30163 32406
rect 30833 32403 30899 32406
rect 4210 32128 4526 32129
rect 0 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1485 32058 1551 32061
rect 0 32056 1551 32058
rect 0 32000 1490 32056
rect 1546 32000 1551 32056
rect 0 31998 1551 32000
rect 0 31968 800 31998
rect 1485 31995 1551 31998
rect 53557 32058 53623 32061
rect 54697 32058 55497 32088
rect 53557 32056 55497 32058
rect 53557 32000 53562 32056
rect 53618 32000 55497 32056
rect 53557 31998 55497 32000
rect 53557 31995 53623 31998
rect 54697 31968 55497 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 53557 30018 53623 30021
rect 54697 30018 55497 30048
rect 53557 30016 55497 30018
rect 53557 29960 53562 30016
rect 53618 29960 55497 30016
rect 53557 29958 55497 29960
rect 53557 29955 53623 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 54697 29928 55497 29958
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 0 29338 800 29368
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 1393 29338 1459 29341
rect 0 29336 1459 29338
rect 0 29280 1398 29336
rect 1454 29280 1459 29336
rect 0 29278 1459 29280
rect 0 29248 800 29278
rect 1393 29275 1459 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 30741 28794 30807 28797
rect 33961 28794 34027 28797
rect 30741 28792 34027 28794
rect 30741 28736 30746 28792
rect 30802 28736 33966 28792
rect 34022 28736 34027 28792
rect 30741 28734 34027 28736
rect 30741 28731 30807 28734
rect 33961 28731 34027 28734
rect 34973 28522 35039 28525
rect 36445 28522 36511 28525
rect 34973 28520 36511 28522
rect 34973 28464 34978 28520
rect 35034 28464 36450 28520
rect 36506 28464 36511 28520
rect 34973 28462 36511 28464
rect 34973 28459 35039 28462
rect 36445 28459 36511 28462
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 53649 27978 53715 27981
rect 54697 27978 55497 28008
rect 53649 27976 55497 27978
rect 53649 27920 53654 27976
rect 53710 27920 55497 27976
rect 53649 27918 55497 27920
rect 53649 27915 53715 27918
rect 54697 27888 55497 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 0 27298 800 27328
rect 1485 27298 1551 27301
rect 0 27296 1551 27298
rect 0 27240 1490 27296
rect 1546 27240 1551 27296
rect 0 27238 1551 27240
rect 0 27208 800 27238
rect 1485 27235 1551 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 0 25258 800 25288
rect 1853 25258 1919 25261
rect 0 25256 1919 25258
rect 0 25200 1858 25256
rect 1914 25200 1919 25256
rect 0 25198 1919 25200
rect 0 25168 800 25198
rect 1853 25195 1919 25198
rect 53557 25258 53623 25261
rect 54697 25258 55497 25288
rect 53557 25256 55497 25258
rect 53557 25200 53562 25256
rect 53618 25200 55497 25256
rect 53557 25198 55497 25200
rect 53557 25195 53623 25198
rect 54697 25168 55497 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 53557 23218 53623 23221
rect 54697 23218 55497 23248
rect 53557 23216 55497 23218
rect 53557 23160 53562 23216
rect 53618 23160 55497 23216
rect 53557 23158 55497 23160
rect 53557 23155 53623 23158
rect 54697 23128 55497 23158
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 0 22538 800 22568
rect 1393 22538 1459 22541
rect 0 22536 1459 22538
rect 0 22480 1398 22536
rect 1454 22480 1459 22536
rect 0 22478 1459 22480
rect 0 22448 800 22478
rect 1393 22475 1459 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 53557 21178 53623 21181
rect 54697 21178 55497 21208
rect 53557 21176 55497 21178
rect 53557 21120 53562 21176
rect 53618 21120 55497 21176
rect 53557 21118 55497 21120
rect 53557 21115 53623 21118
rect 54697 21088 55497 21118
rect 1577 20906 1643 20909
rect 21398 20906 21404 20908
rect 1577 20904 21404 20906
rect 1577 20848 1582 20904
rect 1638 20848 21404 20904
rect 1577 20846 21404 20848
rect 1577 20843 1643 20846
rect 21398 20844 21404 20846
rect 21468 20844 21474 20908
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 0 20498 800 20528
rect 1393 20498 1459 20501
rect 0 20496 1459 20498
rect 0 20440 1398 20496
rect 1454 20440 1459 20496
rect 0 20438 1459 20440
rect 0 20408 800 20438
rect 1393 20435 1459 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 53557 18458 53623 18461
rect 54697 18458 55497 18488
rect 53557 18456 55497 18458
rect 53557 18400 53562 18456
rect 53618 18400 55497 18456
rect 53557 18398 55497 18400
rect 53557 18395 53623 18398
rect 54697 18368 55497 18398
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 0 17778 800 17808
rect 1577 17778 1643 17781
rect 0 17776 1643 17778
rect 0 17720 1582 17776
rect 1638 17720 1643 17776
rect 0 17718 1643 17720
rect 0 17688 800 17718
rect 1577 17715 1643 17718
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 53557 16418 53623 16421
rect 54697 16418 55497 16448
rect 53557 16416 55497 16418
rect 53557 16360 53562 16416
rect 53618 16360 55497 16416
rect 53557 16358 55497 16360
rect 53557 16355 53623 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 54697 16328 55497 16358
rect 50290 16287 50606 16288
rect 4210 15808 4526 15809
rect 0 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1393 15738 1459 15741
rect 0 15736 1459 15738
rect 0 15680 1398 15736
rect 1454 15680 1459 15736
rect 0 15678 1459 15680
rect 0 15648 800 15678
rect 1393 15675 1459 15678
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 0 13698 800 13728
rect 1485 13698 1551 13701
rect 0 13696 1551 13698
rect 0 13640 1490 13696
rect 1546 13640 1551 13696
rect 0 13638 1551 13640
rect 0 13608 800 13638
rect 1485 13635 1551 13638
rect 53649 13698 53715 13701
rect 54697 13698 55497 13728
rect 53649 13696 55497 13698
rect 53649 13640 53654 13696
rect 53710 13640 55497 13696
rect 53649 13638 55497 13640
rect 53649 13635 53715 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 54697 13608 55497 13638
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 53557 11658 53623 11661
rect 54697 11658 55497 11688
rect 53557 11656 55497 11658
rect 53557 11600 53562 11656
rect 53618 11600 55497 11656
rect 53557 11598 55497 11600
rect 53557 11595 53623 11598
rect 54697 11568 55497 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 0 10978 800 11008
rect 1577 10978 1643 10981
rect 0 10976 1643 10978
rect 0 10920 1582 10976
rect 1638 10920 1643 10976
rect 0 10918 1643 10920
rect 0 10888 800 10918
rect 1577 10915 1643 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 53557 9618 53623 9621
rect 54697 9618 55497 9648
rect 53557 9616 55497 9618
rect 53557 9560 53562 9616
rect 53618 9560 55497 9616
rect 53557 9558 55497 9560
rect 53557 9555 53623 9558
rect 54697 9528 55497 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 0 8938 800 8968
rect 1485 8938 1551 8941
rect 0 8936 1551 8938
rect 0 8880 1490 8936
rect 1546 8880 1551 8936
rect 0 8878 1551 8880
rect 0 8848 800 8878
rect 1485 8875 1551 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 0 6898 800 6928
rect 1577 6898 1643 6901
rect 0 6896 1643 6898
rect 0 6840 1582 6896
rect 1638 6840 1643 6896
rect 0 6838 1643 6840
rect 0 6808 800 6838
rect 1577 6835 1643 6838
rect 53649 6898 53715 6901
rect 54697 6898 55497 6928
rect 53649 6896 55497 6898
rect 53649 6840 53654 6896
rect 53710 6840 55497 6896
rect 53649 6838 55497 6840
rect 53649 6835 53715 6838
rect 54697 6808 55497 6838
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 53557 4858 53623 4861
rect 54697 4858 55497 4888
rect 53557 4856 55497 4858
rect 53557 4800 53562 4856
rect 53618 4800 55497 4856
rect 53557 4798 55497 4800
rect 53557 4795 53623 4798
rect 54697 4768 55497 4798
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 0 4178 800 4208
rect 1485 4178 1551 4181
rect 0 4176 1551 4178
rect 0 4120 1490 4176
rect 1546 4120 1551 4176
rect 0 4118 1551 4120
rect 0 4088 800 4118
rect 1485 4115 1551 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 53557 2818 53623 2821
rect 54697 2818 55497 2848
rect 53557 2816 55497 2818
rect 53557 2760 53562 2816
rect 53618 2760 55497 2816
rect 53557 2758 55497 2760
rect 53557 2755 53623 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 54697 2728 55497 2758
rect 34930 2687 35246 2688
rect 24577 2546 24643 2549
rect 30966 2546 30972 2548
rect 24577 2544 30972 2546
rect 24577 2488 24582 2544
rect 24638 2488 30972 2544
rect 24577 2486 30972 2488
rect 24577 2483 24643 2486
rect 30966 2484 30972 2486
rect 31036 2484 31042 2548
rect 9121 2410 9187 2413
rect 20662 2410 20668 2412
rect 9121 2408 20668 2410
rect 9121 2352 9126 2408
rect 9182 2352 20668 2408
rect 9121 2350 20668 2352
rect 9121 2347 9187 2350
rect 20662 2348 20668 2350
rect 20732 2348 20738 2412
rect 23790 2348 23796 2412
rect 23860 2410 23866 2412
rect 45369 2410 45435 2413
rect 23860 2408 45435 2410
rect 23860 2352 45374 2408
rect 45430 2352 45435 2408
rect 23860 2350 45435 2352
rect 23860 2348 23866 2350
rect 45369 2347 45435 2350
rect 19570 2208 19886 2209
rect 0 2138 800 2168
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
rect 1853 2138 1919 2141
rect 0 2136 1919 2138
rect 0 2080 1858 2136
rect 1914 2080 1919 2136
rect 0 2078 1919 2080
rect 0 2048 800 2078
rect 1853 2075 1919 2078
rect 53557 98 53623 101
rect 54697 98 55497 128
rect 53557 96 55497 98
rect 53557 40 53562 96
rect 53618 40 55497 96
rect 53557 38 55497 40
rect 53557 35 53623 38
rect 54697 8 55497 38
<< via3 >>
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 21404 49676 21468 49740
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 23796 48452 23860 48516
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 20668 47424 20732 47428
rect 20668 47368 20718 47424
rect 20718 47368 20732 47424
rect 20668 47364 20732 47368
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 30972 47016 31036 47020
rect 30972 46960 30986 47016
rect 30986 46960 31036 47016
rect 30972 46956 31036 46960
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 21404 20844 21468 20908
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 30972 2484 31036 2548
rect 20668 2348 20732 2412
rect 23796 2348 23860 2412
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 54976 4528 54992
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 54432 19888 54992
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 34928 54976 35248 54992
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 21403 49740 21469 49741
rect 21403 49676 21404 49740
rect 21468 49676 21469 49740
rect 21403 49675 21469 49676
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 20667 47428 20733 47429
rect 20667 47364 20668 47428
rect 20732 47364 20733 47428
rect 20667 47363 20733 47364
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 20670 2413 20730 47363
rect 21406 20909 21466 49675
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 23795 48516 23861 48517
rect 23795 48452 23796 48516
rect 23860 48452 23861 48516
rect 23795 48451 23861 48452
rect 21403 20908 21469 20909
rect 21403 20844 21404 20908
rect 21468 20844 21469 20908
rect 21403 20843 21469 20844
rect 23798 2413 23858 48451
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 30971 47020 31037 47021
rect 30971 46956 30972 47020
rect 31036 46956 31037 47020
rect 30971 46955 31037 46956
rect 30974 2549 31034 46955
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 30971 2548 31037 2549
rect 30971 2484 30972 2548
rect 31036 2484 31037 2548
rect 30971 2483 31037 2484
rect 20667 2412 20733 2413
rect 20667 2348 20668 2412
rect 20732 2348 20733 2412
rect 20667 2347 20733 2348
rect 23795 2412 23861 2413
rect 23795 2348 23796 2412
rect 23860 2348 23861 2412
rect 23795 2347 23861 2348
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2128 35248 2688
rect 50288 54432 50608 54992
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__A dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21344 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__B
timestamp 1649977179
transform -1 0 22080 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__A
timestamp 1649977179
transform 1 0 20056 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__B
timestamp 1649977179
transform -1 0 20792 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A
timestamp 1649977179
transform -1 0 25116 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__A
timestamp 1649977179
transform -1 0 21344 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__B
timestamp 1649977179
transform 1 0 20608 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__A1
timestamp 1649977179
transform -1 0 21344 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__A2
timestamp 1649977179
transform -1 0 24472 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__A
timestamp 1649977179
transform 1 0 20792 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__B
timestamp 1649977179
transform 1 0 22080 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__A
timestamp 1649977179
transform 1 0 21620 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__B
timestamp 1649977179
transform 1 0 21344 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A
timestamp 1649977179
transform 1 0 36064 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__A
timestamp 1649977179
transform 1 0 30636 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__B
timestamp 1649977179
transform -1 0 33120 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__A
timestamp 1649977179
transform 1 0 22264 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__A
timestamp 1649977179
transform 1 0 21160 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__B
timestamp 1649977179
transform 1 0 20148 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A
timestamp 1649977179
transform 1 0 24748 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__B
timestamp 1649977179
transform 1 0 22080 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__B
timestamp 1649977179
transform 1 0 20700 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__A
timestamp 1649977179
transform -1 0 40020 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__B
timestamp 1649977179
transform -1 0 40572 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A
timestamp 1649977179
transform 1 0 30636 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__A
timestamp 1649977179
transform -1 0 33948 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__B1
timestamp 1649977179
transform 1 0 22264 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__A
timestamp 1649977179
transform 1 0 28060 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__A
timestamp 1649977179
transform 1 0 32108 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__B
timestamp 1649977179
transform -1 0 22264 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A
timestamp 1649977179
transform -1 0 35696 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__C1
timestamp 1649977179
transform 1 0 23736 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A2
timestamp 1649977179
transform 1 0 24380 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A
timestamp 1649977179
transform 1 0 28888 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__B
timestamp 1649977179
transform 1 0 24840 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__B
timestamp 1649977179
transform 1 0 24380 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A
timestamp 1649977179
transform -1 0 26312 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__A
timestamp 1649977179
transform 1 0 34040 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__B
timestamp 1649977179
transform 1 0 27048 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__B
timestamp 1649977179
transform 1 0 26220 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__B
timestamp 1649977179
transform 1 0 28428 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A
timestamp 1649977179
transform 1 0 36248 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A1
timestamp 1649977179
transform 1 0 28060 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__B2
timestamp 1649977179
transform -1 0 28060 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__C1
timestamp 1649977179
transform -1 0 28152 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A1
timestamp 1649977179
transform 1 0 26772 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__A
timestamp 1649977179
transform -1 0 33856 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A
timestamp 1649977179
transform -1 0 33304 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__A2
timestamp 1649977179
transform -1 0 22816 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__B1
timestamp 1649977179
transform 1 0 21988 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__C1
timestamp 1649977179
transform -1 0 23000 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__A
timestamp 1649977179
transform 1 0 32108 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__A
timestamp 1649977179
transform -1 0 30636 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__A
timestamp 1649977179
transform -1 0 27140 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__A
timestamp 1649977179
transform 1 0 31924 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__B
timestamp 1649977179
transform 1 0 30268 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__A
timestamp 1649977179
transform 1 0 35052 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__B
timestamp 1649977179
transform 1 0 32844 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__A2
timestamp 1649977179
transform 1 0 28060 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__B1
timestamp 1649977179
transform 1 0 31648 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__B
timestamp 1649977179
transform 1 0 28428 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__C
timestamp 1649977179
transform 1 0 34040 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__A1
timestamp 1649977179
transform 1 0 32108 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__B2
timestamp 1649977179
transform 1 0 28796 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__C1
timestamp 1649977179
transform 1 0 27416 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__A1
timestamp 1649977179
transform -1 0 28980 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__A
timestamp 1649977179
transform -1 0 31188 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__B
timestamp 1649977179
transform -1 0 31556 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__A
timestamp 1649977179
transform 1 0 30820 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__B
timestamp 1649977179
transform 1 0 30268 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A
timestamp 1649977179
transform -1 0 32844 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A
timestamp 1649977179
transform 1 0 28888 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__B1
timestamp 1649977179
transform -1 0 29716 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A
timestamp 1649977179
transform -1 0 36524 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__B
timestamp 1649977179
transform -1 0 35972 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__A
timestamp 1649977179
transform 1 0 35236 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__B
timestamp 1649977179
transform 1 0 32660 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A
timestamp 1649977179
transform 1 0 40388 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__B
timestamp 1649977179
transform -1 0 41124 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A
timestamp 1649977179
transform -1 0 34868 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__B
timestamp 1649977179
transform 1 0 31464 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__C
timestamp 1649977179
transform -1 0 34868 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__D
timestamp 1649977179
transform 1 0 29348 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__A
timestamp 1649977179
transform 1 0 35420 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A1
timestamp 1649977179
transform 1 0 34040 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__A1
timestamp 1649977179
transform -1 0 29624 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__B1
timestamp 1649977179
transform -1 0 30268 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__A
timestamp 1649977179
transform -1 0 35420 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__B
timestamp 1649977179
transform 1 0 35696 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A
timestamp 1649977179
transform 1 0 35236 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__A
timestamp 1649977179
transform -1 0 33764 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__A
timestamp 1649977179
transform -1 0 37352 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__B
timestamp 1649977179
transform 1 0 36616 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__A
timestamp 1649977179
transform 1 0 35696 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__B
timestamp 1649977179
transform 1 0 36248 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__A
timestamp 1649977179
transform 1 0 36340 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A1
timestamp 1649977179
transform 1 0 37260 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__B2
timestamp 1649977179
transform -1 0 37628 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__C1
timestamp 1649977179
transform 1 0 36892 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__A1
timestamp 1649977179
transform 1 0 32476 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__A
timestamp 1649977179
transform 1 0 36064 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__B
timestamp 1649977179
transform 1 0 35788 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__B1
timestamp 1649977179
transform -1 0 36432 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__B2
timestamp 1649977179
transform 1 0 35696 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A
timestamp 1649977179
transform 1 0 37352 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__A
timestamp 1649977179
transform -1 0 37996 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A
timestamp 1649977179
transform 1 0 35788 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__A
timestamp 1649977179
transform 1 0 36708 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__B
timestamp 1649977179
transform 1 0 36156 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__A
timestamp 1649977179
transform 1 0 37260 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__B
timestamp 1649977179
transform 1 0 36156 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A1
timestamp 1649977179
transform 1 0 37260 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__B1
timestamp 1649977179
transform 1 0 36248 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A
timestamp 1649977179
transform 1 0 36800 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__B
timestamp 1649977179
transform 1 0 35972 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A
timestamp 1649977179
transform 1 0 36524 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__A1
timestamp 1649977179
transform 1 0 36064 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__B1
timestamp 1649977179
transform 1 0 37260 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__A1
timestamp 1649977179
transform 1 0 36248 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__A2
timestamp 1649977179
transform -1 0 35696 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__B1
timestamp 1649977179
transform 1 0 36800 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__B2
timestamp 1649977179
transform 1 0 36616 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A1
timestamp 1649977179
transform -1 0 36432 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A2
timestamp 1649977179
transform -1 0 37444 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A
timestamp 1649977179
transform 1 0 40388 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__B
timestamp 1649977179
transform -1 0 39652 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__A
timestamp 1649977179
transform 1 0 38364 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__B
timestamp 1649977179
transform -1 0 40204 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__A
timestamp 1649977179
transform -1 0 39100 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__A
timestamp 1649977179
transform -1 0 38548 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__B1
timestamp 1649977179
transform 1 0 37812 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__A
timestamp 1649977179
transform 1 0 38916 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__B
timestamp 1649977179
transform 1 0 39836 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A
timestamp 1649977179
transform 1 0 36800 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__B
timestamp 1649977179
transform 1 0 37812 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__A
timestamp 1649977179
transform 1 0 35604 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__B
timestamp 1649977179
transform 1 0 34684 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__A
timestamp 1649977179
transform 1 0 37904 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__A
timestamp 1649977179
transform -1 0 37444 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__A1
timestamp 1649977179
transform 1 0 37812 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__B2
timestamp 1649977179
transform -1 0 37444 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__C1
timestamp 1649977179
transform 1 0 37812 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__A
timestamp 1649977179
transform -1 0 39100 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__B
timestamp 1649977179
transform 1 0 40940 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A
timestamp 1649977179
transform 1 0 42596 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__B
timestamp 1649977179
transform -1 0 41768 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A
timestamp 1649977179
transform 1 0 40020 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__A
timestamp 1649977179
transform 1 0 41032 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A
timestamp 1649977179
transform 1 0 40480 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__A
timestamp 1649977179
transform 1 0 40388 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A
timestamp 1649977179
transform 1 0 40388 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__B
timestamp 1649977179
transform 1 0 39836 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__A
timestamp 1649977179
transform 1 0 39008 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__B
timestamp 1649977179
transform -1 0 38640 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__A1
timestamp 1649977179
transform 1 0 37260 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__B2
timestamp 1649977179
transform -1 0 38456 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A1
timestamp 1649977179
transform -1 0 40020 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__A
timestamp 1649977179
transform -1 0 39008 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__A
timestamp 1649977179
transform 1 0 35880 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__B
timestamp 1649977179
transform 1 0 33948 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A
timestamp 1649977179
transform 1 0 39008 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__B
timestamp 1649977179
transform 1 0 38364 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__A
timestamp 1649977179
transform -1 0 39560 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__B
timestamp 1649977179
transform 1 0 38364 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A1
timestamp 1649977179
transform 1 0 37352 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A2
timestamp 1649977179
transform 1 0 38824 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__A
timestamp 1649977179
transform 1 0 39836 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__B
timestamp 1649977179
transform 1 0 39008 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A1
timestamp 1649977179
transform 1 0 40480 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__B1
timestamp 1649977179
transform 1 0 40388 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__B1
timestamp 1649977179
transform 1 0 32568 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A1
timestamp 1649977179
transform -1 0 41216 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A2
timestamp 1649977179
transform -1 0 40664 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__B1
timestamp 1649977179
transform 1 0 40940 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__B2
timestamp 1649977179
transform 1 0 39928 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__A
timestamp 1649977179
transform 1 0 39836 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A
timestamp 1649977179
transform 1 0 42044 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__B
timestamp 1649977179
transform 1 0 41492 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__B1
timestamp 1649977179
transform 1 0 38916 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__A
timestamp 1649977179
transform -1 0 40756 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__A
timestamp 1649977179
transform -1 0 39652 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__A1
timestamp 1649977179
transform -1 0 38088 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__D1
timestamp 1649977179
transform 1 0 38456 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__A
timestamp 1649977179
transform -1 0 35512 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__A
timestamp 1649977179
transform 1 0 41584 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__B
timestamp 1649977179
transform 1 0 41032 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__A1
timestamp 1649977179
transform 1 0 40940 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__A
timestamp 1649977179
transform 1 0 39100 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A
timestamp 1649977179
transform 1 0 38548 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__B1
timestamp 1649977179
transform 1 0 35788 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__B1
timestamp 1649977179
transform -1 0 40020 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__A1
timestamp 1649977179
transform 1 0 34592 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__B2
timestamp 1649977179
transform 1 0 32292 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__A
timestamp 1649977179
transform -1 0 38824 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__B
timestamp 1649977179
transform -1 0 40020 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A
timestamp 1649977179
transform 1 0 38364 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__B
timestamp 1649977179
transform 1 0 37628 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__A1
timestamp 1649977179
transform 1 0 41492 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__A2
timestamp 1649977179
transform 1 0 40940 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__B1
timestamp 1649977179
transform -1 0 41768 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__A1
timestamp 1649977179
transform 1 0 42412 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__A2
timestamp 1649977179
transform -1 0 41676 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__A
timestamp 1649977179
transform 1 0 40388 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A
timestamp 1649977179
transform 1 0 39836 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A
timestamp 1649977179
transform -1 0 39008 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__B
timestamp 1649977179
transform 1 0 38272 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A
timestamp 1649977179
transform 1 0 37076 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__B
timestamp 1649977179
transform 1 0 36432 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A
timestamp 1649977179
transform 1 0 40480 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__B
timestamp 1649977179
transform 1 0 39928 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A1
timestamp 1649977179
transform 1 0 39376 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__B1
timestamp 1649977179
transform 1 0 36524 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__B
timestamp 1649977179
transform 1 0 36064 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A1
timestamp 1649977179
transform 1 0 33212 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A
timestamp 1649977179
transform 1 0 31464 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__A1
timestamp 1649977179
transform 1 0 32844 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__C1
timestamp 1649977179
transform 1 0 33396 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A
timestamp 1649977179
transform -1 0 37444 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__B
timestamp 1649977179
transform -1 0 37904 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__A
timestamp 1649977179
transform 1 0 38180 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__B
timestamp 1649977179
transform 1 0 37168 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A
timestamp 1649977179
transform 1 0 33488 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A
timestamp 1649977179
transform -1 0 30268 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__B1
timestamp 1649977179
transform 1 0 34132 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A
timestamp 1649977179
transform 1 0 34040 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A1
timestamp 1649977179
transform 1 0 32936 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__A
timestamp 1649977179
transform 1 0 38732 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__B
timestamp 1649977179
transform 1 0 38180 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__A
timestamp 1649977179
transform 1 0 37812 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__B
timestamp 1649977179
transform 1 0 38088 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A1
timestamp 1649977179
transform 1 0 30728 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__B2
timestamp 1649977179
transform 1 0 31004 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__A
timestamp 1649977179
transform 1 0 29992 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__A
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__B
timestamp 1649977179
transform 1 0 36432 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A
timestamp 1649977179
transform 1 0 35236 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A
timestamp 1649977179
transform 1 0 28980 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__B
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__A
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__B
timestamp 1649977179
transform -1 0 28152 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__A
timestamp 1649977179
transform 1 0 37996 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__B
timestamp 1649977179
transform 1 0 36616 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A1
timestamp 1649977179
transform 1 0 38916 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A2
timestamp 1649977179
transform 1 0 37260 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A
timestamp 1649977179
transform -1 0 31740 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__B
timestamp 1649977179
transform 1 0 34684 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__A
timestamp 1649977179
transform 1 0 29624 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__A1
timestamp 1649977179
transform 1 0 33580 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__B2
timestamp 1649977179
transform 1 0 28428 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__C1
timestamp 1649977179
transform 1 0 33488 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A1
timestamp 1649977179
transform 1 0 32752 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A
timestamp 1649977179
transform -1 0 28152 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__B
timestamp 1649977179
transform 1 0 28704 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A
timestamp 1649977179
transform 1 0 31188 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__A
timestamp 1649977179
transform 1 0 32108 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__A
timestamp 1649977179
transform -1 0 37996 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__B
timestamp 1649977179
transform 1 0 36156 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__A
timestamp 1649977179
transform 1 0 37168 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__B
timestamp 1649977179
transform -1 0 37904 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__A
timestamp 1649977179
transform 1 0 37536 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__B
timestamp 1649977179
transform -1 0 37168 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__A
timestamp 1649977179
transform 1 0 31372 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__A1
timestamp 1649977179
transform 1 0 34040 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__C1
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A1
timestamp 1649977179
transform 1 0 38364 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A1
timestamp 1649977179
transform 1 0 32660 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__B2
timestamp 1649977179
transform 1 0 31740 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__A
timestamp 1649977179
transform 1 0 28888 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__A
timestamp 1649977179
transform 1 0 36616 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__B
timestamp 1649977179
transform 1 0 35880 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__A
timestamp 1649977179
transform 1 0 14168 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__B
timestamp 1649977179
transform 1 0 15272 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A
timestamp 1649977179
transform -1 0 17664 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__B
timestamp 1649977179
transform 1 0 15824 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__A1
timestamp 1649977179
transform -1 0 15548 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__A2
timestamp 1649977179
transform -1 0 16100 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__A
timestamp 1649977179
transform 1 0 15456 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__B
timestamp 1649977179
transform 1 0 16008 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__A
timestamp 1649977179
transform 1 0 31372 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__A
timestamp 1649977179
transform -1 0 34868 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__A
timestamp 1649977179
transform 1 0 31464 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__A
timestamp 1649977179
transform 1 0 30544 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A
timestamp 1649977179
transform -1 0 24564 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__B
timestamp 1649977179
transform 1 0 21804 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__A
timestamp 1649977179
transform -1 0 19780 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__B
timestamp 1649977179
transform 1 0 22356 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A1
timestamp 1649977179
transform 1 0 28060 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A2
timestamp 1649977179
transform -1 0 29072 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__B1
timestamp 1649977179
transform -1 0 31004 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__C1
timestamp 1649977179
transform 1 0 33396 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__A1
timestamp 1649977179
transform -1 0 31556 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__A2
timestamp 1649977179
transform -1 0 26220 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__A1
timestamp 1649977179
transform 1 0 34040 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__B2
timestamp 1649977179
transform 1 0 35512 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__C1
timestamp 1649977179
transform 1 0 34868 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__A
timestamp 1649977179
transform -1 0 21988 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__B
timestamp 1649977179
transform 1 0 21528 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__A
timestamp 1649977179
transform 1 0 20608 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__B
timestamp 1649977179
transform 1 0 19228 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__B1
timestamp 1649977179
transform 1 0 23736 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__A
timestamp 1649977179
transform 1 0 17112 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__B
timestamp 1649977179
transform 1 0 17664 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__A
timestamp 1649977179
transform -1 0 15180 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__B
timestamp 1649977179
transform -1 0 16560 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__A
timestamp 1649977179
transform -1 0 18400 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__B1
timestamp 1649977179
transform -1 0 18952 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__A1
timestamp 1649977179
transform 1 0 28888 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__A
timestamp 1649977179
transform -1 0 19780 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__A
timestamp 1649977179
transform 1 0 31280 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__B
timestamp 1649977179
transform 1 0 31372 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__C
timestamp 1649977179
transform 1 0 30820 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__A1
timestamp 1649977179
transform 1 0 30176 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__A2
timestamp 1649977179
transform 1 0 30268 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__B1
timestamp 1649977179
transform 1 0 29624 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__B
timestamp 1649977179
transform 1 0 29072 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__B1
timestamp 1649977179
transform 1 0 25760 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__A1
timestamp 1649977179
transform 1 0 28428 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__B1
timestamp 1649977179
transform 1 0 26312 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__A1
timestamp 1649977179
transform 1 0 31556 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__A
timestamp 1649977179
transform 1 0 21252 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__B
timestamp 1649977179
transform -1 0 18768 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__A
timestamp 1649977179
transform 1 0 18768 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__B
timestamp 1649977179
transform -1 0 23000 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__A1
timestamp 1649977179
transform 1 0 18584 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__A2
timestamp 1649977179
transform 1 0 19320 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__A
timestamp 1649977179
transform -1 0 14352 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__B
timestamp 1649977179
transform 1 0 14352 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__A
timestamp 1649977179
transform 1 0 13432 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__B
timestamp 1649977179
transform 1 0 13616 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__A1
timestamp 1649977179
transform 1 0 14444 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__A2
timestamp 1649977179
transform 1 0 13432 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__A
timestamp 1649977179
transform 1 0 19320 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__A
timestamp 1649977179
transform 1 0 19596 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__A1
timestamp 1649977179
transform 1 0 22356 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__B2
timestamp 1649977179
transform 1 0 22632 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__B1
timestamp 1649977179
transform 1 0 28244 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__A
timestamp 1649977179
transform 1 0 21160 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__B
timestamp 1649977179
transform 1 0 20976 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__A
timestamp 1649977179
transform -1 0 22540 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__B
timestamp 1649977179
transform 1 0 22816 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__A
timestamp 1649977179
transform 1 0 24656 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__A
timestamp 1649977179
transform 1 0 26312 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__B
timestamp 1649977179
transform 1 0 25208 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__A1
timestamp 1649977179
transform 1 0 31096 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__B1
timestamp 1649977179
transform 1 0 26128 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__A
timestamp 1649977179
transform 1 0 12972 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__B
timestamp 1649977179
transform 1 0 13708 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__A
timestamp 1649977179
transform 1 0 13524 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__B
timestamp 1649977179
transform 1 0 12880 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__B1
timestamp 1649977179
transform -1 0 16192 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__A
timestamp 1649977179
transform 1 0 19872 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__A1
timestamp 1649977179
transform -1 0 18768 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__A1
timestamp 1649977179
transform 1 0 28520 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__B2
timestamp 1649977179
transform 1 0 26404 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1158__B1
timestamp 1649977179
transform 1 0 25208 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__A1
timestamp 1649977179
transform -1 0 16652 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__A2
timestamp 1649977179
transform 1 0 16008 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__A
timestamp 1649977179
transform 1 0 15180 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__B
timestamp 1649977179
transform 1 0 15456 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__A
timestamp 1649977179
transform 1 0 15364 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__B
timestamp 1649977179
transform -1 0 14996 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__A
timestamp 1649977179
transform 1 0 18860 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__A
timestamp 1649977179
transform 1 0 23828 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__A
timestamp 1649977179
transform 1 0 27968 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__B
timestamp 1649977179
transform 1 0 27140 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__C
timestamp 1649977179
transform -1 0 28336 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__A
timestamp 1649977179
transform 1 0 18584 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__B
timestamp 1649977179
transform 1 0 21988 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__A
timestamp 1649977179
transform -1 0 21344 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__B
timestamp 1649977179
transform 1 0 23368 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__A
timestamp 1649977179
transform 1 0 21804 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__B
timestamp 1649977179
transform 1 0 23184 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__A1
timestamp 1649977179
transform -1 0 25944 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__B2
timestamp 1649977179
transform 1 0 26680 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__C1
timestamp 1649977179
transform 1 0 26312 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__A1
timestamp 1649977179
transform 1 0 26312 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__B1
timestamp 1649977179
transform 1 0 25668 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__A1
timestamp 1649977179
transform 1 0 26312 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__A
timestamp 1649977179
transform 1 0 22816 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__B
timestamp 1649977179
transform 1 0 22540 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__A
timestamp 1649977179
transform 1 0 19964 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__B
timestamp 1649977179
transform 1 0 20608 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__A
timestamp 1649977179
transform -1 0 16192 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__B
timestamp 1649977179
transform -1 0 16744 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__A
timestamp 1649977179
transform 1 0 18308 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__B
timestamp 1649977179
transform 1 0 16928 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__A
timestamp 1649977179
transform 1 0 19412 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__B1
timestamp 1649977179
transform -1 0 18768 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__A1
timestamp 1649977179
transform 1 0 17020 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__A
timestamp 1649977179
transform 1 0 17112 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__A1
timestamp 1649977179
transform 1 0 22264 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__B2
timestamp 1649977179
transform 1 0 23092 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__B1
timestamp 1649977179
transform 1 0 25760 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__A
timestamp 1649977179
transform 1 0 21252 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__B
timestamp 1649977179
transform -1 0 21988 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__A
timestamp 1649977179
transform -1 0 19228 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__B
timestamp 1649977179
transform 1 0 19596 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__A
timestamp 1649977179
transform -1 0 24564 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__B
timestamp 1649977179
transform 1 0 21160 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__A1
timestamp 1649977179
transform 1 0 25208 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__B1
timestamp 1649977179
transform 1 0 25760 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__A
timestamp 1649977179
transform 1 0 27876 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__B
timestamp 1649977179
transform 1 0 27968 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__A
timestamp 1649977179
transform -1 0 15916 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__B
timestamp 1649977179
transform -1 0 17020 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__A
timestamp 1649977179
transform 1 0 16560 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__B
timestamp 1649977179
transform 1 0 19228 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__A
timestamp 1649977179
transform 1 0 16008 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__B1
timestamp 1649977179
transform 1 0 16008 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__B1
timestamp 1649977179
transform 1 0 21712 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__A1
timestamp 1649977179
transform -1 0 25852 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1236__A1
timestamp 1649977179
transform 1 0 23736 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__A
timestamp 1649977179
transform -1 0 24840 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__A
timestamp 1649977179
transform 1 0 20148 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__B
timestamp 1649977179
transform 1 0 22816 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__A
timestamp 1649977179
transform -1 0 22448 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__B
timestamp 1649977179
transform 1 0 23368 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__B1
timestamp 1649977179
transform 1 0 22908 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__A
timestamp 1649977179
transform 1 0 26312 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__A1
timestamp 1649977179
transform -1 0 26496 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__B1
timestamp 1649977179
transform 1 0 27416 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__A
timestamp 1649977179
transform -1 0 16192 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__B
timestamp 1649977179
transform 1 0 16836 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__A
timestamp 1649977179
transform 1 0 16468 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__B
timestamp 1649977179
transform -1 0 15916 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__A
timestamp 1649977179
transform 1 0 17020 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__B1
timestamp 1649977179
transform 1 0 16008 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__B2
timestamp 1649977179
transform 1 0 27508 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__B1
timestamp 1649977179
transform -1 0 22632 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__A
timestamp 1649977179
transform 1 0 15456 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__B
timestamp 1649977179
transform -1 0 16468 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__A
timestamp 1649977179
transform -1 0 17020 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__B
timestamp 1649977179
transform -1 0 17572 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__A
timestamp 1649977179
transform -1 0 16836 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__A
timestamp 1649977179
transform -1 0 21896 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__B
timestamp 1649977179
transform 1 0 22816 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__A
timestamp 1649977179
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__B
timestamp 1649977179
transform 1 0 20884 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__A1
timestamp 1649977179
transform 1 0 23460 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__A2
timestamp 1649977179
transform 1 0 23736 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__A
timestamp 1649977179
transform 1 0 24564 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__A1
timestamp 1649977179
transform 1 0 25116 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__B2
timestamp 1649977179
transform 1 0 24012 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__C1
timestamp 1649977179
transform 1 0 25484 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__A1
timestamp 1649977179
transform 1 0 21896 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__A1
timestamp 1649977179
transform 1 0 26312 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__B1
timestamp 1649977179
transform 1 0 25208 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__A
timestamp 1649977179
transform -1 0 24840 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__B
timestamp 1649977179
transform 1 0 24472 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__A1
timestamp 1649977179
transform 1 0 16284 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__B2
timestamp 1649977179
transform 1 0 16836 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__A1
timestamp 1649977179
transform 1 0 17388 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1298__A
timestamp 1649977179
transform -1 0 17664 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1298__B
timestamp 1649977179
transform -1 0 19596 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__A
timestamp 1649977179
transform -1 0 17112 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__B
timestamp 1649977179
transform 1 0 17848 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__A
timestamp 1649977179
transform -1 0 17020 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__B1
timestamp 1649977179
transform 1 0 18860 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__A
timestamp 1649977179
transform 1 0 21436 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__B
timestamp 1649977179
transform 1 0 24012 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1310__A
timestamp 1649977179
transform 1 0 21160 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1310__B
timestamp 1649977179
transform 1 0 20792 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__A
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__A1
timestamp 1649977179
transform 1 0 25760 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__C1
timestamp 1649977179
transform 1 0 26312 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__A
timestamp 1649977179
transform 1 0 21344 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__B
timestamp 1649977179
transform 1 0 19320 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__A
timestamp 1649977179
transform 1 0 20608 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__B
timestamp 1649977179
transform -1 0 21988 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1321__A
timestamp 1649977179
transform 1 0 26864 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__A
timestamp 1649977179
transform 1 0 16008 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__B
timestamp 1649977179
transform 1 0 16836 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__A
timestamp 1649977179
transform 1 0 15456 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__B
timestamp 1649977179
transform -1 0 16192 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1328__A
timestamp 1649977179
transform -1 0 20148 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1331__A
timestamp 1649977179
transform 1 0 26036 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__A1
timestamp 1649977179
transform 1 0 26588 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__B1
timestamp 1649977179
transform 1 0 27140 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__A1
timestamp 1649977179
transform 1 0 26312 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1334__B1
timestamp 1649977179
transform 1 0 26128 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1335__A
timestamp 1649977179
transform 1 0 23736 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1335__B
timestamp 1649977179
transform 1 0 20240 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__A
timestamp 1649977179
transform -1 0 23920 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__B
timestamp 1649977179
transform 1 0 19688 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1341__A
timestamp 1649977179
transform 1 0 22632 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1343__A
timestamp 1649977179
transform 1 0 18584 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1343__B
timestamp 1649977179
transform -1 0 18216 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__A
timestamp 1649977179
transform 1 0 19780 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__B
timestamp 1649977179
transform -1 0 20516 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1348__A
timestamp 1649977179
transform 1 0 19136 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__B1
timestamp 1649977179
transform -1 0 18768 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1353__A1
timestamp 1649977179
transform -1 0 18768 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__A1
timestamp 1649977179
transform 1 0 19136 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1356__B1
timestamp 1649977179
transform -1 0 18768 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1358__A1
timestamp 1649977179
transform 1 0 20608 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1358__B1
timestamp 1649977179
transform 1 0 28244 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__A1
timestamp 1649977179
transform 1 0 23828 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1360__B1
timestamp 1649977179
transform 1 0 27692 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1361__A
timestamp 1649977179
transform 1 0 21620 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1361__B
timestamp 1649977179
transform 1 0 19412 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1362__A
timestamp 1649977179
transform -1 0 20148 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1362__B
timestamp 1649977179
transform 1 0 19320 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1364__A
timestamp 1649977179
transform -1 0 17664 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1364__B
timestamp 1649977179
transform -1 0 18216 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1367__A
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1370__B1
timestamp 1649977179
transform 1 0 23460 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1376__A
timestamp 1649977179
transform 1 0 24564 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1376__B
timestamp 1649977179
transform 1 0 25116 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1377__A
timestamp 1649977179
transform 1 0 22908 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1377__B
timestamp 1649977179
transform 1 0 24472 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1381__A
timestamp 1649977179
transform -1 0 25576 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1381__B
timestamp 1649977179
transform 1 0 23736 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__A1
timestamp 1649977179
transform 1 0 24380 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__A2
timestamp 1649977179
transform 1 0 27140 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__B1
timestamp 1649977179
transform 1 0 26312 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1383__C
timestamp 1649977179
transform -1 0 25944 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1384__A1
timestamp 1649977179
transform -1 0 23828 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1386__A
timestamp 1649977179
transform 1 0 27600 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1387__A
timestamp 1649977179
transform 1 0 27508 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1387__B
timestamp 1649977179
transform 1 0 26772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1388__A
timestamp 1649977179
transform 1 0 28060 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1388__B
timestamp 1649977179
transform 1 0 27324 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__B1
timestamp 1649977179
transform -1 0 27140 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__A
timestamp 1649977179
transform 1 0 20884 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__B
timestamp 1649977179
transform 1 0 20056 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__A
timestamp 1649977179
transform 1 0 22540 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__B
timestamp 1649977179
transform -1 0 19596 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1398__A
timestamp 1649977179
transform 1 0 22356 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1399__A1
timestamp 1649977179
transform 1 0 20608 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1400__A1
timestamp 1649977179
transform 1 0 21068 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1406__A
timestamp 1649977179
transform 1 0 27600 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1407__A1
timestamp 1649977179
transform 1 0 25116 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1407__B1
timestamp 1649977179
transform 1 0 23092 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1408__A1
timestamp 1649977179
transform -1 0 26128 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__B1
timestamp 1649977179
transform -1 0 28152 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1410__A
timestamp 1649977179
transform 1 0 22908 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__A
timestamp 1649977179
transform 1 0 32660 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__B
timestamp 1649977179
transform 1 0 33488 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1413__A
timestamp 1649977179
transform -1 0 32292 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1413__B
timestamp 1649977179
transform -1 0 33396 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1415__A
timestamp 1649977179
transform 1 0 21988 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1415__B
timestamp 1649977179
transform -1 0 21988 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1418__A
timestamp 1649977179
transform 1 0 31924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1419__A
timestamp 1649977179
transform 1 0 29072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1421__B1
timestamp 1649977179
transform -1 0 27968 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1423__A
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1424__A
timestamp 1649977179
transform -1 0 29716 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1425__A
timestamp 1649977179
transform 1 0 32476 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1425__B
timestamp 1649977179
transform 1 0 29992 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1426__A
timestamp 1649977179
transform 1 0 32384 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1426__B
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1430__B1
timestamp 1649977179
transform 1 0 28244 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1431__A1
timestamp 1649977179
transform 1 0 28612 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__B1
timestamp 1649977179
transform 1 0 29348 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1433__A
timestamp 1649977179
transform -1 0 34500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1433__B
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__A
timestamp 1649977179
transform 1 0 31464 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1437__C1
timestamp 1649977179
transform 1 0 33764 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1440__A
timestamp 1649977179
transform -1 0 31188 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1444__A
timestamp 1649977179
transform -1 0 32016 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1445__C1
timestamp 1649977179
transform 1 0 34040 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1449__A
timestamp 1649977179
transform 1 0 22908 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__A2
timestamp 1649977179
transform -1 0 27140 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__C1
timestamp 1649977179
transform 1 0 23920 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__A1
timestamp 1649977179
transform -1 0 28244 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1452__A1
timestamp 1649977179
transform 1 0 22356 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1452__A2
timestamp 1649977179
transform -1 0 21988 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1452__B1
timestamp 1649977179
transform 1 0 21712 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1453__A2
timestamp 1649977179
transform -1 0 22356 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1453__C1
timestamp 1649977179
transform 1 0 22724 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1649977179
transform -1 0 35420 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 52992 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 52992 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 52992 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 1748 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 50508 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 1564 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 52992 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 40940 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 1748 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 1748 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 14536 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 2668 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 6532 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 1564 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 1748 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 52992 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 24840 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 47932 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 1748 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 1748 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 1748 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 32292 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 22172 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 52256 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 2300 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 52992 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 35052 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 18768 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 52992 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 23920 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 1564 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 52992 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 22172 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 52992 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 52992 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 23276 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 45172 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 52992 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 7452 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 1748 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 27416 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 1748 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 35052 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 11684 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 27416 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 1748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 1564 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 8464 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 2852 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 48668 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 38364 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 25484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 52992 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 52992 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 1748 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 52992 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 11684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 19412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 1564 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform -1 0 52992 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1649977179
transform -1 0 29992 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1649977179
transform -1 0 45172 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1649977179
transform -1 0 43424 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1649977179
transform -1 0 3956 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1649977179
transform -1 0 11960 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1649977179
transform -1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1649977179
transform -1 0 1564 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1649977179
transform -1 0 1564 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1649977179
transform -1 0 53728 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output70_A
timestamp 1649977179
transform -1 0 15180 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output71_A
timestamp 1649977179
transform 1 0 36616 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output72_A
timestamp 1649977179
transform 1 0 13340 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output73_A
timestamp 1649977179
transform -1 0 52992 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output74_A
timestamp 1649977179
transform 1 0 52808 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output75_A
timestamp 1649977179
transform -1 0 52992 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output76_A
timestamp 1649977179
transform -1 0 40296 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output77_A
timestamp 1649977179
transform -1 0 17756 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output78_A
timestamp 1649977179
transform -1 0 52992 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output79_A
timestamp 1649977179
transform 1 0 52808 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output80_A
timestamp 1649977179
transform -1 0 51244 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output82_A
timestamp 1649977179
transform 1 0 2116 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output83_A
timestamp 1649977179
transform -1 0 52992 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output84_A
timestamp 1649977179
transform -1 0 2300 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output85_A
timestamp 1649977179
transform 1 0 2116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output86_A
timestamp 1649977179
transform 1 0 35972 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output87_A
timestamp 1649977179
transform 1 0 2116 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output88_A
timestamp 1649977179
transform 1 0 42688 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output89_A
timestamp 1649977179
transform -1 0 47104 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output90_A
timestamp 1649977179
transform -1 0 2300 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output91_A
timestamp 1649977179
transform 1 0 4692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output92_A
timestamp 1649977179
transform 1 0 17572 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output93_A
timestamp 1649977179
transform 1 0 51428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output94_A
timestamp 1649977179
transform 1 0 52808 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output95_A
timestamp 1649977179
transform 1 0 52808 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output96_A
timestamp 1649977179
transform 1 0 2116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output97_A
timestamp 1649977179
transform 1 0 2116 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output98_A
timestamp 1649977179
transform -1 0 52992 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output99_A
timestamp 1649977179
transform 1 0 6716 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output100_A
timestamp 1649977179
transform -1 0 52992 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output101_A
timestamp 1649977179
transform 1 0 52808 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1649977179
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35
timestamp 1649977179
transform 1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63
timestamp 1649977179
transform 1 0 6900 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_75
timestamp 1649977179
transform 1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1649977179
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_89 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9292 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1649977179
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115
timestamp 1649977179
transform 1 0 11684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_127
timestamp 1649977179
transform 1 0 12788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_133
timestamp 1649977179
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1649977179
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1649977179
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154
timestamp 1649977179
transform 1 0 15272 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1649977179
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1649977179
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_233
timestamp 1649977179
transform 1 0 22540 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_245
timestamp 1649977179
transform 1 0 23644 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1649977179
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_257
timestamp 1649977179
transform 1 0 24748 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_265
timestamp 1649977179
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1649977179
transform 1 0 26220 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1649977179
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_281
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1649977179
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_294
timestamp 1649977179
transform 1 0 28152 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1649977179
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_314
timestamp 1649977179
transform 1 0 29992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_328
timestamp 1649977179
transform 1 0 31280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_343
timestamp 1649977179
transform 1 0 32660 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_355
timestamp 1649977179
transform 1 0 33764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1649977179
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_365
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_373
timestamp 1649977179
transform 1 0 35420 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_385
timestamp 1649977179
transform 1 0 36524 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_388
timestamp 1649977179
transform 1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_397
timestamp 1649977179
transform 1 0 37628 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_405
timestamp 1649977179
transform 1 0 38364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_413
timestamp 1649977179
transform 1 0 39100 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1649977179
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_421
timestamp 1649977179
transform 1 0 39836 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_429
timestamp 1649977179
transform 1 0 40572 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_433
timestamp 1649977179
transform 1 0 40940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_443
timestamp 1649977179
transform 1 0 41860 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1649977179
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_449
timestamp 1649977179
transform 1 0 42412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_454
timestamp 1649977179
transform 1 0 42872 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_462
timestamp 1649977179
transform 1 0 43608 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_474
timestamp 1649977179
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_477
timestamp 1649977179
transform 1 0 44988 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_483
timestamp 1649977179
transform 1 0 45540 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_495
timestamp 1649977179
transform 1 0 46644 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_503
timestamp 1649977179
transform 1 0 47380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_505
timestamp 1649977179
transform 1 0 47564 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_515
timestamp 1649977179
transform 1 0 48484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_527
timestamp 1649977179
transform 1 0 49588 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_531
timestamp 1649977179
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_533
timestamp 1649977179
transform 1 0 50140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_543
timestamp 1649977179
transform 1 0 51060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_553
timestamp 1649977179
transform 1 0 51980 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_559
timestamp 1649977179
transform 1 0 52532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_561
timestamp 1649977179
transform 1 0 52716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_565
timestamp 1649977179
transform 1 0 53084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_572
timestamp 1649977179
transform 1 0 53728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1649977179
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_19
timestamp 1649977179
transform 1 0 2852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_31
timestamp 1649977179
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_43
timestamp 1649977179
transform 1 0 5060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_59
timestamp 1649977179
transform 1 0 6532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_71
timestamp 1649977179
transform 1 0 7636 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_83
timestamp 1649977179
transform 1 0 8740 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_95
timestamp 1649977179
transform 1 0 9844 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1649977179
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_135
timestamp 1649977179
transform 1 0 13524 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_147
timestamp 1649977179
transform 1 0 14628 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp 1649977179
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_193
timestamp 1649977179
transform 1 0 18860 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_199
timestamp 1649977179
transform 1 0 19412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_211
timestamp 1649977179
transform 1 0 20516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1649977179
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_229
timestamp 1649977179
transform 1 0 22172 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_241
timestamp 1649977179
transform 1 0 23276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_253
timestamp 1649977179
transform 1 0 24380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_265
timestamp 1649977179
transform 1 0 25484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_277
timestamp 1649977179
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1649977179
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1649977179
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1649977179
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1649977179
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1649977179
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_339
timestamp 1649977179
transform 1 0 32292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_351
timestamp 1649977179
transform 1 0 33396 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_363
timestamp 1649977179
transform 1 0 34500 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_369
timestamp 1649977179
transform 1 0 35052 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_381
timestamp 1649977179
transform 1 0 36156 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_389
timestamp 1649977179
transform 1 0 36892 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1649977179
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1649977179
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1649977179
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1649977179
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1649977179
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1649977179
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1649977179
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1649977179
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_473
timestamp 1649977179
transform 1 0 44620 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_479
timestamp 1649977179
transform 1 0 45172 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_491
timestamp 1649977179
transform 1 0 46276 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1649977179
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_505
timestamp 1649977179
transform 1 0 47564 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_509
timestamp 1649977179
transform 1 0 47932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_521
timestamp 1649977179
transform 1 0 49036 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_533
timestamp 1649977179
transform 1 0 50140 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_537
timestamp 1649977179
transform 1 0 50508 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_545
timestamp 1649977179
transform 1 0 51244 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_549
timestamp 1649977179
transform 1 0 51612 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_553
timestamp 1649977179
transform 1 0 51980 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_556
timestamp 1649977179
transform 1 0 52256 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_561
timestamp 1649977179
transform 1 0 52716 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_564
timestamp 1649977179
transform 1 0 52992 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_572
timestamp 1649977179
transform 1 0 53728 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_7
timestamp 1649977179
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_13
timestamp 1649977179
transform 1 0 2300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_25
timestamp 1649977179
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1649977179
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1649977179
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1649977179
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1649977179
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1649977179
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1649977179
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1649977179
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1649977179
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1649977179
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1649977179
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1649977179
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1649977179
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1649977179
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1649977179
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1649977179
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1649977179
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1649977179
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1649977179
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1649977179
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1649977179
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1649977179
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1649977179
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1649977179
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1649977179
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1649977179
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1649977179
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1649977179
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1649977179
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1649977179
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1649977179
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1649977179
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1649977179
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_557
timestamp 1649977179
transform 1 0 52348 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_561
timestamp 1649977179
transform 1 0 52716 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_564
timestamp 1649977179
transform 1 0 52992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_572
timestamp 1649977179
transform 1 0 53728 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1649977179
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1649977179
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1649977179
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1649977179
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1649977179
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1649977179
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1649977179
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1649977179
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1649977179
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1649977179
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1649977179
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1649977179
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1649977179
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1649977179
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1649977179
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1649977179
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1649977179
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1649977179
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1649977179
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1649977179
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1649977179
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1649977179
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1649977179
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1649977179
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1649977179
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1649977179
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1649977179
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1649977179
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1649977179
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1649977179
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_573
timestamp 1649977179
transform 1 0 53820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_7
timestamp 1649977179
transform 1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_13
timestamp 1649977179
transform 1 0 2300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1649977179
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1649977179
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1649977179
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1649977179
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1649977179
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1649977179
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1649977179
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1649977179
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1649977179
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1649977179
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1649977179
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1649977179
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1649977179
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1649977179
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1649977179
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1649977179
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1649977179
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1649977179
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1649977179
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1649977179
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1649977179
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1649977179
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1649977179
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1649977179
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1649977179
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1649977179
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1649977179
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1649977179
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1649977179
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1649977179
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1649977179
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1649977179
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1649977179
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_569
timestamp 1649977179
transform 1 0 53452 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_575
timestamp 1649977179
transform 1 0 54004 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1649977179
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1649977179
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1649977179
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1649977179
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1649977179
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1649977179
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1649977179
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1649977179
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1649977179
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1649977179
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1649977179
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1649977179
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1649977179
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1649977179
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1649977179
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1649977179
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1649977179
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1649977179
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1649977179
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1649977179
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1649977179
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1649977179
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1649977179
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1649977179
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1649977179
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1649977179
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1649977179
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1649977179
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1649977179
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1649977179
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_561
timestamp 1649977179
transform 1 0 52716 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_564
timestamp 1649977179
transform 1 0 52992 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_572
timestamp 1649977179
transform 1 0 53728 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1649977179
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1649977179
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1649977179
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1649977179
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1649977179
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1649977179
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1649977179
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1649977179
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1649977179
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1649977179
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1649977179
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1649977179
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1649977179
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1649977179
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1649977179
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1649977179
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1649977179
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1649977179
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1649977179
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1649977179
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1649977179
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1649977179
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1649977179
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1649977179
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1649977179
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1649977179
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1649977179
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1649977179
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1649977179
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_569
timestamp 1649977179
transform 1 0 53452 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_575
timestamp 1649977179
transform 1 0 54004 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1649977179
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1649977179
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1649977179
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1649977179
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1649977179
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1649977179
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1649977179
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1649977179
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1649977179
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1649977179
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1649977179
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1649977179
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1649977179
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1649977179
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1649977179
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1649977179
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1649977179
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1649977179
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1649977179
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1649977179
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1649977179
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1649977179
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1649977179
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1649977179
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1649977179
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1649977179
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_573
timestamp 1649977179
transform 1 0 53820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7
timestamp 1649977179
transform 1 0 1748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_19
timestamp 1649977179
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1649977179
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1649977179
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1649977179
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1649977179
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1649977179
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1649977179
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1649977179
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1649977179
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1649977179
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1649977179
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1649977179
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1649977179
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1649977179
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1649977179
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1649977179
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1649977179
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1649977179
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1649977179
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1649977179
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1649977179
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1649977179
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1649977179
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1649977179
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1649977179
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1649977179
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1649977179
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1649977179
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1649977179
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1649977179
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1649977179
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1649977179
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1649977179
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_569
timestamp 1649977179
transform 1 0 53452 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_575
timestamp 1649977179
transform 1 0 54004 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_11
timestamp 1649977179
transform 1 0 2116 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_23
timestamp 1649977179
transform 1 0 3220 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_35
timestamp 1649977179
transform 1 0 4324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp 1649977179
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1649977179
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1649977179
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1649977179
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1649977179
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1649977179
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1649977179
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1649977179
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1649977179
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1649977179
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1649977179
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1649977179
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1649977179
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1649977179
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1649977179
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1649977179
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1649977179
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1649977179
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1649977179
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1649977179
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1649977179
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1649977179
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1649977179
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1649977179
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1649977179
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1649977179
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1649977179
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1649977179
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1649977179
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1649977179
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1649977179
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_561
timestamp 1649977179
transform 1 0 52716 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_564
timestamp 1649977179
transform 1 0 52992 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_572
timestamp 1649977179
transform 1 0 53728 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1649977179
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1649977179
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1649977179
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1649977179
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1649977179
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1649977179
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1649977179
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1649977179
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1649977179
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1649977179
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1649977179
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1649977179
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1649977179
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1649977179
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1649977179
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1649977179
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1649977179
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1649977179
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1649977179
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1649977179
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1649977179
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1649977179
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1649977179
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1649977179
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1649977179
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1649977179
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1649977179
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1649977179
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1649977179
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1649977179
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1649977179
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1649977179
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1649977179
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_569
timestamp 1649977179
transform 1 0 53452 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_575
timestamp 1649977179
transform 1 0 54004 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1649977179
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1649977179
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1649977179
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1649977179
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1649977179
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1649977179
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1649977179
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1649977179
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1649977179
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1649977179
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1649977179
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1649977179
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1649977179
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1649977179
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1649977179
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1649977179
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1649977179
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1649977179
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1649977179
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1649977179
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1649977179
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1649977179
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1649977179
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1649977179
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1649977179
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1649977179
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1649977179
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1649977179
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1649977179
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1649977179
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1649977179
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_573
timestamp 1649977179
transform 1 0 53820 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_7
timestamp 1649977179
transform 1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_13
timestamp 1649977179
transform 1 0 2300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_25
timestamp 1649977179
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1649977179
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1649977179
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1649977179
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1649977179
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1649977179
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1649977179
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1649977179
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1649977179
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1649977179
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1649977179
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1649977179
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1649977179
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1649977179
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1649977179
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1649977179
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1649977179
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1649977179
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1649977179
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1649977179
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1649977179
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1649977179
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1649977179
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1649977179
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1649977179
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1649977179
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1649977179
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1649977179
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1649977179
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1649977179
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1649977179
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1649977179
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1649977179
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_569
timestamp 1649977179
transform 1 0 53452 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_575
timestamp 1649977179
transform 1 0 54004 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1649977179
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1649977179
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1649977179
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1649977179
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1649977179
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1649977179
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1649977179
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1649977179
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1649977179
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1649977179
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1649977179
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1649977179
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1649977179
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1649977179
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1649977179
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1649977179
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1649977179
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1649977179
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1649977179
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1649977179
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1649977179
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1649977179
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1649977179
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1649977179
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1649977179
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1649977179
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1649977179
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1649977179
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1649977179
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1649977179
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_573
timestamp 1649977179
transform 1 0 53820 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1649977179
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1649977179
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1649977179
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1649977179
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1649977179
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1649977179
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1649977179
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1649977179
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1649977179
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1649977179
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1649977179
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1649977179
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1649977179
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1649977179
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1649977179
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1649977179
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1649977179
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1649977179
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1649977179
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1649977179
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1649977179
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1649977179
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1649977179
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1649977179
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1649977179
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1649977179
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1649977179
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1649977179
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1649977179
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1649977179
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1649977179
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_557
timestamp 1649977179
transform 1 0 52348 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_561
timestamp 1649977179
transform 1 0 52716 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_564
timestamp 1649977179
transform 1 0 52992 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_572
timestamp 1649977179
transform 1 0 53728 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_7
timestamp 1649977179
transform 1 0 1748 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_19
timestamp 1649977179
transform 1 0 2852 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_31
timestamp 1649977179
transform 1 0 3956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_43
timestamp 1649977179
transform 1 0 5060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1649977179
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1649977179
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1649977179
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1649977179
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1649977179
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1649977179
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1649977179
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1649977179
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1649977179
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1649977179
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1649977179
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1649977179
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1649977179
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1649977179
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1649977179
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1649977179
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1649977179
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1649977179
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1649977179
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1649977179
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1649977179
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1649977179
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1649977179
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1649977179
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1649977179
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1649977179
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1649977179
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1649977179
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1649977179
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1649977179
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1649977179
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1649977179
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1649977179
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_573
timestamp 1649977179
transform 1 0 53820 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_13
timestamp 1649977179
transform 1 0 2300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_25
timestamp 1649977179
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1649977179
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1649977179
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1649977179
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1649977179
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1649977179
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1649977179
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1649977179
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1649977179
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1649977179
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1649977179
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1649977179
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1649977179
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1649977179
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1649977179
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1649977179
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1649977179
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1649977179
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1649977179
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1649977179
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1649977179
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1649977179
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1649977179
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1649977179
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1649977179
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1649977179
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1649977179
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1649977179
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1649977179
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1649977179
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1649977179
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1649977179
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1649977179
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1649977179
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_569
timestamp 1649977179
transform 1 0 53452 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_575
timestamp 1649977179
transform 1 0 54004 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1649977179
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1649977179
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1649977179
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1649977179
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1649977179
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1649977179
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1649977179
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1649977179
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1649977179
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1649977179
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1649977179
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1649977179
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1649977179
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1649977179
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1649977179
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1649977179
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1649977179
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1649977179
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1649977179
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1649977179
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1649977179
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1649977179
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1649977179
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1649977179
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1649977179
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1649977179
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1649977179
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1649977179
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1649977179
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_561
timestamp 1649977179
transform 1 0 52716 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_564
timestamp 1649977179
transform 1 0 52992 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_572
timestamp 1649977179
transform 1 0 53728 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1649977179
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1649977179
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1649977179
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1649977179
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1649977179
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1649977179
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1649977179
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1649977179
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1649977179
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1649977179
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1649977179
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1649977179
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1649977179
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1649977179
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1649977179
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1649977179
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1649977179
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1649977179
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1649977179
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1649977179
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1649977179
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1649977179
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1649977179
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1649977179
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1649977179
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1649977179
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1649977179
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1649977179
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1649977179
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1649977179
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1649977179
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_569
timestamp 1649977179
transform 1 0 53452 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_575
timestamp 1649977179
transform 1 0 54004 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1649977179
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1649977179
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1649977179
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1649977179
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1649977179
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1649977179
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1649977179
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1649977179
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1649977179
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1649977179
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1649977179
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1649977179
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1649977179
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1649977179
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1649977179
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1649977179
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1649977179
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1649977179
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1649977179
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1649977179
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1649977179
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1649977179
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1649977179
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1649977179
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1649977179
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1649977179
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1649977179
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1649977179
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1649977179
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1649977179
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1649977179
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1649977179
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1649977179
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_573
timestamp 1649977179
transform 1 0 53820 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1649977179
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1649977179
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1649977179
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1649977179
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1649977179
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1649977179
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1649977179
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1649977179
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1649977179
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1649977179
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1649977179
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1649977179
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1649977179
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1649977179
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1649977179
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1649977179
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1649977179
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1649977179
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1649977179
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1649977179
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1649977179
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1649977179
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1649977179
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1649977179
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1649977179
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1649977179
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1649977179
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1649977179
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1649977179
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1649977179
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1649977179
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1649977179
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1649977179
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_569
timestamp 1649977179
transform 1 0 53452 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_575
timestamp 1649977179
transform 1 0 54004 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_7
timestamp 1649977179
transform 1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_13
timestamp 1649977179
transform 1 0 2300 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_25
timestamp 1649977179
transform 1 0 3404 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_37
timestamp 1649977179
transform 1 0 4508 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_49
timestamp 1649977179
transform 1 0 5612 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1649977179
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1649977179
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1649977179
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1649977179
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1649977179
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1649977179
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1649977179
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1649977179
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1649977179
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1649977179
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1649977179
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1649977179
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1649977179
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1649977179
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1649977179
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1649977179
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1649977179
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1649977179
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1649977179
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1649977179
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1649977179
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1649977179
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1649977179
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1649977179
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1649977179
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1649977179
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1649977179
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1649977179
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1649977179
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1649977179
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1649977179
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1649977179
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_561
timestamp 1649977179
transform 1 0 52716 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_564
timestamp 1649977179
transform 1 0 52992 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_572
timestamp 1649977179
transform 1 0 53728 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1649977179
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1649977179
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1649977179
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1649977179
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1649977179
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1649977179
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1649977179
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1649977179
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1649977179
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1649977179
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1649977179
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1649977179
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1649977179
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1649977179
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1649977179
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1649977179
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1649977179
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1649977179
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1649977179
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1649977179
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1649977179
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1649977179
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1649977179
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1649977179
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1649977179
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1649977179
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1649977179
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1649977179
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1649977179
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1649977179
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1649977179
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1649977179
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_569
timestamp 1649977179
transform 1 0 53452 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_575
timestamp 1649977179
transform 1 0 54004 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1649977179
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1649977179
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1649977179
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1649977179
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1649977179
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1649977179
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1649977179
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1649977179
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1649977179
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1649977179
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1649977179
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1649977179
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1649977179
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1649977179
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1649977179
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1649977179
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1649977179
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1649977179
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1649977179
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1649977179
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1649977179
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1649977179
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1649977179
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1649977179
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1649977179
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1649977179
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1649977179
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1649977179
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1649977179
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1649977179
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1649977179
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1649977179
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_573
timestamp 1649977179
transform 1 0 53820 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_5
timestamp 1649977179
transform 1 0 1564 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_17
timestamp 1649977179
transform 1 0 2668 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_25
timestamp 1649977179
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1649977179
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1649977179
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1649977179
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1649977179
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1649977179
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1649977179
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1649977179
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1649977179
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1649977179
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1649977179
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1649977179
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1649977179
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1649977179
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1649977179
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1649977179
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1649977179
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1649977179
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1649977179
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1649977179
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1649977179
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1649977179
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1649977179
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1649977179
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1649977179
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1649977179
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1649977179
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1649977179
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1649977179
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1649977179
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1649977179
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1649977179
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1649977179
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_569
timestamp 1649977179
transform 1 0 53452 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_575
timestamp 1649977179
transform 1 0 54004 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_7
timestamp 1649977179
transform 1 0 1748 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_19
timestamp 1649977179
transform 1 0 2852 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_31
timestamp 1649977179
transform 1 0 3956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_43
timestamp 1649977179
transform 1 0 5060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1649977179
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1649977179
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1649977179
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1649977179
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1649977179
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1649977179
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1649977179
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1649977179
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1649977179
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1649977179
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1649977179
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1649977179
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1649977179
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1649977179
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1649977179
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1649977179
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1649977179
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1649977179
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1649977179
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1649977179
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1649977179
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1649977179
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1649977179
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1649977179
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1649977179
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1649977179
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1649977179
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1649977179
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1649977179
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1649977179
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1649977179
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1649977179
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1649977179
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_573
timestamp 1649977179
transform 1 0 53820 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1649977179
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1649977179
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1649977179
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1649977179
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1649977179
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1649977179
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1649977179
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1649977179
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1649977179
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1649977179
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1649977179
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1649977179
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1649977179
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1649977179
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1649977179
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1649977179
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1649977179
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1649977179
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1649977179
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1649977179
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1649977179
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1649977179
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1649977179
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1649977179
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1649977179
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1649977179
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1649977179
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1649977179
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1649977179
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1649977179
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1649977179
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_557
timestamp 1649977179
transform 1 0 52348 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_561
timestamp 1649977179
transform 1 0 52716 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_564
timestamp 1649977179
transform 1 0 52992 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_572
timestamp 1649977179
transform 1 0 53728 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1649977179
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1649977179
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1649977179
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1649977179
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1649977179
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1649977179
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1649977179
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1649977179
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1649977179
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1649977179
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1649977179
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1649977179
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1649977179
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1649977179
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1649977179
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1649977179
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1649977179
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1649977179
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1649977179
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1649977179
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1649977179
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1649977179
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1649977179
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1649977179
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1649977179
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1649977179
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1649977179
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1649977179
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1649977179
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1649977179
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1649977179
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1649977179
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1649977179
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1649977179
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_573
timestamp 1649977179
transform 1 0 53820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_7
timestamp 1649977179
transform 1 0 1748 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_19
timestamp 1649977179
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1649977179
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1649977179
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1649977179
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1649977179
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1649977179
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1649977179
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1649977179
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1649977179
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1649977179
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1649977179
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1649977179
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1649977179
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1649977179
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1649977179
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1649977179
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1649977179
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1649977179
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1649977179
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1649977179
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1649977179
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1649977179
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1649977179
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1649977179
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1649977179
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1649977179
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1649977179
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1649977179
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1649977179
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1649977179
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1649977179
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1649977179
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1649977179
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1649977179
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1649977179
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_569
timestamp 1649977179
transform 1 0 53452 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_575
timestamp 1649977179
transform 1 0 54004 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_13
timestamp 1649977179
transform 1 0 2300 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_25
timestamp 1649977179
transform 1 0 3404 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_37
timestamp 1649977179
transform 1 0 4508 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_49
timestamp 1649977179
transform 1 0 5612 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1649977179
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1649977179
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1649977179
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1649977179
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1649977179
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1649977179
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1649977179
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1649977179
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1649977179
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1649977179
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1649977179
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1649977179
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1649977179
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1649977179
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1649977179
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1649977179
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1649977179
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1649977179
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1649977179
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1649977179
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1649977179
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1649977179
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1649977179
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1649977179
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1649977179
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1649977179
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1649977179
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1649977179
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1649977179
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1649977179
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1649977179
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1649977179
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_573
timestamp 1649977179
transform 1 0 53820 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1649977179
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1649977179
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1649977179
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1649977179
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1649977179
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1649977179
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1649977179
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1649977179
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1649977179
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1649977179
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1649977179
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1649977179
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1649977179
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1649977179
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1649977179
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1649977179
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1649977179
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1649977179
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1649977179
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1649977179
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1649977179
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1649977179
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1649977179
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1649977179
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1649977179
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1649977179
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1649977179
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1649977179
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1649977179
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1649977179
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1649977179
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1649977179
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_557
timestamp 1649977179
transform 1 0 52348 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_561
timestamp 1649977179
transform 1 0 52716 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_564
timestamp 1649977179
transform 1 0 52992 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_572
timestamp 1649977179
transform 1 0 53728 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1649977179
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1649977179
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1649977179
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1649977179
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1649977179
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1649977179
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1649977179
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1649977179
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1649977179
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1649977179
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1649977179
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1649977179
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1649977179
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1649977179
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1649977179
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1649977179
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1649977179
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1649977179
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1649977179
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1649977179
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1649977179
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1649977179
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1649977179
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1649977179
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1649977179
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1649977179
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1649977179
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1649977179
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1649977179
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1649977179
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1649977179
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1649977179
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1649977179
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_573
timestamp 1649977179
transform 1 0 53820 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1649977179
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1649977179
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1649977179
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1649977179
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1649977179
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1649977179
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1649977179
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1649977179
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1649977179
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1649977179
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1649977179
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1649977179
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1649977179
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1649977179
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1649977179
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1649977179
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1649977179
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1649977179
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1649977179
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1649977179
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1649977179
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1649977179
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1649977179
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1649977179
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1649977179
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1649977179
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1649977179
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1649977179
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1649977179
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1649977179
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1649977179
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1649977179
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1649977179
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1649977179
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_569
timestamp 1649977179
transform 1 0 53452 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_575
timestamp 1649977179
transform 1 0 54004 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_5
timestamp 1649977179
transform 1 0 1564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_17
timestamp 1649977179
transform 1 0 2668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_29
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_41
timestamp 1649977179
transform 1 0 4876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_53
timestamp 1649977179
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1649977179
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1649977179
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1649977179
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1649977179
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1649977179
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1649977179
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1649977179
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1649977179
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1649977179
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1649977179
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1649977179
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1649977179
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1649977179
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1649977179
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1649977179
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1649977179
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1649977179
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1649977179
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1649977179
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1649977179
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1649977179
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1649977179
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1649977179
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1649977179
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1649977179
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1649977179
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1649977179
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1649977179
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1649977179
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1649977179
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1649977179
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1649977179
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1649977179
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1649977179
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1649977179
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_573
timestamp 1649977179
transform 1 0 53820 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_7
timestamp 1649977179
transform 1 0 1748 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_19
timestamp 1649977179
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1649977179
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1649977179
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1649977179
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1649977179
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1649977179
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1649977179
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1649977179
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1649977179
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1649977179
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1649977179
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1649977179
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1649977179
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1649977179
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1649977179
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1649977179
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1649977179
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1649977179
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1649977179
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1649977179
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1649977179
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1649977179
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1649977179
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1649977179
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1649977179
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1649977179
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1649977179
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1649977179
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1649977179
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1649977179
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1649977179
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1649977179
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1649977179
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1649977179
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1649977179
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1649977179
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1649977179
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1649977179
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1649977179
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1649977179
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1649977179
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1649977179
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1649977179
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1649977179
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1649977179
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1649977179
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_569
timestamp 1649977179
transform 1 0 53452 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_575
timestamp 1649977179
transform 1 0 54004 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1649977179
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1649977179
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1649977179
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1649977179
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1649977179
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1649977179
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1649977179
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1649977179
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1649977179
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1649977179
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1649977179
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1649977179
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1649977179
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1649977179
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1649977179
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1649977179
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1649977179
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1649977179
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1649977179
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1649977179
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1649977179
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1649977179
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1649977179
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1649977179
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1649977179
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1649977179
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1649977179
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1649977179
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1649977179
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1649977179
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1649977179
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1649977179
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1649977179
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1649977179
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1649977179
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1649977179
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1649977179
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1649977179
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1649977179
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1649977179
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1649977179
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1649977179
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1649977179
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1649977179
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1649977179
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1649977179
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1649977179
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_561
timestamp 1649977179
transform 1 0 52716 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_564
timestamp 1649977179
transform 1 0 52992 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_572
timestamp 1649977179
transform 1 0 53728 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_5
timestamp 1649977179
transform 1 0 1564 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_17
timestamp 1649977179
transform 1 0 2668 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_25
timestamp 1649977179
transform 1 0 3404 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1649977179
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1649977179
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1649977179
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1649977179
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1649977179
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1649977179
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1649977179
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1649977179
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1649977179
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1649977179
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1649977179
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1649977179
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1649977179
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1649977179
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1649977179
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1649977179
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1649977179
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1649977179
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1649977179
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1649977179
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1649977179
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1649977179
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1649977179
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1649977179
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1649977179
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1649977179
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1649977179
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1649977179
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1649977179
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1649977179
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1649977179
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1649977179
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1649977179
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1649977179
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1649977179
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1649977179
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1649977179
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1649977179
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1649977179
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1649977179
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1649977179
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1649977179
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1649977179
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1649977179
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1649977179
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_569
timestamp 1649977179
transform 1 0 53452 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_575
timestamp 1649977179
transform 1 0 54004 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_9
timestamp 1649977179
transform 1 0 1932 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_21
timestamp 1649977179
transform 1 0 3036 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_33
timestamp 1649977179
transform 1 0 4140 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_45
timestamp 1649977179
transform 1 0 5244 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp 1649977179
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1649977179
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1649977179
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1649977179
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1649977179
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1649977179
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1649977179
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1649977179
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1649977179
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1649977179
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1649977179
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1649977179
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1649977179
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1649977179
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1649977179
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1649977179
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1649977179
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1649977179
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1649977179
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1649977179
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1649977179
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1649977179
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1649977179
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1649977179
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1649977179
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1649977179
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1649977179
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1649977179
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1649977179
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1649977179
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1649977179
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1649977179
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1649977179
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1649977179
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1649977179
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1649977179
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1649977179
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1649977179
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1649977179
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1649977179
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1649977179
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1649977179
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1649977179
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1649977179
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1649977179
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1649977179
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1649977179
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_573
timestamp 1649977179
transform 1 0 53820 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1649977179
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1649977179
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1649977179
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1649977179
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1649977179
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1649977179
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1649977179
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1649977179
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1649977179
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1649977179
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1649977179
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1649977179
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1649977179
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_209
timestamp 1649977179
transform 1 0 20332 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_217
timestamp 1649977179
transform 1 0 21068 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_229
timestamp 1649977179
transform 1 0 22172 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_241
timestamp 1649977179
transform 1 0 23276 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_249
timestamp 1649977179
transform 1 0 24012 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1649977179
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1649977179
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1649977179
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1649977179
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1649977179
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1649977179
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1649977179
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1649977179
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1649977179
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1649977179
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1649977179
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1649977179
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1649977179
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1649977179
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1649977179
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1649977179
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1649977179
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1649977179
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1649977179
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1649977179
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1649977179
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1649977179
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1649977179
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1649977179
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1649977179
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1649977179
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1649977179
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1649977179
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1649977179
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1649977179
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_569
timestamp 1649977179
transform 1 0 53452 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_575
timestamp 1649977179
transform 1 0 54004 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1649977179
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1649977179
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1649977179
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1649977179
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1649977179
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1649977179
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1649977179
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1649977179
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1649977179
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1649977179
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1649977179
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1649977179
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1649977179
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1649977179
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_205
timestamp 1649977179
transform 1 0 19964 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_208
timestamp 1649977179
transform 1 0 20240 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_215
timestamp 1649977179
transform 1 0 20884 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1649977179
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_227
timestamp 1649977179
transform 1 0 21988 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_239
timestamp 1649977179
transform 1 0 23092 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_251
timestamp 1649977179
transform 1 0 24196 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_263
timestamp 1649977179
transform 1 0 25300 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_275
timestamp 1649977179
transform 1 0 26404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1649977179
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1649977179
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_305
timestamp 1649977179
transform 1 0 29164 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_313
timestamp 1649977179
transform 1 0 29900 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_316
timestamp 1649977179
transform 1 0 30176 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_328
timestamp 1649977179
transform 1 0 31280 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1649977179
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1649977179
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1649977179
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1649977179
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1649977179
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1649977179
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1649977179
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1649977179
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1649977179
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1649977179
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1649977179
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1649977179
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1649977179
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1649977179
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1649977179
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1649977179
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1649977179
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1649977179
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1649977179
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1649977179
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1649977179
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1649977179
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1649977179
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_561
timestamp 1649977179
transform 1 0 52716 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_564
timestamp 1649977179
transform 1 0 52992 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_572
timestamp 1649977179
transform 1 0 53728 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1649977179
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1649977179
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1649977179
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1649977179
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1649977179
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1649977179
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1649977179
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1649977179
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1649977179
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1649977179
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1649977179
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1649977179
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1649977179
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1649977179
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1649977179
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_201
timestamp 1649977179
transform 1 0 19596 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_207
timestamp 1649977179
transform 1 0 20148 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_216
timestamp 1649977179
transform 1 0 20976 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_223
timestamp 1649977179
transform 1 0 21620 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_229
timestamp 1649977179
transform 1 0 22172 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_235
timestamp 1649977179
transform 1 0 22724 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_247
timestamp 1649977179
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1649977179
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1649977179
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_277
timestamp 1649977179
transform 1 0 26588 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_281
timestamp 1649977179
transform 1 0 26956 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_287
timestamp 1649977179
transform 1 0 27508 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_299
timestamp 1649977179
transform 1 0 28612 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1649977179
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_309
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_313
timestamp 1649977179
transform 1 0 29900 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_321
timestamp 1649977179
transform 1 0 30636 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_327
timestamp 1649977179
transform 1 0 31188 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_339
timestamp 1649977179
transform 1 0 32292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_351
timestamp 1649977179
transform 1 0 33396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1649977179
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1649977179
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1649977179
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1649977179
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1649977179
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1649977179
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1649977179
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1649977179
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1649977179
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1649977179
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1649977179
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1649977179
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1649977179
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1649977179
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1649977179
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1649977179
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1649977179
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1649977179
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1649977179
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1649977179
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1649977179
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_569
timestamp 1649977179
transform 1 0 53452 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_575
timestamp 1649977179
transform 1 0 54004 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_7
timestamp 1649977179
transform 1 0 1748 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_19
timestamp 1649977179
transform 1 0 2852 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_31
timestamp 1649977179
transform 1 0 3956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_43
timestamp 1649977179
transform 1 0 5060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1649977179
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1649977179
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1649977179
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1649977179
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1649977179
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1649977179
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1649977179
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1649977179
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1649977179
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1649977179
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1649977179
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_193
timestamp 1649977179
transform 1 0 18860 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_197
timestamp 1649977179
transform 1 0 19228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_200
timestamp 1649977179
transform 1 0 19504 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_209
timestamp 1649977179
transform 1 0 20332 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1649977179
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_228
timestamp 1649977179
transform 1 0 22080 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_240
timestamp 1649977179
transform 1 0 23184 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_252
timestamp 1649977179
transform 1 0 24288 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_256
timestamp 1649977179
transform 1 0 24656 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_260
timestamp 1649977179
transform 1 0 25024 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_263
timestamp 1649977179
transform 1 0 25300 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_269
timestamp 1649977179
transform 1 0 25852 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_272
timestamp 1649977179
transform 1 0 26128 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_283
timestamp 1649977179
transform 1 0 27140 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_289
timestamp 1649977179
transform 1 0 27692 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_295
timestamp 1649977179
transform 1 0 28244 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_303
timestamp 1649977179
transform 1 0 28980 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_306
timestamp 1649977179
transform 1 0 29256 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_317
timestamp 1649977179
transform 1 0 30268 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_328
timestamp 1649977179
transform 1 0 31280 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_339
timestamp 1649977179
transform 1 0 32292 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_351
timestamp 1649977179
transform 1 0 33396 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_363
timestamp 1649977179
transform 1 0 34500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_375
timestamp 1649977179
transform 1 0 35604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_387
timestamp 1649977179
transform 1 0 36708 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1649977179
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1649977179
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1649977179
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1649977179
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1649977179
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1649977179
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1649977179
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1649977179
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1649977179
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1649977179
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1649977179
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1649977179
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1649977179
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1649977179
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1649977179
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1649977179
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1649977179
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1649977179
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1649977179
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_573
timestamp 1649977179
transform 1 0 53820 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_11
timestamp 1649977179
transform 1 0 2116 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_23
timestamp 1649977179
transform 1 0 3220 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1649977179
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1649977179
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1649977179
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1649977179
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1649977179
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1649977179
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1649977179
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1649977179
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1649977179
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1649977179
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1649977179
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1649977179
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1649977179
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1649977179
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_201
timestamp 1649977179
transform 1 0 19596 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_208
timestamp 1649977179
transform 1 0 20240 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_219
timestamp 1649977179
transform 1 0 21252 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_225
timestamp 1649977179
transform 1 0 21804 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_239
timestamp 1649977179
transform 1 0 23092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1649977179
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_257
timestamp 1649977179
transform 1 0 24748 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_263
timestamp 1649977179
transform 1 0 25300 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_267
timestamp 1649977179
transform 1 0 25668 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_270
timestamp 1649977179
transform 1 0 25944 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_277
timestamp 1649977179
transform 1 0 26588 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_284
timestamp 1649977179
transform 1 0 27232 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_290
timestamp 1649977179
transform 1 0 27784 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_294
timestamp 1649977179
transform 1 0 28152 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_297
timestamp 1649977179
transform 1 0 28428 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_304
timestamp 1649977179
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_312
timestamp 1649977179
transform 1 0 29808 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_324
timestamp 1649977179
transform 1 0 30912 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_331
timestamp 1649977179
transform 1 0 31556 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_337
timestamp 1649977179
transform 1 0 32108 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_343
timestamp 1649977179
transform 1 0 32660 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_355
timestamp 1649977179
transform 1 0 33764 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1649977179
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1649977179
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1649977179
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1649977179
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1649977179
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1649977179
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1649977179
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1649977179
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1649977179
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1649977179
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1649977179
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1649977179
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1649977179
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1649977179
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1649977179
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1649977179
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1649977179
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1649977179
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1649977179
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1649977179
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_557
timestamp 1649977179
transform 1 0 52348 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_561
timestamp 1649977179
transform 1 0 52716 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_564
timestamp 1649977179
transform 1 0 52992 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_572
timestamp 1649977179
transform 1 0 53728 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1649977179
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1649977179
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1649977179
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1649977179
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1649977179
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1649977179
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1649977179
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1649977179
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1649977179
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1649977179
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1649977179
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1649977179
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1649977179
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1649977179
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1649977179
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1649977179
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_193
timestamp 1649977179
transform 1 0 18860 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_201
timestamp 1649977179
transform 1 0 19596 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_208
timestamp 1649977179
transform 1 0 20240 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_215
timestamp 1649977179
transform 1 0 20884 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1649977179
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_227
timestamp 1649977179
transform 1 0 21988 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_233
timestamp 1649977179
transform 1 0 22540 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_239
timestamp 1649977179
transform 1 0 23092 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_245
timestamp 1649977179
transform 1 0 23644 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_254
timestamp 1649977179
transform 1 0 24472 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_261
timestamp 1649977179
transform 1 0 25116 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_269
timestamp 1649977179
transform 1 0 25852 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_275
timestamp 1649977179
transform 1 0 26404 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1649977179
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_288
timestamp 1649977179
transform 1 0 27600 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_294
timestamp 1649977179
transform 1 0 28152 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_303
timestamp 1649977179
transform 1 0 28980 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_311
timestamp 1649977179
transform 1 0 29716 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_317
timestamp 1649977179
transform 1 0 30268 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_328
timestamp 1649977179
transform 1 0 31280 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_339
timestamp 1649977179
transform 1 0 32292 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_345
timestamp 1649977179
transform 1 0 32844 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_351
timestamp 1649977179
transform 1 0 33396 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_357
timestamp 1649977179
transform 1 0 33948 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_363
timestamp 1649977179
transform 1 0 34500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_375
timestamp 1649977179
transform 1 0 35604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_387
timestamp 1649977179
transform 1 0 36708 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1649977179
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1649977179
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1649977179
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1649977179
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1649977179
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1649977179
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1649977179
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1649977179
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1649977179
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1649977179
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1649977179
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1649977179
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1649977179
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1649977179
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1649977179
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1649977179
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1649977179
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1649977179
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1649977179
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_573
timestamp 1649977179
transform 1 0 53820 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1649977179
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1649977179
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1649977179
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1649977179
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1649977179
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1649977179
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1649977179
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1649977179
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1649977179
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1649977179
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1649977179
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1649977179
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1649977179
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1649977179
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1649977179
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1649977179
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_197
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_203
timestamp 1649977179
transform 1 0 19780 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_211
timestamp 1649977179
transform 1 0 20516 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_219
timestamp 1649977179
transform 1 0 21252 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_230
timestamp 1649977179
transform 1 0 22264 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_237
timestamp 1649977179
transform 1 0 22908 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_245
timestamp 1649977179
transform 1 0 23644 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1649977179
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_256
timestamp 1649977179
transform 1 0 24656 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_266
timestamp 1649977179
transform 1 0 25576 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_277
timestamp 1649977179
transform 1 0 26588 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_289
timestamp 1649977179
transform 1 0 27692 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_296
timestamp 1649977179
transform 1 0 28336 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_304
timestamp 1649977179
transform 1 0 29072 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_314
timestamp 1649977179
transform 1 0 29992 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_323
timestamp 1649977179
transform 1 0 30820 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_330
timestamp 1649977179
transform 1 0 31464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_336
timestamp 1649977179
transform 1 0 32016 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_342
timestamp 1649977179
transform 1 0 32568 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_348
timestamp 1649977179
transform 1 0 33120 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_354
timestamp 1649977179
transform 1 0 33672 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_360
timestamp 1649977179
transform 1 0 34224 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_367
timestamp 1649977179
transform 1 0 34868 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_373
timestamp 1649977179
transform 1 0 35420 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_376
timestamp 1649977179
transform 1 0 35696 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_382
timestamp 1649977179
transform 1 0 36248 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_394
timestamp 1649977179
transform 1 0 37352 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_406
timestamp 1649977179
transform 1 0 38456 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_418
timestamp 1649977179
transform 1 0 39560 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1649977179
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1649977179
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1649977179
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1649977179
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1649977179
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1649977179
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1649977179
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1649977179
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1649977179
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1649977179
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1649977179
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1649977179
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1649977179
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1649977179
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1649977179
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_569
timestamp 1649977179
transform 1 0 53452 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_575
timestamp 1649977179
transform 1 0 54004 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1649977179
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1649977179
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1649977179
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1649977179
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1649977179
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1649977179
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1649977179
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1649977179
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1649977179
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1649977179
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1649977179
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1649977179
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1649977179
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1649977179
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1649977179
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1649977179
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_193
timestamp 1649977179
transform 1 0 18860 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_201
timestamp 1649977179
transform 1 0 19596 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_205
timestamp 1649977179
transform 1 0 19964 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_211
timestamp 1649977179
transform 1 0 20516 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_215
timestamp 1649977179
transform 1 0 20884 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1649977179
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_235
timestamp 1649977179
transform 1 0 22724 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_241
timestamp 1649977179
transform 1 0 23276 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_247
timestamp 1649977179
transform 1 0 23828 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_254
timestamp 1649977179
transform 1 0 24472 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_260
timestamp 1649977179
transform 1 0 25024 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_266
timestamp 1649977179
transform 1 0 25576 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1649977179
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_287
timestamp 1649977179
transform 1 0 27508 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_295
timestamp 1649977179
transform 1 0 28244 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_301
timestamp 1649977179
transform 1 0 28796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_310
timestamp 1649977179
transform 1 0 29624 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_314
timestamp 1649977179
transform 1 0 29992 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_319
timestamp 1649977179
transform 1 0 30452 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_326
timestamp 1649977179
transform 1 0 31096 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_332
timestamp 1649977179
transform 1 0 31648 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_343
timestamp 1649977179
transform 1 0 32660 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_347
timestamp 1649977179
transform 1 0 33028 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_361
timestamp 1649977179
transform 1 0 34316 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_377
timestamp 1649977179
transform 1 0 35788 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_383
timestamp 1649977179
transform 1 0 36340 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1649977179
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1649977179
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1649977179
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1649977179
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1649977179
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1649977179
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1649977179
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1649977179
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1649977179
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1649977179
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1649977179
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1649977179
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1649977179
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1649977179
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1649977179
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1649977179
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1649977179
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1649977179
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1649977179
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_573
timestamp 1649977179
transform 1 0 53820 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_7
timestamp 1649977179
transform 1 0 1748 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_13
timestamp 1649977179
transform 1 0 2300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_25
timestamp 1649977179
transform 1 0 3404 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1649977179
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1649977179
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1649977179
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1649977179
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1649977179
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1649977179
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1649977179
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1649977179
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1649977179
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1649977179
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1649977179
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1649977179
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1649977179
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1649977179
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_205
timestamp 1649977179
transform 1 0 19964 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_211
timestamp 1649977179
transform 1 0 20516 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_214
timestamp 1649977179
transform 1 0 20792 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_225
timestamp 1649977179
transform 1 0 21804 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_238
timestamp 1649977179
transform 1 0 23000 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1649977179
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_258
timestamp 1649977179
transform 1 0 24840 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_270
timestamp 1649977179
transform 1 0 25944 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_279
timestamp 1649977179
transform 1 0 26772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_285
timestamp 1649977179
transform 1 0 27324 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_289
timestamp 1649977179
transform 1 0 27692 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_292
timestamp 1649977179
transform 1 0 27968 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 1649977179
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_311
timestamp 1649977179
transform 1 0 29716 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_322
timestamp 1649977179
transform 1 0 30728 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_331
timestamp 1649977179
transform 1 0 31556 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_351
timestamp 1649977179
transform 1 0 33396 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1649977179
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1649977179
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_374
timestamp 1649977179
transform 1 0 35512 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_380
timestamp 1649977179
transform 1 0 36064 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_386
timestamp 1649977179
transform 1 0 36616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_392
timestamp 1649977179
transform 1 0 37168 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_398
timestamp 1649977179
transform 1 0 37720 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_410
timestamp 1649977179
transform 1 0 38824 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_418
timestamp 1649977179
transform 1 0 39560 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1649977179
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1649977179
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1649977179
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1649977179
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1649977179
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1649977179
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1649977179
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1649977179
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1649977179
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1649977179
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1649977179
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1649977179
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1649977179
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1649977179
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1649977179
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_569
timestamp 1649977179
transform 1 0 53452 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_572
timestamp 1649977179
transform 1 0 53728 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1649977179
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1649977179
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1649977179
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1649977179
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1649977179
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1649977179
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1649977179
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1649977179
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1649977179
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1649977179
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1649977179
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1649977179
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1649977179
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1649977179
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1649977179
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1649977179
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1649977179
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_181
timestamp 1649977179
transform 1 0 17756 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_189
timestamp 1649977179
transform 1 0 18492 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_192
timestamp 1649977179
transform 1 0 18768 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_198
timestamp 1649977179
transform 1 0 19320 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_207
timestamp 1649977179
transform 1 0 20148 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_216
timestamp 1649977179
transform 1 0 20976 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_231
timestamp 1649977179
transform 1 0 22356 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_243
timestamp 1649977179
transform 1 0 23460 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_251
timestamp 1649977179
transform 1 0 24196 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_259
timestamp 1649977179
transform 1 0 24932 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_270
timestamp 1649977179
transform 1 0 25944 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1649977179
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_285
timestamp 1649977179
transform 1 0 27324 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_289
timestamp 1649977179
transform 1 0 27692 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_294
timestamp 1649977179
transform 1 0 28152 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_303
timestamp 1649977179
transform 1 0 28980 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_309
timestamp 1649977179
transform 1 0 29532 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_320
timestamp 1649977179
transform 1 0 30544 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1649977179
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_353
timestamp 1649977179
transform 1 0 33580 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_370
timestamp 1649977179
transform 1 0 35144 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_377
timestamp 1649977179
transform 1 0 35788 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_384
timestamp 1649977179
transform 1 0 36432 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_395
timestamp 1649977179
transform 1 0 37444 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_401
timestamp 1649977179
transform 1 0 37996 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_413
timestamp 1649977179
transform 1 0 39100 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_425
timestamp 1649977179
transform 1 0 40204 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_437
timestamp 1649977179
transform 1 0 41308 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_445
timestamp 1649977179
transform 1 0 42044 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1649977179
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1649977179
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1649977179
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1649977179
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1649977179
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1649977179
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1649977179
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1649977179
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1649977179
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1649977179
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1649977179
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1649977179
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_561
timestamp 1649977179
transform 1 0 52716 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_572
timestamp 1649977179
transform 1 0 53728 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1649977179
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1649977179
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1649977179
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1649977179
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1649977179
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1649977179
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1649977179
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1649977179
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1649977179
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1649977179
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1649977179
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1649977179
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1649977179
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1649977179
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_177
timestamp 1649977179
transform 1 0 17388 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_185
timestamp 1649977179
transform 1 0 18124 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1649977179
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_197
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_205
timestamp 1649977179
transform 1 0 19964 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_209
timestamp 1649977179
transform 1 0 20332 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_215
timestamp 1649977179
transform 1 0 20884 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_224
timestamp 1649977179
transform 1 0 21712 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_236
timestamp 1649977179
transform 1 0 22816 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1649977179
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1649977179
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_253
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_257
timestamp 1649977179
transform 1 0 24748 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_265
timestamp 1649977179
transform 1 0 25484 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_273
timestamp 1649977179
transform 1 0 26220 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_291
timestamp 1649977179
transform 1 0 27876 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1649977179
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1649977179
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_313
timestamp 1649977179
transform 1 0 29900 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_321
timestamp 1649977179
transform 1 0 30636 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_342
timestamp 1649977179
transform 1 0 32568 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_352
timestamp 1649977179
transform 1 0 33488 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_356
timestamp 1649977179
transform 1 0 33856 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_360
timestamp 1649977179
transform 1 0 34224 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_373
timestamp 1649977179
transform 1 0 35420 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_382
timestamp 1649977179
transform 1 0 36248 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_388
timestamp 1649977179
transform 1 0 36800 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_394
timestamp 1649977179
transform 1 0 37352 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_400
timestamp 1649977179
transform 1 0 37904 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_412
timestamp 1649977179
transform 1 0 39008 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1649977179
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1649977179
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1649977179
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1649977179
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1649977179
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1649977179
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1649977179
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1649977179
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1649977179
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1649977179
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1649977179
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1649977179
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1649977179
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1649977179
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1649977179
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_569
timestamp 1649977179
transform 1 0 53452 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_575
timestamp 1649977179
transform 1 0 54004 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_5
timestamp 1649977179
transform 1 0 1564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_17
timestamp 1649977179
transform 1 0 2668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_29
timestamp 1649977179
transform 1 0 3772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_41
timestamp 1649977179
transform 1 0 4876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 1649977179
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1649977179
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1649977179
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1649977179
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1649977179
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1649977179
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1649977179
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1649977179
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1649977179
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1649977179
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1649977179
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_169
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_177
timestamp 1649977179
transform 1 0 17388 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_180
timestamp 1649977179
transform 1 0 17664 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_186
timestamp 1649977179
transform 1 0 18216 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_192
timestamp 1649977179
transform 1 0 18768 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_199
timestamp 1649977179
transform 1 0 19412 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_208
timestamp 1649977179
transform 1 0 20240 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_216
timestamp 1649977179
transform 1 0 20976 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_234
timestamp 1649977179
transform 1 0 22632 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_242
timestamp 1649977179
transform 1 0 23368 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_246
timestamp 1649977179
transform 1 0 23736 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_249
timestamp 1649977179
transform 1 0 24012 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_255
timestamp 1649977179
transform 1 0 24564 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_264
timestamp 1649977179
transform 1 0 25392 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_275
timestamp 1649977179
transform 1 0 26404 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1649977179
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_284
timestamp 1649977179
transform 1 0 27232 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_290
timestamp 1649977179
transform 1 0 27784 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_296
timestamp 1649977179
transform 1 0 28336 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_314
timestamp 1649977179
transform 1 0 29992 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_320
timestamp 1649977179
transform 1 0 30544 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_323
timestamp 1649977179
transform 1 0 30820 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 1649977179
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_346
timestamp 1649977179
transform 1 0 32936 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_352
timestamp 1649977179
transform 1 0 33488 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_356
timestamp 1649977179
transform 1 0 33856 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_373
timestamp 1649977179
transform 1 0 35420 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1649977179
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1649977179
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1649977179
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1649977179
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1649977179
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1649977179
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1649977179
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1649977179
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1649977179
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1649977179
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1649977179
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1649977179
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1649977179
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1649977179
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1649977179
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1649977179
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1649977179
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1649977179
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1649977179
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1649977179
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1649977179
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_573
timestamp 1649977179
transform 1 0 53820 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_7
timestamp 1649977179
transform 1 0 1748 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_19
timestamp 1649977179
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1649977179
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1649977179
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1649977179
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1649977179
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1649977179
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1649977179
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1649977179
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1649977179
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1649977179
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1649977179
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1649977179
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1649977179
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1649977179
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_177
timestamp 1649977179
transform 1 0 17388 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_183
timestamp 1649977179
transform 1 0 17940 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_186
timestamp 1649977179
transform 1 0 18216 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_192
timestamp 1649977179
transform 1 0 18768 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_197
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_204
timestamp 1649977179
transform 1 0 19872 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_214
timestamp 1649977179
transform 1 0 20792 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_224
timestamp 1649977179
transform 1 0 21712 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_231
timestamp 1649977179
transform 1 0 22356 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_239
timestamp 1649977179
transform 1 0 23092 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_246
timestamp 1649977179
transform 1 0 23736 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_257
timestamp 1649977179
transform 1 0 24748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_267
timestamp 1649977179
transform 1 0 25668 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_273
timestamp 1649977179
transform 1 0 26220 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_296
timestamp 1649977179
transform 1 0 28336 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_300
timestamp 1649977179
transform 1 0 28704 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_304
timestamp 1649977179
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_311
timestamp 1649977179
transform 1 0 29716 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_317
timestamp 1649977179
transform 1 0 30268 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_323
timestamp 1649977179
transform 1 0 30820 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_331
timestamp 1649977179
transform 1 0 31556 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_341
timestamp 1649977179
transform 1 0 32476 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_348
timestamp 1649977179
transform 1 0 33120 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_354
timestamp 1649977179
transform 1 0 33672 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_360
timestamp 1649977179
transform 1 0 34224 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_378
timestamp 1649977179
transform 1 0 35880 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_388
timestamp 1649977179
transform 1 0 36800 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_400
timestamp 1649977179
transform 1 0 37904 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_412
timestamp 1649977179
transform 1 0 39008 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1649977179
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1649977179
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1649977179
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1649977179
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1649977179
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1649977179
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1649977179
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1649977179
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1649977179
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1649977179
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1649977179
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1649977179
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1649977179
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1649977179
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1649977179
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_569
timestamp 1649977179
transform 1 0 53452 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_575
timestamp 1649977179
transform 1 0 54004 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1649977179
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1649977179
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1649977179
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1649977179
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1649977179
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1649977179
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1649977179
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1649977179
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1649977179
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1649977179
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1649977179
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1649977179
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1649977179
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1649977179
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1649977179
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_181
timestamp 1649977179
transform 1 0 17756 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_184
timestamp 1649977179
transform 1 0 18032 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_192
timestamp 1649977179
transform 1 0 18768 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_198
timestamp 1649977179
transform 1 0 19320 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_204
timestamp 1649977179
transform 1 0 19872 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_210
timestamp 1649977179
transform 1 0 20424 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1649977179
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1649977179
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_228
timestamp 1649977179
transform 1 0 22080 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_236
timestamp 1649977179
transform 1 0 22816 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_240
timestamp 1649977179
transform 1 0 23184 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_247
timestamp 1649977179
transform 1 0 23828 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_254
timestamp 1649977179
transform 1 0 24472 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_263
timestamp 1649977179
transform 1 0 25300 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_272
timestamp 1649977179
transform 1 0 26128 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_300
timestamp 1649977179
transform 1 0 28704 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_312
timestamp 1649977179
transform 1 0 29808 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_324
timestamp 1649977179
transform 1 0 30912 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_327
timestamp 1649977179
transform 1 0 31188 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1649977179
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_354
timestamp 1649977179
transform 1 0 33672 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_360
timestamp 1649977179
transform 1 0 34224 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_51_372
timestamp 1649977179
transform 1 0 35328 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_380
timestamp 1649977179
transform 1 0 36064 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_384
timestamp 1649977179
transform 1 0 36432 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_395
timestamp 1649977179
transform 1 0 37444 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_407
timestamp 1649977179
transform 1 0 38548 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_419
timestamp 1649977179
transform 1 0 39652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_431
timestamp 1649977179
transform 1 0 40756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_443
timestamp 1649977179
transform 1 0 41860 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1649977179
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1649977179
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1649977179
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1649977179
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1649977179
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1649977179
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1649977179
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1649977179
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1649977179
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1649977179
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1649977179
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1649977179
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1649977179
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_561
timestamp 1649977179
transform 1 0 52716 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_564
timestamp 1649977179
transform 1 0 52992 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_572
timestamp 1649977179
transform 1 0 53728 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1649977179
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1649977179
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1649977179
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1649977179
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1649977179
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1649977179
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1649977179
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1649977179
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1649977179
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1649977179
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1649977179
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1649977179
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1649977179
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1649977179
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_165
timestamp 1649977179
transform 1 0 16284 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_171
timestamp 1649977179
transform 1 0 16836 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_174
timestamp 1649977179
transform 1 0 17112 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_180
timestamp 1649977179
transform 1 0 17664 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_191
timestamp 1649977179
transform 1 0 18676 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1649977179
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_197
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_200
timestamp 1649977179
transform 1 0 19504 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_210
timestamp 1649977179
transform 1 0 20424 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_218
timestamp 1649977179
transform 1 0 21160 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_225
timestamp 1649977179
transform 1 0 21804 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_233
timestamp 1649977179
transform 1 0 22540 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_236
timestamp 1649977179
transform 1 0 22816 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_244
timestamp 1649977179
transform 1 0 23552 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_260
timestamp 1649977179
transform 1 0 25024 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_268
timestamp 1649977179
transform 1 0 25760 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_273
timestamp 1649977179
transform 1 0 26220 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_279
timestamp 1649977179
transform 1 0 26772 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_285
timestamp 1649977179
transform 1 0 27324 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_291
timestamp 1649977179
transform 1 0 27876 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_297
timestamp 1649977179
transform 1 0 28428 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_305
timestamp 1649977179
transform 1 0 29164 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_328
timestamp 1649977179
transform 1 0 31280 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_334
timestamp 1649977179
transform 1 0 31832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_340
timestamp 1649977179
transform 1 0 32384 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_346
timestamp 1649977179
transform 1 0 32936 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1649977179
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1649977179
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_367
timestamp 1649977179
transform 1 0 34868 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_373
timestamp 1649977179
transform 1 0 35420 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_377
timestamp 1649977179
transform 1 0 35788 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_388
timestamp 1649977179
transform 1 0 36800 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_394
timestamp 1649977179
transform 1 0 37352 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_400
timestamp 1649977179
transform 1 0 37904 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_412
timestamp 1649977179
transform 1 0 39008 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1649977179
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1649977179
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1649977179
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1649977179
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1649977179
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1649977179
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1649977179
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1649977179
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1649977179
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1649977179
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1649977179
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1649977179
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1649977179
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1649977179
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1649977179
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_569
timestamp 1649977179
transform 1 0 53452 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_575
timestamp 1649977179
transform 1 0 54004 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1649977179
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1649977179
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1649977179
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1649977179
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1649977179
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1649977179
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1649977179
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1649977179
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1649977179
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1649977179
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1649977179
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1649977179
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1649977179
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_161
timestamp 1649977179
transform 1 0 15916 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_164
timestamp 1649977179
transform 1 0 16192 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_169
timestamp 1649977179
transform 1 0 16652 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_175
timestamp 1649977179
transform 1 0 17204 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_182
timestamp 1649977179
transform 1 0 17848 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_194
timestamp 1649977179
transform 1 0 18952 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_205
timestamp 1649977179
transform 1 0 19964 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_216
timestamp 1649977179
transform 1 0 20976 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_225
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_229
timestamp 1649977179
transform 1 0 22172 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_237
timestamp 1649977179
transform 1 0 22908 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_250
timestamp 1649977179
transform 1 0 24104 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_257
timestamp 1649977179
transform 1 0 24748 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_263
timestamp 1649977179
transform 1 0 25300 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_271
timestamp 1649977179
transform 1 0 26036 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1649977179
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_300
timestamp 1649977179
transform 1 0 28704 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_306
timestamp 1649977179
transform 1 0 29256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_310
timestamp 1649977179
transform 1 0 29624 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_316
timestamp 1649977179
transform 1 0 30176 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_324
timestamp 1649977179
transform 1 0 30912 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_332
timestamp 1649977179
transform 1 0 31648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_342
timestamp 1649977179
transform 1 0 32568 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_351
timestamp 1649977179
transform 1 0 33396 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_363
timestamp 1649977179
transform 1 0 34500 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_374
timestamp 1649977179
transform 1 0 35512 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1649977179
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1649977179
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_399
timestamp 1649977179
transform 1 0 37812 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1649977179
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1649977179
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1649977179
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1649977179
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1649977179
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1649977179
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1649977179
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1649977179
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1649977179
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1649977179
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1649977179
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1649977179
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1649977179
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1649977179
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1649977179
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1649977179
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1649977179
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1649977179
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_573
timestamp 1649977179
transform 1 0 53820 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1649977179
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1649977179
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1649977179
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1649977179
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1649977179
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1649977179
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1649977179
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1649977179
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1649977179
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1649977179
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1649977179
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1649977179
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_153
timestamp 1649977179
transform 1 0 15180 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_158
timestamp 1649977179
transform 1 0 15640 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_164
timestamp 1649977179
transform 1 0 16192 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_171
timestamp 1649977179
transform 1 0 16836 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_180
timestamp 1649977179
transform 1 0 17664 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_190
timestamp 1649977179
transform 1 0 18584 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_54_202
timestamp 1649977179
transform 1 0 19688 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_214
timestamp 1649977179
transform 1 0 20792 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_218
timestamp 1649977179
transform 1 0 21160 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_224
timestamp 1649977179
transform 1 0 21712 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_233
timestamp 1649977179
transform 1 0 22540 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_239
timestamp 1649977179
transform 1 0 23092 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_244
timestamp 1649977179
transform 1 0 23552 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_54_260
timestamp 1649977179
transform 1 0 25024 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_270
timestamp 1649977179
transform 1 0 25944 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_276
timestamp 1649977179
transform 1 0 26496 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_282
timestamp 1649977179
transform 1 0 27048 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_294
timestamp 1649977179
transform 1 0 28152 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1649977179
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_309
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_312
timestamp 1649977179
transform 1 0 29808 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_323
timestamp 1649977179
transform 1 0 30820 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_334
timestamp 1649977179
transform 1 0 31832 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_343
timestamp 1649977179
transform 1 0 32660 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_350
timestamp 1649977179
transform 1 0 33304 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_360
timestamp 1649977179
transform 1 0 34224 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_367
timestamp 1649977179
transform 1 0 34868 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_373
timestamp 1649977179
transform 1 0 35420 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_389
timestamp 1649977179
transform 1 0 36892 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_401
timestamp 1649977179
transform 1 0 37996 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_407
timestamp 1649977179
transform 1 0 38548 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1649977179
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1649977179
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1649977179
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1649977179
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1649977179
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1649977179
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1649977179
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1649977179
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1649977179
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1649977179
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1649977179
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1649977179
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1649977179
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1649977179
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1649977179
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1649977179
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_569
timestamp 1649977179
transform 1 0 53452 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_575
timestamp 1649977179
transform 1 0 54004 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_7
timestamp 1649977179
transform 1 0 1748 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_13
timestamp 1649977179
transform 1 0 2300 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_25
timestamp 1649977179
transform 1 0 3404 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_37
timestamp 1649977179
transform 1 0 4508 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_49
timestamp 1649977179
transform 1 0 5612 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1649977179
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1649977179
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1649977179
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1649977179
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1649977179
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1649977179
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1649977179
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1649977179
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1649977179
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1649977179
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1649977179
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1649977179
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_173
timestamp 1649977179
transform 1 0 17020 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_181
timestamp 1649977179
transform 1 0 17756 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_190
timestamp 1649977179
transform 1 0 18584 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_199
timestamp 1649977179
transform 1 0 19412 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_207
timestamp 1649977179
transform 1 0 20148 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_211
timestamp 1649977179
transform 1 0 20516 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_219
timestamp 1649977179
transform 1 0 21252 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1649977179
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_225
timestamp 1649977179
transform 1 0 21804 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_229
timestamp 1649977179
transform 1 0 22172 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_236
timestamp 1649977179
transform 1 0 22816 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_247
timestamp 1649977179
transform 1 0 23828 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_257
timestamp 1649977179
transform 1 0 24748 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_268
timestamp 1649977179
transform 1 0 25760 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_274
timestamp 1649977179
transform 1 0 26312 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_283
timestamp 1649977179
transform 1 0 27140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_295
timestamp 1649977179
transform 1 0 28244 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_299
timestamp 1649977179
transform 1 0 28612 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_305
timestamp 1649977179
transform 1 0 29164 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_312
timestamp 1649977179
transform 1 0 29808 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_324
timestamp 1649977179
transform 1 0 30912 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_332
timestamp 1649977179
transform 1 0 31648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_341
timestamp 1649977179
transform 1 0 32476 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_349
timestamp 1649977179
transform 1 0 33212 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_355
timestamp 1649977179
transform 1 0 33764 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_361
timestamp 1649977179
transform 1 0 34316 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_367
timestamp 1649977179
transform 1 0 34868 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_378
timestamp 1649977179
transform 1 0 35880 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1649977179
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1649977179
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_398
timestamp 1649977179
transform 1 0 37720 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_404
timestamp 1649977179
transform 1 0 38272 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_410
timestamp 1649977179
transform 1 0 38824 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_422
timestamp 1649977179
transform 1 0 39928 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_434
timestamp 1649977179
transform 1 0 41032 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_446
timestamp 1649977179
transform 1 0 42136 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1649977179
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1649977179
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1649977179
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1649977179
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1649977179
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1649977179
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1649977179
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1649977179
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1649977179
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1649977179
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1649977179
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1649977179
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_561
timestamp 1649977179
transform 1 0 52716 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_564
timestamp 1649977179
transform 1 0 52992 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_572
timestamp 1649977179
transform 1 0 53728 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1649977179
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1649977179
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1649977179
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1649977179
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1649977179
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1649977179
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1649977179
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1649977179
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1649977179
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1649977179
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1649977179
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1649977179
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1649977179
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_165
timestamp 1649977179
transform 1 0 16284 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_56_173
timestamp 1649977179
transform 1 0 17020 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_181
timestamp 1649977179
transform 1 0 17756 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_188
timestamp 1649977179
transform 1 0 18400 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_202
timestamp 1649977179
transform 1 0 19688 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_209
timestamp 1649977179
transform 1 0 20332 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_213
timestamp 1649977179
transform 1 0 20700 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_216
timestamp 1649977179
transform 1 0 20976 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_222
timestamp 1649977179
transform 1 0 21528 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_231
timestamp 1649977179
transform 1 0 22356 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_242
timestamp 1649977179
transform 1 0 23368 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_248
timestamp 1649977179
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_260
timestamp 1649977179
transform 1 0 25024 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_272
timestamp 1649977179
transform 1 0 26128 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_293
timestamp 1649977179
transform 1 0 28060 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_304
timestamp 1649977179
transform 1 0 29072 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_311
timestamp 1649977179
transform 1 0 29716 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_320
timestamp 1649977179
transform 1 0 30544 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_329
timestamp 1649977179
transform 1 0 31372 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_342
timestamp 1649977179
transform 1 0 32568 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_348
timestamp 1649977179
transform 1 0 33120 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_354
timestamp 1649977179
transform 1 0 33672 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_360
timestamp 1649977179
transform 1 0 34224 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_373
timestamp 1649977179
transform 1 0 35420 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_382
timestamp 1649977179
transform 1 0 36248 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_389
timestamp 1649977179
transform 1 0 36892 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_395
timestamp 1649977179
transform 1 0 37444 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_401
timestamp 1649977179
transform 1 0 37996 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_407
timestamp 1649977179
transform 1 0 38548 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1649977179
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1649977179
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_423
timestamp 1649977179
transform 1 0 40020 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_429
timestamp 1649977179
transform 1 0 40572 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_441
timestamp 1649977179
transform 1 0 41676 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_453
timestamp 1649977179
transform 1 0 42780 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_465
timestamp 1649977179
transform 1 0 43884 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_473
timestamp 1649977179
transform 1 0 44620 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1649977179
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1649977179
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1649977179
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1649977179
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1649977179
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1649977179
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1649977179
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1649977179
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1649977179
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_569
timestamp 1649977179
transform 1 0 53452 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_575
timestamp 1649977179
transform 1 0 54004 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1649977179
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1649977179
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1649977179
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1649977179
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1649977179
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1649977179
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1649977179
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1649977179
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1649977179
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1649977179
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1649977179
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1649977179
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1649977179
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1649977179
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1649977179
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_169
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_173
timestamp 1649977179
transform 1 0 17020 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_179
timestamp 1649977179
transform 1 0 17572 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_186
timestamp 1649977179
transform 1 0 18216 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_192
timestamp 1649977179
transform 1 0 18768 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_195
timestamp 1649977179
transform 1 0 19044 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_201
timestamp 1649977179
transform 1 0 19596 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_207
timestamp 1649977179
transform 1 0 20148 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_211
timestamp 1649977179
transform 1 0 20516 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_214
timestamp 1649977179
transform 1 0 20792 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1649977179
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_227
timestamp 1649977179
transform 1 0 21988 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_231
timestamp 1649977179
transform 1 0 22356 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_235
timestamp 1649977179
transform 1 0 22724 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_245
timestamp 1649977179
transform 1 0 23644 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_251
timestamp 1649977179
transform 1 0 24196 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_255
timestamp 1649977179
transform 1 0 24564 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_258
timestamp 1649977179
transform 1 0 24840 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_264
timestamp 1649977179
transform 1 0 25392 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_270
timestamp 1649977179
transform 1 0 25944 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_276
timestamp 1649977179
transform 1 0 26496 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_288
timestamp 1649977179
transform 1 0 27600 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_294
timestamp 1649977179
transform 1 0 28152 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_303
timestamp 1649977179
transform 1 0 28980 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_315
timestamp 1649977179
transform 1 0 30084 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_324
timestamp 1649977179
transform 1 0 30912 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_331
timestamp 1649977179
transform 1 0 31556 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1649977179
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_339
timestamp 1649977179
transform 1 0 32292 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_347
timestamp 1649977179
transform 1 0 33028 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_353
timestamp 1649977179
transform 1 0 33580 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_357
timestamp 1649977179
transform 1 0 33948 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_365
timestamp 1649977179
transform 1 0 34684 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_374
timestamp 1649977179
transform 1 0 35512 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_383
timestamp 1649977179
transform 1 0 36340 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1649977179
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_400
timestamp 1649977179
transform 1 0 37904 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_408
timestamp 1649977179
transform 1 0 38640 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_414
timestamp 1649977179
transform 1 0 39192 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_423
timestamp 1649977179
transform 1 0 40020 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_429
timestamp 1649977179
transform 1 0 40572 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_435
timestamp 1649977179
transform 1 0 41124 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1649977179
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1649977179
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1649977179
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1649977179
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1649977179
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1649977179
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1649977179
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1649977179
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1649977179
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1649977179
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1649977179
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1649977179
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1649977179
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1649977179
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_573
timestamp 1649977179
transform 1 0 53820 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_3
timestamp 1649977179
transform 1 0 1380 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_7
timestamp 1649977179
transform 1 0 1748 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_19
timestamp 1649977179
transform 1 0 2852 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1649977179
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1649977179
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1649977179
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1649977179
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1649977179
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1649977179
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1649977179
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1649977179
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1649977179
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1649977179
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1649977179
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1649977179
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1649977179
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_167
timestamp 1649977179
transform 1 0 16468 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_173
timestamp 1649977179
transform 1 0 17020 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_179
timestamp 1649977179
transform 1 0 17572 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_188
timestamp 1649977179
transform 1 0 18400 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_199
timestamp 1649977179
transform 1 0 19412 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_207
timestamp 1649977179
transform 1 0 20148 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_217
timestamp 1649977179
transform 1 0 21068 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_223
timestamp 1649977179
transform 1 0 21620 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_230
timestamp 1649977179
transform 1 0 22264 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_237
timestamp 1649977179
transform 1 0 22908 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_248
timestamp 1649977179
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_253
timestamp 1649977179
transform 1 0 24380 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_256
timestamp 1649977179
transform 1 0 24656 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_267
timestamp 1649977179
transform 1 0 25668 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_276
timestamp 1649977179
transform 1 0 26496 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_284
timestamp 1649977179
transform 1 0 27232 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_292
timestamp 1649977179
transform 1 0 27968 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_303
timestamp 1649977179
transform 1 0 28980 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1649977179
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_316
timestamp 1649977179
transform 1 0 30176 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_322
timestamp 1649977179
transform 1 0 30728 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_332
timestamp 1649977179
transform 1 0 31648 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_340
timestamp 1649977179
transform 1 0 32384 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_346
timestamp 1649977179
transform 1 0 32936 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_360
timestamp 1649977179
transform 1 0 34224 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_372
timestamp 1649977179
transform 1 0 35328 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_381
timestamp 1649977179
transform 1 0 36156 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_387
timestamp 1649977179
transform 1 0 36708 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_393
timestamp 1649977179
transform 1 0 37260 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_399
timestamp 1649977179
transform 1 0 37812 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_405
timestamp 1649977179
transform 1 0 38364 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_411
timestamp 1649977179
transform 1 0 38916 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1649977179
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_423
timestamp 1649977179
transform 1 0 40020 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_435
timestamp 1649977179
transform 1 0 41124 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_447
timestamp 1649977179
transform 1 0 42228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_459
timestamp 1649977179
transform 1 0 43332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_471
timestamp 1649977179
transform 1 0 44436 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1649977179
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1649977179
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1649977179
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1649977179
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1649977179
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1649977179
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1649977179
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1649977179
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1649977179
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1649977179
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_569
timestamp 1649977179
transform 1 0 53452 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_575
timestamp 1649977179
transform 1 0 54004 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_3
timestamp 1649977179
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_11
timestamp 1649977179
transform 1 0 2116 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_23
timestamp 1649977179
transform 1 0 3220 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_35
timestamp 1649977179
transform 1 0 4324 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_47
timestamp 1649977179
transform 1 0 5428 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1649977179
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1649977179
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1649977179
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1649977179
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1649977179
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1649977179
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1649977179
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1649977179
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_149
timestamp 1649977179
transform 1 0 14812 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_155
timestamp 1649977179
transform 1 0 15364 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_158
timestamp 1649977179
transform 1 0 15640 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_164
timestamp 1649977179
transform 1 0 16192 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_171
timestamp 1649977179
transform 1 0 16836 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_180
timestamp 1649977179
transform 1 0 17664 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_189
timestamp 1649977179
transform 1 0 18492 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_198
timestamp 1649977179
transform 1 0 19320 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_209
timestamp 1649977179
transform 1 0 20332 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_215
timestamp 1649977179
transform 1 0 20884 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_220
timestamp 1649977179
transform 1 0 21344 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_225
timestamp 1649977179
transform 1 0 21804 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_234
timestamp 1649977179
transform 1 0 22632 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_242
timestamp 1649977179
transform 1 0 23368 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_245
timestamp 1649977179
transform 1 0 23644 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_251
timestamp 1649977179
transform 1 0 24196 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_257
timestamp 1649977179
transform 1 0 24748 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_269
timestamp 1649977179
transform 1 0 25852 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_273
timestamp 1649977179
transform 1 0 26220 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_276
timestamp 1649977179
transform 1 0 26496 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_284
timestamp 1649977179
transform 1 0 27232 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_292
timestamp 1649977179
transform 1 0 27968 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_295
timestamp 1649977179
transform 1 0 28244 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_306
timestamp 1649977179
transform 1 0 29256 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_317
timestamp 1649977179
transform 1 0 30268 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_324
timestamp 1649977179
transform 1 0 30912 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_332
timestamp 1649977179
transform 1 0 31648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_345
timestamp 1649977179
transform 1 0 32844 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_354
timestamp 1649977179
transform 1 0 33672 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_358
timestamp 1649977179
transform 1 0 34040 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_366
timestamp 1649977179
transform 1 0 34776 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_373
timestamp 1649977179
transform 1 0 35420 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_380
timestamp 1649977179
transform 1 0 36064 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_386
timestamp 1649977179
transform 1 0 36616 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_393
timestamp 1649977179
transform 1 0 37260 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_397
timestamp 1649977179
transform 1 0 37628 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_403
timestamp 1649977179
transform 1 0 38180 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_409
timestamp 1649977179
transform 1 0 38732 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_415
timestamp 1649977179
transform 1 0 39284 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_427
timestamp 1649977179
transform 1 0 40388 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_439
timestamp 1649977179
transform 1 0 41492 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1649977179
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1649977179
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1649977179
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1649977179
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1649977179
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1649977179
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1649977179
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1649977179
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1649977179
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1649977179
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1649977179
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1649977179
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1649977179
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1649977179
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_573
timestamp 1649977179
transform 1 0 53820 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1649977179
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1649977179
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1649977179
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1649977179
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1649977179
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1649977179
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1649977179
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1649977179
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1649977179
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1649977179
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1649977179
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1649977179
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1649977179
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1649977179
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_153
timestamp 1649977179
transform 1 0 15180 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_161
timestamp 1649977179
transform 1 0 15916 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_167
timestamp 1649977179
transform 1 0 16468 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_174
timestamp 1649977179
transform 1 0 17112 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_185
timestamp 1649977179
transform 1 0 18124 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_192
timestamp 1649977179
transform 1 0 18768 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1649977179
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_207
timestamp 1649977179
transform 1 0 20148 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_213
timestamp 1649977179
transform 1 0 20700 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_220
timestamp 1649977179
transform 1 0 21344 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_229
timestamp 1649977179
transform 1 0 22172 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_238
timestamp 1649977179
transform 1 0 23000 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_248
timestamp 1649977179
transform 1 0 23920 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_253
timestamp 1649977179
transform 1 0 24380 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_260
timestamp 1649977179
transform 1 0 25024 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_264
timestamp 1649977179
transform 1 0 25392 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_267
timestamp 1649977179
transform 1 0 25668 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_273
timestamp 1649977179
transform 1 0 26220 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_296
timestamp 1649977179
transform 1 0 28336 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_302
timestamp 1649977179
transform 1 0 28888 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_309
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_314
timestamp 1649977179
transform 1 0 29992 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_318
timestamp 1649977179
transform 1 0 30360 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_336
timestamp 1649977179
transform 1 0 32016 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1649977179
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1649977179
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_369
timestamp 1649977179
transform 1 0 35052 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_376
timestamp 1649977179
transform 1 0 35696 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_382
timestamp 1649977179
transform 1 0 36248 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_388
timestamp 1649977179
transform 1 0 36800 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_394
timestamp 1649977179
transform 1 0 37352 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_400
timestamp 1649977179
transform 1 0 37904 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_406
timestamp 1649977179
transform 1 0 38456 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_412
timestamp 1649977179
transform 1 0 39008 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_423
timestamp 1649977179
transform 1 0 40020 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_435
timestamp 1649977179
transform 1 0 41124 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_447
timestamp 1649977179
transform 1 0 42228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_459
timestamp 1649977179
transform 1 0 43332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_471
timestamp 1649977179
transform 1 0 44436 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1649977179
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1649977179
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1649977179
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1649977179
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1649977179
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1649977179
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1649977179
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1649977179
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1649977179
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_557
timestamp 1649977179
transform 1 0 52348 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_561
timestamp 1649977179
transform 1 0 52716 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_564
timestamp 1649977179
transform 1 0 52992 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_572
timestamp 1649977179
transform 1 0 53728 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1649977179
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_7
timestamp 1649977179
transform 1 0 1748 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_19
timestamp 1649977179
transform 1 0 2852 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_31
timestamp 1649977179
transform 1 0 3956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_43
timestamp 1649977179
transform 1 0 5060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1649977179
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1649977179
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1649977179
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1649977179
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1649977179
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1649977179
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1649977179
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1649977179
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1649977179
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1649977179
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1649977179
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_161
timestamp 1649977179
transform 1 0 15916 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_164
timestamp 1649977179
transform 1 0 16192 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_169
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_173
timestamp 1649977179
transform 1 0 17020 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_180
timestamp 1649977179
transform 1 0 17664 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_190
timestamp 1649977179
transform 1 0 18584 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_194
timestamp 1649977179
transform 1 0 18952 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_199
timestamp 1649977179
transform 1 0 19412 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_208
timestamp 1649977179
transform 1 0 20240 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_220
timestamp 1649977179
transform 1 0 21344 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_232
timestamp 1649977179
transform 1 0 22448 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_238
timestamp 1649977179
transform 1 0 23000 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_244
timestamp 1649977179
transform 1 0 23552 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_255
timestamp 1649977179
transform 1 0 24564 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_263
timestamp 1649977179
transform 1 0 25300 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_275
timestamp 1649977179
transform 1 0 26404 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1649977179
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_286
timestamp 1649977179
transform 1 0 27416 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_294
timestamp 1649977179
transform 1 0 28152 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_298
timestamp 1649977179
transform 1 0 28520 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_319
timestamp 1649977179
transform 1 0 30452 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_325
timestamp 1649977179
transform 1 0 31004 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_331
timestamp 1649977179
transform 1 0 31556 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1649977179
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_345
timestamp 1649977179
transform 1 0 32844 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_351
timestamp 1649977179
transform 1 0 33396 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_362
timestamp 1649977179
transform 1 0 34408 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_373
timestamp 1649977179
transform 1 0 35420 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_379
timestamp 1649977179
transform 1 0 35972 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_383
timestamp 1649977179
transform 1 0 36340 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_388
timestamp 1649977179
transform 1 0 36800 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_398
timestamp 1649977179
transform 1 0 37720 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_405
timestamp 1649977179
transform 1 0 38364 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_412
timestamp 1649977179
transform 1 0 39008 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_418
timestamp 1649977179
transform 1 0 39560 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_424
timestamp 1649977179
transform 1 0 40112 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_430
timestamp 1649977179
transform 1 0 40664 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_442
timestamp 1649977179
transform 1 0 41768 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1649977179
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1649977179
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1649977179
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1649977179
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1649977179
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1649977179
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1649977179
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1649977179
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1649977179
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1649977179
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1649977179
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1649977179
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1649977179
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_573
timestamp 1649977179
transform 1 0 53820 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_3
timestamp 1649977179
transform 1 0 1380 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_11
timestamp 1649977179
transform 1 0 2116 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_23
timestamp 1649977179
transform 1 0 3220 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1649977179
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1649977179
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1649977179
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1649977179
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1649977179
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1649977179
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1649977179
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1649977179
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1649977179
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1649977179
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1649977179
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1649977179
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1649977179
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_165
timestamp 1649977179
transform 1 0 16284 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_169
timestamp 1649977179
transform 1 0 16652 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_175
timestamp 1649977179
transform 1 0 17204 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_187
timestamp 1649977179
transform 1 0 18308 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1649977179
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_201
timestamp 1649977179
transform 1 0 19596 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_209
timestamp 1649977179
transform 1 0 20332 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_215
timestamp 1649977179
transform 1 0 20884 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_224
timestamp 1649977179
transform 1 0 21712 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_231
timestamp 1649977179
transform 1 0 22356 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_239
timestamp 1649977179
transform 1 0 23092 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_248
timestamp 1649977179
transform 1 0 23920 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1649977179
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_258
timestamp 1649977179
transform 1 0 24840 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_281
timestamp 1649977179
transform 1 0 26956 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_304
timestamp 1649977179
transform 1 0 29072 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_316
timestamp 1649977179
transform 1 0 30176 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_327
timestamp 1649977179
transform 1 0 31188 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_333
timestamp 1649977179
transform 1 0 31740 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_339
timestamp 1649977179
transform 1 0 32292 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_347
timestamp 1649977179
transform 1 0 33028 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_360
timestamp 1649977179
transform 1 0 34224 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_369
timestamp 1649977179
transform 1 0 35052 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_377
timestamp 1649977179
transform 1 0 35788 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_385
timestamp 1649977179
transform 1 0 36524 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_393
timestamp 1649977179
transform 1 0 37260 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_405
timestamp 1649977179
transform 1 0 38364 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_412
timestamp 1649977179
transform 1 0 39008 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_423
timestamp 1649977179
transform 1 0 40020 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_429
timestamp 1649977179
transform 1 0 40572 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_441
timestamp 1649977179
transform 1 0 41676 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_453
timestamp 1649977179
transform 1 0 42780 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_465
timestamp 1649977179
transform 1 0 43884 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_473
timestamp 1649977179
transform 1 0 44620 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1649977179
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1649977179
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1649977179
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1649977179
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1649977179
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1649977179
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1649977179
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1649977179
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1649977179
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_569
timestamp 1649977179
transform 1 0 53452 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_575
timestamp 1649977179
transform 1 0 54004 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1649977179
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1649977179
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1649977179
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1649977179
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1649977179
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1649977179
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1649977179
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1649977179
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1649977179
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1649977179
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1649977179
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1649977179
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1649977179
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1649977179
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1649977179
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1649977179
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1649977179
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_169
timestamp 1649977179
transform 1 0 16652 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_181
timestamp 1649977179
transform 1 0 17756 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_191
timestamp 1649977179
transform 1 0 18676 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_197
timestamp 1649977179
transform 1 0 19228 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_203
timestamp 1649977179
transform 1 0 19780 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_209
timestamp 1649977179
transform 1 0 20332 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1649977179
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1649977179
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_225
timestamp 1649977179
transform 1 0 21804 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_228
timestamp 1649977179
transform 1 0 22080 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_234
timestamp 1649977179
transform 1 0 22632 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_241
timestamp 1649977179
transform 1 0 23276 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_248
timestamp 1649977179
transform 1 0 23920 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_259
timestamp 1649977179
transform 1 0 24932 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_263
timestamp 1649977179
transform 1 0 25300 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_270
timestamp 1649977179
transform 1 0 25944 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1649977179
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_285
timestamp 1649977179
transform 1 0 27324 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_295
timestamp 1649977179
transform 1 0 28244 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_319
timestamp 1649977179
transform 1 0 30452 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_326
timestamp 1649977179
transform 1 0 31096 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_332
timestamp 1649977179
transform 1 0 31648 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_339
timestamp 1649977179
transform 1 0 32292 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_345
timestamp 1649977179
transform 1 0 32844 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_349
timestamp 1649977179
transform 1 0 33212 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_355
timestamp 1649977179
transform 1 0 33764 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_364
timestamp 1649977179
transform 1 0 34592 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_373
timestamp 1649977179
transform 1 0 35420 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_388
timestamp 1649977179
transform 1 0 36800 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_393
timestamp 1649977179
transform 1 0 37260 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_410
timestamp 1649977179
transform 1 0 38824 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_420
timestamp 1649977179
transform 1 0 39744 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_432
timestamp 1649977179
transform 1 0 40848 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_444
timestamp 1649977179
transform 1 0 41952 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1649977179
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1649977179
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1649977179
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1649977179
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1649977179
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1649977179
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1649977179
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1649977179
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1649977179
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1649977179
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1649977179
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1649977179
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1649977179
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_573
timestamp 1649977179
transform 1 0 53820 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1649977179
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1649977179
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1649977179
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1649977179
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1649977179
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1649977179
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1649977179
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1649977179
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1649977179
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1649977179
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1649977179
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1649977179
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1649977179
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1649977179
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_153
timestamp 1649977179
transform 1 0 15180 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_161
timestamp 1649977179
transform 1 0 15916 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_164
timestamp 1649977179
transform 1 0 16192 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_170
timestamp 1649977179
transform 1 0 16744 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_183
timestamp 1649977179
transform 1 0 17940 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_187
timestamp 1649977179
transform 1 0 18308 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_192
timestamp 1649977179
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_202
timestamp 1649977179
transform 1 0 19688 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_209
timestamp 1649977179
transform 1 0 20332 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_213
timestamp 1649977179
transform 1 0 20700 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_217
timestamp 1649977179
transform 1 0 21068 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_223
timestamp 1649977179
transform 1 0 21620 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_226
timestamp 1649977179
transform 1 0 21896 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_232
timestamp 1649977179
transform 1 0 22448 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_239
timestamp 1649977179
transform 1 0 23092 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_248
timestamp 1649977179
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_261
timestamp 1649977179
transform 1 0 25116 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_269
timestamp 1649977179
transform 1 0 25852 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_277
timestamp 1649977179
transform 1 0 26588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_283
timestamp 1649977179
transform 1 0 27140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_289
timestamp 1649977179
transform 1 0 27692 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_295
timestamp 1649977179
transform 1 0 28244 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_299
timestamp 1649977179
transform 1 0 28612 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1649977179
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_317
timestamp 1649977179
transform 1 0 30268 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_329
timestamp 1649977179
transform 1 0 31372 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_335
timestamp 1649977179
transform 1 0 31924 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_341
timestamp 1649977179
transform 1 0 32476 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_347
timestamp 1649977179
transform 1 0 33028 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_353
timestamp 1649977179
transform 1 0 33580 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_360
timestamp 1649977179
transform 1 0 34224 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_368
timestamp 1649977179
transform 1 0 34960 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_374
timestamp 1649977179
transform 1 0 35512 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_382
timestamp 1649977179
transform 1 0 36248 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_386
timestamp 1649977179
transform 1 0 36616 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_398
timestamp 1649977179
transform 1 0 37720 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_408
timestamp 1649977179
transform 1 0 38640 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_414
timestamp 1649977179
transform 1 0 39192 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1649977179
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1649977179
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1649977179
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1649977179
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1649977179
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1649977179
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1649977179
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1649977179
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1649977179
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1649977179
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1649977179
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1649977179
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1649977179
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1649977179
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_557
timestamp 1649977179
transform 1 0 52348 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_561
timestamp 1649977179
transform 1 0 52716 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_564
timestamp 1649977179
transform 1 0 52992 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_572
timestamp 1649977179
transform 1 0 53728 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1649977179
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1649977179
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1649977179
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1649977179
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1649977179
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1649977179
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1649977179
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1649977179
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1649977179
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1649977179
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1649977179
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1649977179
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1649977179
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1649977179
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1649977179
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_149
timestamp 1649977179
transform 1 0 14812 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_155
timestamp 1649977179
transform 1 0 15364 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_158
timestamp 1649977179
transform 1 0 15640 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_164
timestamp 1649977179
transform 1 0 16192 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_169
timestamp 1649977179
transform 1 0 16652 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_173
timestamp 1649977179
transform 1 0 17020 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_183
timestamp 1649977179
transform 1 0 17940 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_187
timestamp 1649977179
transform 1 0 18308 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_193
timestamp 1649977179
transform 1 0 18860 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_201
timestamp 1649977179
transform 1 0 19596 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_208
timestamp 1649977179
transform 1 0 20240 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_220
timestamp 1649977179
transform 1 0 21344 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_229
timestamp 1649977179
transform 1 0 22172 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_235
timestamp 1649977179
transform 1 0 22724 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_238
timestamp 1649977179
transform 1 0 23000 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_245
timestamp 1649977179
transform 1 0 23644 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_255
timestamp 1649977179
transform 1 0 24564 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_266
timestamp 1649977179
transform 1 0 25576 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_276
timestamp 1649977179
transform 1 0 26496 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_298
timestamp 1649977179
transform 1 0 28520 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_304
timestamp 1649977179
transform 1 0 29072 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_325
timestamp 1649977179
transform 1 0 31004 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_331
timestamp 1649977179
transform 1 0 31556 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1649977179
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_343
timestamp 1649977179
transform 1 0 32660 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_351
timestamp 1649977179
transform 1 0 33396 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_360
timestamp 1649977179
transform 1 0 34224 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_366
timestamp 1649977179
transform 1 0 34776 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_375
timestamp 1649977179
transform 1 0 35604 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_379
timestamp 1649977179
transform 1 0 35972 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_383
timestamp 1649977179
transform 1 0 36340 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1649977179
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_393
timestamp 1649977179
transform 1 0 37260 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_401
timestamp 1649977179
transform 1 0 37996 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_407
timestamp 1649977179
transform 1 0 38548 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_413
timestamp 1649977179
transform 1 0 39100 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_425
timestamp 1649977179
transform 1 0 40204 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_437
timestamp 1649977179
transform 1 0 41308 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_445
timestamp 1649977179
transform 1 0 42044 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1649977179
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1649977179
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1649977179
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1649977179
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1649977179
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1649977179
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1649977179
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1649977179
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1649977179
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1649977179
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1649977179
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1649977179
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1649977179
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_573
timestamp 1649977179
transform 1 0 53820 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_3
timestamp 1649977179
transform 1 0 1380 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_7
timestamp 1649977179
transform 1 0 1748 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_19
timestamp 1649977179
transform 1 0 2852 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1649977179
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1649977179
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1649977179
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1649977179
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1649977179
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1649977179
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1649977179
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1649977179
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1649977179
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1649977179
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1649977179
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1649977179
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1649977179
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1649977179
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_155
timestamp 1649977179
transform 1 0 15364 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_161
timestamp 1649977179
transform 1 0 15916 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_170
timestamp 1649977179
transform 1 0 16744 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_174
timestamp 1649977179
transform 1 0 17112 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_181
timestamp 1649977179
transform 1 0 17756 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_188
timestamp 1649977179
transform 1 0 18400 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_200
timestamp 1649977179
transform 1 0 19504 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_204
timestamp 1649977179
transform 1 0 19872 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_211
timestamp 1649977179
transform 1 0 20516 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_221
timestamp 1649977179
transform 1 0 21436 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_230
timestamp 1649977179
transform 1 0 22264 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_239
timestamp 1649977179
transform 1 0 23092 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_245
timestamp 1649977179
transform 1 0 23644 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_248
timestamp 1649977179
transform 1 0 23920 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_258
timestamp 1649977179
transform 1 0 24840 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_265
timestamp 1649977179
transform 1 0 25484 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_274
timestamp 1649977179
transform 1 0 26312 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_282
timestamp 1649977179
transform 1 0 27048 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_288
timestamp 1649977179
transform 1 0 27600 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_294
timestamp 1649977179
transform 1 0 28152 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_304
timestamp 1649977179
transform 1 0 29072 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_309
timestamp 1649977179
transform 1 0 29532 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_317
timestamp 1649977179
transform 1 0 30268 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_329
timestamp 1649977179
transform 1 0 31372 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_338
timestamp 1649977179
transform 1 0 32200 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_66_355
timestamp 1649977179
transform 1 0 33764 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1649977179
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_365
timestamp 1649977179
transform 1 0 34684 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_371
timestamp 1649977179
transform 1 0 35236 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_379
timestamp 1649977179
transform 1 0 35972 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_386
timestamp 1649977179
transform 1 0 36616 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_396
timestamp 1649977179
transform 1 0 37536 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_402
timestamp 1649977179
transform 1 0 38088 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_408
timestamp 1649977179
transform 1 0 38640 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_414
timestamp 1649977179
transform 1 0 39192 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_423
timestamp 1649977179
transform 1 0 40020 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_435
timestamp 1649977179
transform 1 0 41124 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_447
timestamp 1649977179
transform 1 0 42228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_459
timestamp 1649977179
transform 1 0 43332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_471
timestamp 1649977179
transform 1 0 44436 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1649977179
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1649977179
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1649977179
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1649977179
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1649977179
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1649977179
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1649977179
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1649977179
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1649977179
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1649977179
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_569
timestamp 1649977179
transform 1 0 53452 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_575
timestamp 1649977179
transform 1 0 54004 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_3
timestamp 1649977179
transform 1 0 1380 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_11
timestamp 1649977179
transform 1 0 2116 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_23
timestamp 1649977179
transform 1 0 3220 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_35
timestamp 1649977179
transform 1 0 4324 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_47
timestamp 1649977179
transform 1 0 5428 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1649977179
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1649977179
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1649977179
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1649977179
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1649977179
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1649977179
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1649977179
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1649977179
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1649977179
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1649977179
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1649977179
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_164
timestamp 1649977179
transform 1 0 16192 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_174
timestamp 1649977179
transform 1 0 17112 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_184
timestamp 1649977179
transform 1 0 18032 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_192
timestamp 1649977179
transform 1 0 18768 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_196
timestamp 1649977179
transform 1 0 19136 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_199
timestamp 1649977179
transform 1 0 19412 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_208
timestamp 1649977179
transform 1 0 20240 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_220
timestamp 1649977179
transform 1 0 21344 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_232
timestamp 1649977179
transform 1 0 22448 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_238
timestamp 1649977179
transform 1 0 23000 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_242
timestamp 1649977179
transform 1 0 23368 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_252
timestamp 1649977179
transform 1 0 24288 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_258
timestamp 1649977179
transform 1 0 24840 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_264
timestamp 1649977179
transform 1 0 25392 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_270
timestamp 1649977179
transform 1 0 25944 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_276
timestamp 1649977179
transform 1 0 26496 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_287
timestamp 1649977179
transform 1 0 27508 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_293
timestamp 1649977179
transform 1 0 28060 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_301
timestamp 1649977179
transform 1 0 28796 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_304
timestamp 1649977179
transform 1 0 29072 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_314
timestamp 1649977179
transform 1 0 29992 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_326
timestamp 1649977179
transform 1 0 31096 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_332
timestamp 1649977179
transform 1 0 31648 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_354
timestamp 1649977179
transform 1 0 33672 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_363
timestamp 1649977179
transform 1 0 34500 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_374
timestamp 1649977179
transform 1 0 35512 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_380
timestamp 1649977179
transform 1 0 36064 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_388
timestamp 1649977179
transform 1 0 36800 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_398
timestamp 1649977179
transform 1 0 37720 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_413
timestamp 1649977179
transform 1 0 39100 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_419
timestamp 1649977179
transform 1 0 39652 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_425
timestamp 1649977179
transform 1 0 40204 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_431
timestamp 1649977179
transform 1 0 40756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_443
timestamp 1649977179
transform 1 0 41860 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1649977179
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1649977179
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1649977179
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1649977179
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1649977179
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1649977179
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1649977179
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1649977179
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1649977179
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1649977179
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1649977179
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1649977179
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1649977179
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1649977179
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_573
timestamp 1649977179
transform 1 0 53820 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1649977179
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1649977179
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1649977179
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1649977179
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1649977179
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1649977179
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1649977179
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1649977179
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1649977179
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1649977179
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1649977179
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1649977179
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1649977179
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1649977179
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1649977179
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_141
timestamp 1649977179
transform 1 0 14076 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_151
timestamp 1649977179
transform 1 0 14996 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_157
timestamp 1649977179
transform 1 0 15548 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_164
timestamp 1649977179
transform 1 0 16192 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_174
timestamp 1649977179
transform 1 0 17112 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_186
timestamp 1649977179
transform 1 0 18216 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_192
timestamp 1649977179
transform 1 0 18768 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_197
timestamp 1649977179
transform 1 0 19228 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_201
timestamp 1649977179
transform 1 0 19596 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_206
timestamp 1649977179
transform 1 0 20056 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_213
timestamp 1649977179
transform 1 0 20700 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_221
timestamp 1649977179
transform 1 0 21436 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_227
timestamp 1649977179
transform 1 0 21988 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_236
timestamp 1649977179
transform 1 0 22816 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_248
timestamp 1649977179
transform 1 0 23920 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_262
timestamp 1649977179
transform 1 0 25208 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_266
timestamp 1649977179
transform 1 0 25576 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_269
timestamp 1649977179
transform 1 0 25852 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_277
timestamp 1649977179
transform 1 0 26588 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_300
timestamp 1649977179
transform 1 0 28704 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_309
timestamp 1649977179
transform 1 0 29532 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_313
timestamp 1649977179
transform 1 0 29900 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_325
timestamp 1649977179
transform 1 0 31004 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_334
timestamp 1649977179
transform 1 0 31832 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_344
timestamp 1649977179
transform 1 0 32752 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_353
timestamp 1649977179
transform 1 0 33580 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_359
timestamp 1649977179
transform 1 0 34132 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1649977179
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_369
timestamp 1649977179
transform 1 0 35052 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_376
timestamp 1649977179
transform 1 0 35696 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_380
timestamp 1649977179
transform 1 0 36064 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_386
timestamp 1649977179
transform 1 0 36616 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_392
timestamp 1649977179
transform 1 0 37168 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_399
timestamp 1649977179
transform 1 0 37812 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_416
timestamp 1649977179
transform 1 0 39376 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_423
timestamp 1649977179
transform 1 0 40020 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_429
timestamp 1649977179
transform 1 0 40572 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_435
timestamp 1649977179
transform 1 0 41124 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_441
timestamp 1649977179
transform 1 0 41676 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_453
timestamp 1649977179
transform 1 0 42780 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_465
timestamp 1649977179
transform 1 0 43884 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_473
timestamp 1649977179
transform 1 0 44620 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1649977179
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1649977179
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1649977179
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1649977179
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1649977179
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1649977179
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1649977179
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1649977179
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1649977179
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_569
timestamp 1649977179
transform 1 0 53452 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_575
timestamp 1649977179
transform 1 0 54004 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1649977179
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1649977179
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1649977179
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1649977179
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1649977179
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1649977179
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1649977179
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1649977179
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1649977179
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1649977179
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1649977179
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1649977179
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1649977179
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1649977179
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1649977179
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1649977179
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_161
timestamp 1649977179
transform 1 0 15916 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_164
timestamp 1649977179
transform 1 0 16192 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_169
timestamp 1649977179
transform 1 0 16652 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_178
timestamp 1649977179
transform 1 0 17480 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_188
timestamp 1649977179
transform 1 0 18400 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_197
timestamp 1649977179
transform 1 0 19228 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_204
timestamp 1649977179
transform 1 0 19872 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_69_214
timestamp 1649977179
transform 1 0 20792 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_220
timestamp 1649977179
transform 1 0 21344 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_225
timestamp 1649977179
transform 1 0 21804 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_232
timestamp 1649977179
transform 1 0 22448 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_242
timestamp 1649977179
transform 1 0 23368 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_252
timestamp 1649977179
transform 1 0 24288 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_261
timestamp 1649977179
transform 1 0 25116 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_269
timestamp 1649977179
transform 1 0 25852 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_273
timestamp 1649977179
transform 1 0 26220 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_276
timestamp 1649977179
transform 1 0 26496 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_281
timestamp 1649977179
transform 1 0 26956 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_286
timestamp 1649977179
transform 1 0 27416 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_306
timestamp 1649977179
transform 1 0 29256 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_312
timestamp 1649977179
transform 1 0 29808 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_320
timestamp 1649977179
transform 1 0 30544 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_327
timestamp 1649977179
transform 1 0 31188 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1649977179
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_339
timestamp 1649977179
transform 1 0 32292 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_69_351
timestamp 1649977179
transform 1 0 33396 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_359
timestamp 1649977179
transform 1 0 34132 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_365
timestamp 1649977179
transform 1 0 34684 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_373
timestamp 1649977179
transform 1 0 35420 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_377
timestamp 1649977179
transform 1 0 35788 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_384
timestamp 1649977179
transform 1 0 36432 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_393
timestamp 1649977179
transform 1 0 37260 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_398
timestamp 1649977179
transform 1 0 37720 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_412
timestamp 1649977179
transform 1 0 39008 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_424
timestamp 1649977179
transform 1 0 40112 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_430
timestamp 1649977179
transform 1 0 40664 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_436
timestamp 1649977179
transform 1 0 41216 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_442
timestamp 1649977179
transform 1 0 41768 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1649977179
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1649977179
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1649977179
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1649977179
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1649977179
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1649977179
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1649977179
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1649977179
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1649977179
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1649977179
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1649977179
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1649977179
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_561
timestamp 1649977179
transform 1 0 52716 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_564
timestamp 1649977179
transform 1 0 52992 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_572
timestamp 1649977179
transform 1 0 53728 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1649977179
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1649977179
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1649977179
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1649977179
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1649977179
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1649977179
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1649977179
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1649977179
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1649977179
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1649977179
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1649977179
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1649977179
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1649977179
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1649977179
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1649977179
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1649977179
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_153
timestamp 1649977179
transform 1 0 15180 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_158
timestamp 1649977179
transform 1 0 15640 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_164
timestamp 1649977179
transform 1 0 16192 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_170
timestamp 1649977179
transform 1 0 16744 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_176
timestamp 1649977179
transform 1 0 17296 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_184
timestamp 1649977179
transform 1 0 18032 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_191
timestamp 1649977179
transform 1 0 18676 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1649977179
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_197
timestamp 1649977179
transform 1 0 19228 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_201
timestamp 1649977179
transform 1 0 19596 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_207
timestamp 1649977179
transform 1 0 20148 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_216
timestamp 1649977179
transform 1 0 20976 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_226
timestamp 1649977179
transform 1 0 21896 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_232
timestamp 1649977179
transform 1 0 22448 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_239
timestamp 1649977179
transform 1 0 23092 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_248
timestamp 1649977179
transform 1 0 23920 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_260
timestamp 1649977179
transform 1 0 25024 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_266
timestamp 1649977179
transform 1 0 25576 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_269
timestamp 1649977179
transform 1 0 25852 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_282
timestamp 1649977179
transform 1 0 27048 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_70_304
timestamp 1649977179
transform 1 0 29072 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_316
timestamp 1649977179
transform 1 0 30176 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_325
timestamp 1649977179
transform 1 0 31004 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_334
timestamp 1649977179
transform 1 0 31832 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_341
timestamp 1649977179
transform 1 0 32476 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_347
timestamp 1649977179
transform 1 0 33028 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_355
timestamp 1649977179
transform 1 0 33764 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1649977179
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_368
timestamp 1649977179
transform 1 0 34960 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_375
timestamp 1649977179
transform 1 0 35604 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_379
timestamp 1649977179
transform 1 0 35972 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_397
timestamp 1649977179
transform 1 0 37628 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_70_416
timestamp 1649977179
transform 1 0 39376 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_424
timestamp 1649977179
transform 1 0 40112 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_430
timestamp 1649977179
transform 1 0 40664 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_436
timestamp 1649977179
transform 1 0 41216 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_442
timestamp 1649977179
transform 1 0 41768 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_454
timestamp 1649977179
transform 1 0 42872 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_466
timestamp 1649977179
transform 1 0 43976 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_474
timestamp 1649977179
transform 1 0 44712 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1649977179
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1649977179
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1649977179
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1649977179
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1649977179
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1649977179
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1649977179
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1649977179
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1649977179
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_569
timestamp 1649977179
transform 1 0 53452 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_575
timestamp 1649977179
transform 1 0 54004 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_7
timestamp 1649977179
transform 1 0 1748 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_13
timestamp 1649977179
transform 1 0 2300 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_25
timestamp 1649977179
transform 1 0 3404 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_37
timestamp 1649977179
transform 1 0 4508 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_49
timestamp 1649977179
transform 1 0 5612 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1649977179
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1649977179
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1649977179
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1649977179
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1649977179
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1649977179
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1649977179
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1649977179
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1649977179
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1649977179
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1649977179
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_161
timestamp 1649977179
transform 1 0 15916 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_164
timestamp 1649977179
transform 1 0 16192 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_71_169
timestamp 1649977179
transform 1 0 16652 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_174
timestamp 1649977179
transform 1 0 17112 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_184
timestamp 1649977179
transform 1 0 18032 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_193
timestamp 1649977179
transform 1 0 18860 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_214
timestamp 1649977179
transform 1 0 20792 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_220
timestamp 1649977179
transform 1 0 21344 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_225
timestamp 1649977179
transform 1 0 21804 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_229
timestamp 1649977179
transform 1 0 22172 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_235
timestamp 1649977179
transform 1 0 22724 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_241
timestamp 1649977179
transform 1 0 23276 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_248
timestamp 1649977179
transform 1 0 23920 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_256
timestamp 1649977179
transform 1 0 24656 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_263
timestamp 1649977179
transform 1 0 25300 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_267
timestamp 1649977179
transform 1 0 25668 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_270
timestamp 1649977179
transform 1 0 25944 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_276
timestamp 1649977179
transform 1 0 26496 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_300
timestamp 1649977179
transform 1 0 28704 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_308
timestamp 1649977179
transform 1 0 29440 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_318
timestamp 1649977179
transform 1 0 30360 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1649977179
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1649977179
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_337
timestamp 1649977179
transform 1 0 32108 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_343
timestamp 1649977179
transform 1 0 32660 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_347
timestamp 1649977179
transform 1 0 33028 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_356
timestamp 1649977179
transform 1 0 33856 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_365
timestamp 1649977179
transform 1 0 34684 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_378
timestamp 1649977179
transform 1 0 35880 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_388
timestamp 1649977179
transform 1 0 36800 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_393
timestamp 1649977179
transform 1 0 37260 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_397
timestamp 1649977179
transform 1 0 37628 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_406
timestamp 1649977179
transform 1 0 38456 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_417
timestamp 1649977179
transform 1 0 39468 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_423
timestamp 1649977179
transform 1 0 40020 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_429
timestamp 1649977179
transform 1 0 40572 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_435
timestamp 1649977179
transform 1 0 41124 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1649977179
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1649977179
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_451
timestamp 1649977179
transform 1 0 42596 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_463
timestamp 1649977179
transform 1 0 43700 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_475
timestamp 1649977179
transform 1 0 44804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_487
timestamp 1649977179
transform 1 0 45908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_499
timestamp 1649977179
transform 1 0 47012 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1649977179
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1649977179
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1649977179
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1649977179
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1649977179
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1649977179
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1649977179
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1649977179
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_573
timestamp 1649977179
transform 1 0 53820 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1649977179
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1649977179
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1649977179
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1649977179
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1649977179
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1649977179
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1649977179
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1649977179
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1649977179
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1649977179
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1649977179
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1649977179
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1649977179
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1649977179
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1649977179
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_72_141
timestamp 1649977179
transform 1 0 14076 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_72_146
timestamp 1649977179
transform 1 0 14536 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_154
timestamp 1649977179
transform 1 0 15272 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_157
timestamp 1649977179
transform 1 0 15548 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_163
timestamp 1649977179
transform 1 0 16100 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_169
timestamp 1649977179
transform 1 0 16652 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_175
timestamp 1649977179
transform 1 0 17204 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_185
timestamp 1649977179
transform 1 0 18124 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_189
timestamp 1649977179
transform 1 0 18492 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_192
timestamp 1649977179
transform 1 0 18768 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_197
timestamp 1649977179
transform 1 0 19228 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_203
timestamp 1649977179
transform 1 0 19780 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_219
timestamp 1649977179
transform 1 0 21252 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_230
timestamp 1649977179
transform 1 0 22264 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_238
timestamp 1649977179
transform 1 0 23000 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_244
timestamp 1649977179
transform 1 0 23552 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_253
timestamp 1649977179
transform 1 0 24380 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_261
timestamp 1649977179
transform 1 0 25116 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_270
timestamp 1649977179
transform 1 0 25944 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_278
timestamp 1649977179
transform 1 0 26680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_286
timestamp 1649977179
transform 1 0 27416 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_293
timestamp 1649977179
transform 1 0 28060 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_301
timestamp 1649977179
transform 1 0 28796 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_304
timestamp 1649977179
transform 1 0 29072 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_309
timestamp 1649977179
transform 1 0 29532 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_333
timestamp 1649977179
transform 1 0 31740 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_354
timestamp 1649977179
transform 1 0 33672 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_360
timestamp 1649977179
transform 1 0 34224 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_370
timestamp 1649977179
transform 1 0 35144 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_376
timestamp 1649977179
transform 1 0 35696 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_387
timestamp 1649977179
transform 1 0 36708 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_398
timestamp 1649977179
transform 1 0 37720 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_407
timestamp 1649977179
transform 1 0 38548 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_414
timestamp 1649977179
transform 1 0 39192 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_423
timestamp 1649977179
transform 1 0 40020 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_429
timestamp 1649977179
transform 1 0 40572 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_435
timestamp 1649977179
transform 1 0 41124 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_441
timestamp 1649977179
transform 1 0 41676 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_447
timestamp 1649977179
transform 1 0 42228 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_453
timestamp 1649977179
transform 1 0 42780 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_465
timestamp 1649977179
transform 1 0 43884 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_473
timestamp 1649977179
transform 1 0 44620 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1649977179
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1649977179
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1649977179
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1649977179
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1649977179
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1649977179
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1649977179
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1649977179
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_557
timestamp 1649977179
transform 1 0 52348 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_561
timestamp 1649977179
transform 1 0 52716 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_564
timestamp 1649977179
transform 1 0 52992 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_572
timestamp 1649977179
transform 1 0 53728 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1649977179
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1649977179
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1649977179
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1649977179
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1649977179
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1649977179
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1649977179
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1649977179
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1649977179
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1649977179
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1649977179
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1649977179
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1649977179
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_125
timestamp 1649977179
transform 1 0 12604 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_133
timestamp 1649977179
transform 1 0 13340 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_138
timestamp 1649977179
transform 1 0 13800 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_144
timestamp 1649977179
transform 1 0 14352 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_151
timestamp 1649977179
transform 1 0 14996 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_159
timestamp 1649977179
transform 1 0 15732 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_164
timestamp 1649977179
transform 1 0 16192 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_174
timestamp 1649977179
transform 1 0 17112 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_181
timestamp 1649977179
transform 1 0 17756 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_189
timestamp 1649977179
transform 1 0 18492 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_195
timestamp 1649977179
transform 1 0 19044 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_204
timestamp 1649977179
transform 1 0 19872 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_216
timestamp 1649977179
transform 1 0 20976 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_73_232
timestamp 1649977179
transform 1 0 22448 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_243
timestamp 1649977179
transform 1 0 23460 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_249
timestamp 1649977179
transform 1 0 24012 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_256
timestamp 1649977179
transform 1 0 24656 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_264
timestamp 1649977179
transform 1 0 25392 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_270
timestamp 1649977179
transform 1 0 25944 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_276
timestamp 1649977179
transform 1 0 26496 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_281
timestamp 1649977179
transform 1 0 26956 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_286
timestamp 1649977179
transform 1 0 27416 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_295
timestamp 1649977179
transform 1 0 28244 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_303
timestamp 1649977179
transform 1 0 28980 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_307
timestamp 1649977179
transform 1 0 29348 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_325
timestamp 1649977179
transform 1 0 31004 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_331
timestamp 1649977179
transform 1 0 31556 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1649977179
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_340
timestamp 1649977179
transform 1 0 32384 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_353
timestamp 1649977179
transform 1 0 33580 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_364
timestamp 1649977179
transform 1 0 34592 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_373
timestamp 1649977179
transform 1 0 35420 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_377
timestamp 1649977179
transform 1 0 35788 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1649977179
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1649977179
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_399
timestamp 1649977179
transform 1 0 37812 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_406
timestamp 1649977179
transform 1 0 38456 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_412
timestamp 1649977179
transform 1 0 39008 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_418
timestamp 1649977179
transform 1 0 39560 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_424
timestamp 1649977179
transform 1 0 40112 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_430
timestamp 1649977179
transform 1 0 40664 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_436
timestamp 1649977179
transform 1 0 41216 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_442
timestamp 1649977179
transform 1 0 41768 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1649977179
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1649977179
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1649977179
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1649977179
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1649977179
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1649977179
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1649977179
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1649977179
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1649977179
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1649977179
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1649977179
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1649977179
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1649977179
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_573
timestamp 1649977179
transform 1 0 53820 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1649977179
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1649977179
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1649977179
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1649977179
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1649977179
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1649977179
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1649977179
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1649977179
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1649977179
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1649977179
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1649977179
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1649977179
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_121
timestamp 1649977179
transform 1 0 12236 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_127
timestamp 1649977179
transform 1 0 12788 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_130
timestamp 1649977179
transform 1 0 13064 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_136
timestamp 1649977179
transform 1 0 13616 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_144
timestamp 1649977179
transform 1 0 14352 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_153
timestamp 1649977179
transform 1 0 15180 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_165
timestamp 1649977179
transform 1 0 16284 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_176
timestamp 1649977179
transform 1 0 17296 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_185
timestamp 1649977179
transform 1 0 18124 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_189
timestamp 1649977179
transform 1 0 18492 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_192
timestamp 1649977179
transform 1 0 18768 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_197
timestamp 1649977179
transform 1 0 19228 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_200
timestamp 1649977179
transform 1 0 19504 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_210
timestamp 1649977179
transform 1 0 20424 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_221
timestamp 1649977179
transform 1 0 21436 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_227
timestamp 1649977179
transform 1 0 21988 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_233
timestamp 1649977179
transform 1 0 22540 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_240
timestamp 1649977179
transform 1 0 23184 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_248
timestamp 1649977179
transform 1 0 23920 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_258
timestamp 1649977179
transform 1 0 24840 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_265
timestamp 1649977179
transform 1 0 25484 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_271
timestamp 1649977179
transform 1 0 26036 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_274
timestamp 1649977179
transform 1 0 26312 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_280
timestamp 1649977179
transform 1 0 26864 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_291
timestamp 1649977179
transform 1 0 27876 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_304
timestamp 1649977179
transform 1 0 29072 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_316
timestamp 1649977179
transform 1 0 30176 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_322
timestamp 1649977179
transform 1 0 30728 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_328
timestamp 1649977179
transform 1 0 31280 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_74_339
timestamp 1649977179
transform 1 0 32292 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_348
timestamp 1649977179
transform 1 0 33120 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_354
timestamp 1649977179
transform 1 0 33672 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_359
timestamp 1649977179
transform 1 0 34132 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1649977179
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_368
timestamp 1649977179
transform 1 0 34960 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_375
timestamp 1649977179
transform 1 0 35604 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_384
timestamp 1649977179
transform 1 0 36432 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_393
timestamp 1649977179
transform 1 0 37260 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_400
timestamp 1649977179
transform 1 0 37904 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_406
timestamp 1649977179
transform 1 0 38456 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_412
timestamp 1649977179
transform 1 0 39008 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_74_423
timestamp 1649977179
transform 1 0 40020 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_429
timestamp 1649977179
transform 1 0 40572 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_435
timestamp 1649977179
transform 1 0 41124 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_447
timestamp 1649977179
transform 1 0 42228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_459
timestamp 1649977179
transform 1 0 43332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_471
timestamp 1649977179
transform 1 0 44436 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1649977179
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1649977179
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1649977179
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1649977179
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1649977179
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1649977179
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1649977179
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1649977179
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1649977179
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1649977179
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_569
timestamp 1649977179
transform 1 0 53452 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_575
timestamp 1649977179
transform 1 0 54004 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_3
timestamp 1649977179
transform 1 0 1380 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_7
timestamp 1649977179
transform 1 0 1748 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_19
timestamp 1649977179
transform 1 0 2852 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_31
timestamp 1649977179
transform 1 0 3956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_43
timestamp 1649977179
transform 1 0 5060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1649977179
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1649977179
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1649977179
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1649977179
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1649977179
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1649977179
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1649977179
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1649977179
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_125
timestamp 1649977179
transform 1 0 12604 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_131
timestamp 1649977179
transform 1 0 13156 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_137
timestamp 1649977179
transform 1 0 13708 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_146
timestamp 1649977179
transform 1 0 14536 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_158
timestamp 1649977179
transform 1 0 15640 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_164
timestamp 1649977179
transform 1 0 16192 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_176
timestamp 1649977179
transform 1 0 17296 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_185
timestamp 1649977179
transform 1 0 18124 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_193
timestamp 1649977179
transform 1 0 18860 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_75_205
timestamp 1649977179
transform 1 0 19964 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_213
timestamp 1649977179
transform 1 0 20700 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_220
timestamp 1649977179
transform 1 0 21344 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_225
timestamp 1649977179
transform 1 0 21804 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_229
timestamp 1649977179
transform 1 0 22172 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_238
timestamp 1649977179
transform 1 0 23000 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_250
timestamp 1649977179
transform 1 0 24104 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_260
timestamp 1649977179
transform 1 0 25024 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_269
timestamp 1649977179
transform 1 0 25852 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_273
timestamp 1649977179
transform 1 0 26220 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_276
timestamp 1649977179
transform 1 0 26496 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_281
timestamp 1649977179
transform 1 0 26956 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_290
timestamp 1649977179
transform 1 0 27784 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_298
timestamp 1649977179
transform 1 0 28520 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_319
timestamp 1649977179
transform 1 0 30452 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_330
timestamp 1649977179
transform 1 0 31464 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_337
timestamp 1649977179
transform 1 0 32108 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_348
timestamp 1649977179
transform 1 0 33120 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_356
timestamp 1649977179
transform 1 0 33856 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_363
timestamp 1649977179
transform 1 0 34500 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_369
timestamp 1649977179
transform 1 0 35052 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_373
timestamp 1649977179
transform 1 0 35420 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_377
timestamp 1649977179
transform 1 0 35788 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1649977179
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1649977179
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_395
timestamp 1649977179
transform 1 0 37444 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_401
timestamp 1649977179
transform 1 0 37996 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_407
timestamp 1649977179
transform 1 0 38548 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_413
timestamp 1649977179
transform 1 0 39100 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_419
timestamp 1649977179
transform 1 0 39652 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_425
timestamp 1649977179
transform 1 0 40204 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_437
timestamp 1649977179
transform 1 0 41308 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_445
timestamp 1649977179
transform 1 0 42044 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1649977179
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1649977179
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1649977179
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1649977179
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1649977179
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1649977179
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1649977179
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1649977179
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1649977179
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1649977179
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1649977179
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1649977179
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1649977179
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_573
timestamp 1649977179
transform 1 0 53820 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_3
timestamp 1649977179
transform 1 0 1380 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_11
timestamp 1649977179
transform 1 0 2116 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_23
timestamp 1649977179
transform 1 0 3220 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1649977179
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1649977179
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1649977179
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1649977179
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1649977179
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1649977179
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1649977179
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1649977179
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1649977179
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1649977179
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1649977179
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_133
timestamp 1649977179
transform 1 0 13340 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_136
timestamp 1649977179
transform 1 0 13616 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_141
timestamp 1649977179
transform 1 0 14076 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_144
timestamp 1649977179
transform 1 0 14352 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_151
timestamp 1649977179
transform 1 0 14996 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_159
timestamp 1649977179
transform 1 0 15732 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_168
timestamp 1649977179
transform 1 0 16560 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_179
timestamp 1649977179
transform 1 0 17572 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1649977179
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1649977179
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_76_197
timestamp 1649977179
transform 1 0 19228 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_76_204
timestamp 1649977179
transform 1 0 19872 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_214
timestamp 1649977179
transform 1 0 20792 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_222
timestamp 1649977179
transform 1 0 21528 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_229
timestamp 1649977179
transform 1 0 22172 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_238
timestamp 1649977179
transform 1 0 23000 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_248
timestamp 1649977179
transform 1 0 23920 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_255
timestamp 1649977179
transform 1 0 24564 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_259
timestamp 1649977179
transform 1 0 24932 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_266
timestamp 1649977179
transform 1 0 25576 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_277
timestamp 1649977179
transform 1 0 26588 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_300
timestamp 1649977179
transform 1 0 28704 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_326
timestamp 1649977179
transform 1 0 31096 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_347
timestamp 1649977179
transform 1 0 33028 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_356
timestamp 1649977179
transform 1 0 33856 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_367
timestamp 1649977179
transform 1 0 34868 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_373
timestamp 1649977179
transform 1 0 35420 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_384
timestamp 1649977179
transform 1 0 36432 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_390
timestamp 1649977179
transform 1 0 36984 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_396
timestamp 1649977179
transform 1 0 37536 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_402
timestamp 1649977179
transform 1 0 38088 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_408
timestamp 1649977179
transform 1 0 38640 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_414
timestamp 1649977179
transform 1 0 39192 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1649977179
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1649977179
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1649977179
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1649977179
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1649977179
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1649977179
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1649977179
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1649977179
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1649977179
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1649977179
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1649977179
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1649977179
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1649977179
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1649977179
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_557
timestamp 1649977179
transform 1 0 52348 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_561
timestamp 1649977179
transform 1 0 52716 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_564
timestamp 1649977179
transform 1 0 52992 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_572
timestamp 1649977179
transform 1 0 53728 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1649977179
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1649977179
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1649977179
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1649977179
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1649977179
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1649977179
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1649977179
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1649977179
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1649977179
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1649977179
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1649977179
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1649977179
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1649977179
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1649977179
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_139
timestamp 1649977179
transform 1 0 13892 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_77_147
timestamp 1649977179
transform 1 0 14628 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_153
timestamp 1649977179
transform 1 0 15180 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_160
timestamp 1649977179
transform 1 0 15824 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_77_172
timestamp 1649977179
transform 1 0 16928 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_181
timestamp 1649977179
transform 1 0 17756 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_187
timestamp 1649977179
transform 1 0 18308 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_192
timestamp 1649977179
transform 1 0 18768 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_201
timestamp 1649977179
transform 1 0 19596 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_205
timestamp 1649977179
transform 1 0 19964 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_211
timestamp 1649977179
transform 1 0 20516 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_220
timestamp 1649977179
transform 1 0 21344 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_230
timestamp 1649977179
transform 1 0 22264 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_237
timestamp 1649977179
transform 1 0 22908 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_246
timestamp 1649977179
transform 1 0 23736 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_257
timestamp 1649977179
transform 1 0 24748 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_267
timestamp 1649977179
transform 1 0 25668 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_276
timestamp 1649977179
transform 1 0 26496 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_281
timestamp 1649977179
transform 1 0 26956 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_285
timestamp 1649977179
transform 1 0 27324 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_293
timestamp 1649977179
transform 1 0 28060 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_77_319
timestamp 1649977179
transform 1 0 30452 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1649977179
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1649977179
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_340
timestamp 1649977179
transform 1 0 32384 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_353
timestamp 1649977179
transform 1 0 33580 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_77_363
timestamp 1649977179
transform 1 0 34500 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_371
timestamp 1649977179
transform 1 0 35236 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_377
timestamp 1649977179
transform 1 0 35788 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_386
timestamp 1649977179
transform 1 0 36616 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_77_395
timestamp 1649977179
transform 1 0 37444 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_401
timestamp 1649977179
transform 1 0 37996 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_407
timestamp 1649977179
transform 1 0 38548 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_413
timestamp 1649977179
transform 1 0 39100 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_425
timestamp 1649977179
transform 1 0 40204 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_437
timestamp 1649977179
transform 1 0 41308 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_445
timestamp 1649977179
transform 1 0 42044 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1649977179
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1649977179
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1649977179
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1649977179
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1649977179
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1649977179
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1649977179
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1649977179
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1649977179
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1649977179
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1649977179
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1649977179
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1649977179
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_573
timestamp 1649977179
transform 1 0 53820 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1649977179
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1649977179
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1649977179
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1649977179
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1649977179
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1649977179
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1649977179
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1649977179
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1649977179
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1649977179
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1649977179
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1649977179
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1649977179
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1649977179
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1649977179
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1649977179
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_153
timestamp 1649977179
transform 1 0 15180 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_156
timestamp 1649977179
transform 1 0 15456 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_162
timestamp 1649977179
transform 1 0 16008 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_168
timestamp 1649977179
transform 1 0 16560 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_176
timestamp 1649977179
transform 1 0 17296 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_183
timestamp 1649977179
transform 1 0 17940 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_189
timestamp 1649977179
transform 1 0 18492 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_192
timestamp 1649977179
transform 1 0 18768 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_199
timestamp 1649977179
transform 1 0 19412 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_208
timestamp 1649977179
transform 1 0 20240 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_219
timestamp 1649977179
transform 1 0 21252 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_226
timestamp 1649977179
transform 1 0 21896 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_230
timestamp 1649977179
transform 1 0 22264 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_236
timestamp 1649977179
transform 1 0 22816 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_240
timestamp 1649977179
transform 1 0 23184 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_248
timestamp 1649977179
transform 1 0 23920 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_260
timestamp 1649977179
transform 1 0 25024 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_268
timestamp 1649977179
transform 1 0 25760 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_274
timestamp 1649977179
transform 1 0 26312 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_277
timestamp 1649977179
transform 1 0 26588 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_285
timestamp 1649977179
transform 1 0 27324 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_293
timestamp 1649977179
transform 1 0 28060 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_296
timestamp 1649977179
transform 1 0 28336 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_304
timestamp 1649977179
transform 1 0 29072 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_328
timestamp 1649977179
transform 1 0 31280 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_337
timestamp 1649977179
transform 1 0 32108 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_341
timestamp 1649977179
transform 1 0 32476 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_345
timestamp 1649977179
transform 1 0 32844 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_355
timestamp 1649977179
transform 1 0 33764 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1649977179
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_372
timestamp 1649977179
transform 1 0 35328 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_382
timestamp 1649977179
transform 1 0 36248 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_389
timestamp 1649977179
transform 1 0 36892 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_395
timestamp 1649977179
transform 1 0 37444 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_401
timestamp 1649977179
transform 1 0 37996 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_407
timestamp 1649977179
transform 1 0 38548 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1649977179
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1649977179
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1649977179
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1649977179
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1649977179
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1649977179
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1649977179
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1649977179
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1649977179
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1649977179
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1649977179
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1649977179
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1649977179
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1649977179
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1649977179
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1649977179
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1649977179
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_569
timestamp 1649977179
transform 1 0 53452 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_575
timestamp 1649977179
transform 1 0 54004 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_3
timestamp 1649977179
transform 1 0 1380 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_7
timestamp 1649977179
transform 1 0 1748 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_19
timestamp 1649977179
transform 1 0 2852 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_31
timestamp 1649977179
transform 1 0 3956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_43
timestamp 1649977179
transform 1 0 5060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1649977179
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1649977179
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1649977179
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1649977179
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1649977179
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1649977179
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1649977179
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1649977179
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1649977179
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1649977179
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1649977179
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1649977179
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1649977179
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_169
timestamp 1649977179
transform 1 0 16652 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_173
timestamp 1649977179
transform 1 0 17020 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_176
timestamp 1649977179
transform 1 0 17296 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_182
timestamp 1649977179
transform 1 0 17848 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_188
timestamp 1649977179
transform 1 0 18400 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_194
timestamp 1649977179
transform 1 0 18952 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_201
timestamp 1649977179
transform 1 0 19596 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_209
timestamp 1649977179
transform 1 0 20332 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_216
timestamp 1649977179
transform 1 0 20976 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_227
timestamp 1649977179
transform 1 0 21988 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_233
timestamp 1649977179
transform 1 0 22540 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_240
timestamp 1649977179
transform 1 0 23184 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_248
timestamp 1649977179
transform 1 0 23920 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_258
timestamp 1649977179
transform 1 0 24840 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_264
timestamp 1649977179
transform 1 0 25392 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_270
timestamp 1649977179
transform 1 0 25944 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_276
timestamp 1649977179
transform 1 0 26496 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_79_281
timestamp 1649977179
transform 1 0 26956 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_288
timestamp 1649977179
transform 1 0 27600 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_294
timestamp 1649977179
transform 1 0 28152 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_300
timestamp 1649977179
transform 1 0 28704 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_306
timestamp 1649977179
transform 1 0 29256 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_312
timestamp 1649977179
transform 1 0 29808 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_318
timestamp 1649977179
transform 1 0 30360 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_326
timestamp 1649977179
transform 1 0 31096 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1649977179
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1649977179
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_79_337
timestamp 1649977179
transform 1 0 32108 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_342
timestamp 1649977179
transform 1 0 32568 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_350
timestamp 1649977179
transform 1 0 33304 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_356
timestamp 1649977179
transform 1 0 33856 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_360
timestamp 1649977179
transform 1 0 34224 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_369
timestamp 1649977179
transform 1 0 35052 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_378
timestamp 1649977179
transform 1 0 35880 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_384
timestamp 1649977179
transform 1 0 36432 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_395
timestamp 1649977179
transform 1 0 37444 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_401
timestamp 1649977179
transform 1 0 37996 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_413
timestamp 1649977179
transform 1 0 39100 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_425
timestamp 1649977179
transform 1 0 40204 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_437
timestamp 1649977179
transform 1 0 41308 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_445
timestamp 1649977179
transform 1 0 42044 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1649977179
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1649977179
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1649977179
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1649977179
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1649977179
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1649977179
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1649977179
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1649977179
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1649977179
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1649977179
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1649977179
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1649977179
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1649977179
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_573
timestamp 1649977179
transform 1 0 53820 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_3
timestamp 1649977179
transform 1 0 1380 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_11
timestamp 1649977179
transform 1 0 2116 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_23
timestamp 1649977179
transform 1 0 3220 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1649977179
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1649977179
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1649977179
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1649977179
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1649977179
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1649977179
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1649977179
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1649977179
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1649977179
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1649977179
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1649977179
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1649977179
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1649977179
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1649977179
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1649977179
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1649977179
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_177
timestamp 1649977179
transform 1 0 17388 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_180
timestamp 1649977179
transform 1 0 17664 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_188
timestamp 1649977179
transform 1 0 18400 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_192
timestamp 1649977179
transform 1 0 18768 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_197
timestamp 1649977179
transform 1 0 19228 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_203
timestamp 1649977179
transform 1 0 19780 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_210
timestamp 1649977179
transform 1 0 20424 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_218
timestamp 1649977179
transform 1 0 21160 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_224
timestamp 1649977179
transform 1 0 21712 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_230
timestamp 1649977179
transform 1 0 22264 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_236
timestamp 1649977179
transform 1 0 22816 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_242
timestamp 1649977179
transform 1 0 23368 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_248
timestamp 1649977179
transform 1 0 23920 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_255
timestamp 1649977179
transform 1 0 24564 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_261
timestamp 1649977179
transform 1 0 25116 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_268
timestamp 1649977179
transform 1 0 25760 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_293
timestamp 1649977179
transform 1 0 28060 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_299
timestamp 1649977179
transform 1 0 28612 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1649977179
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_313
timestamp 1649977179
transform 1 0 29900 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_319
timestamp 1649977179
transform 1 0 30452 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_325
timestamp 1649977179
transform 1 0 31004 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_331
timestamp 1649977179
transform 1 0 31556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_342
timestamp 1649977179
transform 1 0 32568 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_351
timestamp 1649977179
transform 1 0 33396 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_355
timestamp 1649977179
transform 1 0 33764 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_360
timestamp 1649977179
transform 1 0 34224 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_371
timestamp 1649977179
transform 1 0 35236 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_378
timestamp 1649977179
transform 1 0 35880 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_384
timestamp 1649977179
transform 1 0 36432 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_390
timestamp 1649977179
transform 1 0 36984 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_396
timestamp 1649977179
transform 1 0 37536 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_408
timestamp 1649977179
transform 1 0 38640 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1649977179
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1649977179
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1649977179
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1649977179
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1649977179
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1649977179
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1649977179
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1649977179
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1649977179
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1649977179
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1649977179
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1649977179
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1649977179
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1649977179
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1649977179
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_569
timestamp 1649977179
transform 1 0 53452 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_575
timestamp 1649977179
transform 1 0 54004 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1649977179
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1649977179
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1649977179
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1649977179
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1649977179
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1649977179
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1649977179
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1649977179
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1649977179
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1649977179
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1649977179
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1649977179
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1649977179
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1649977179
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1649977179
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1649977179
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1649977179
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1649977179
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1649977179
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_181
timestamp 1649977179
transform 1 0 17756 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_189
timestamp 1649977179
transform 1 0 18492 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_194
timestamp 1649977179
transform 1 0 18952 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_200
timestamp 1649977179
transform 1 0 19504 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_206
timestamp 1649977179
transform 1 0 20056 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_214
timestamp 1649977179
transform 1 0 20792 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_220
timestamp 1649977179
transform 1 0 21344 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_225
timestamp 1649977179
transform 1 0 21804 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_229
timestamp 1649977179
transform 1 0 22172 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_232
timestamp 1649977179
transform 1 0 22448 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_238
timestamp 1649977179
transform 1 0 23000 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_245
timestamp 1649977179
transform 1 0 23644 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_256
timestamp 1649977179
transform 1 0 24656 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_264
timestamp 1649977179
transform 1 0 25392 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_272
timestamp 1649977179
transform 1 0 26128 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_81_287
timestamp 1649977179
transform 1 0 27508 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_81_297
timestamp 1649977179
transform 1 0 28428 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_306
timestamp 1649977179
transform 1 0 29256 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_317
timestamp 1649977179
transform 1 0 30268 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_324
timestamp 1649977179
transform 1 0 30912 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_330
timestamp 1649977179
transform 1 0 31464 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_344
timestamp 1649977179
transform 1 0 32752 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_354
timestamp 1649977179
transform 1 0 33672 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_360
timestamp 1649977179
transform 1 0 34224 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_369
timestamp 1649977179
transform 1 0 35052 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_375
timestamp 1649977179
transform 1 0 35604 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_381
timestamp 1649977179
transform 1 0 36156 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_387
timestamp 1649977179
transform 1 0 36708 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1649977179
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_395
timestamp 1649977179
transform 1 0 37444 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_401
timestamp 1649977179
transform 1 0 37996 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_413
timestamp 1649977179
transform 1 0 39100 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_425
timestamp 1649977179
transform 1 0 40204 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_437
timestamp 1649977179
transform 1 0 41308 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_445
timestamp 1649977179
transform 1 0 42044 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1649977179
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1649977179
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1649977179
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1649977179
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1649977179
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1649977179
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1649977179
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1649977179
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1649977179
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1649977179
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1649977179
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1649977179
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_81_561
timestamp 1649977179
transform 1 0 52716 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_564
timestamp 1649977179
transform 1 0 52992 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_572
timestamp 1649977179
transform 1 0 53728 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1649977179
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1649977179
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1649977179
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1649977179
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1649977179
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1649977179
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1649977179
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1649977179
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1649977179
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1649977179
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1649977179
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1649977179
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1649977179
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1649977179
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1649977179
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1649977179
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1649977179
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1649977179
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1649977179
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1649977179
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1649977179
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_197
timestamp 1649977179
transform 1 0 19228 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_203
timestamp 1649977179
transform 1 0 19780 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_209
timestamp 1649977179
transform 1 0 20332 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_215
timestamp 1649977179
transform 1 0 20884 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_221
timestamp 1649977179
transform 1 0 21436 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_227
timestamp 1649977179
transform 1 0 21988 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_233
timestamp 1649977179
transform 1 0 22540 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_237
timestamp 1649977179
transform 1 0 22908 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1649977179
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1649977179
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_255
timestamp 1649977179
transform 1 0 24564 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_267
timestamp 1649977179
transform 1 0 25668 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_279
timestamp 1649977179
transform 1 0 26772 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_287
timestamp 1649977179
transform 1 0 27508 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_295
timestamp 1649977179
transform 1 0 28244 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_304
timestamp 1649977179
transform 1 0 29072 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_82_309
timestamp 1649977179
transform 1 0 29532 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_318
timestamp 1649977179
transform 1 0 30360 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_327
timestamp 1649977179
transform 1 0 31188 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_333
timestamp 1649977179
transform 1 0 31740 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_337
timestamp 1649977179
transform 1 0 32108 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_342
timestamp 1649977179
transform 1 0 32568 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_354
timestamp 1649977179
transform 1 0 33672 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_360
timestamp 1649977179
transform 1 0 34224 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_367
timestamp 1649977179
transform 1 0 34868 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_373
timestamp 1649977179
transform 1 0 35420 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_379
timestamp 1649977179
transform 1 0 35972 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_385
timestamp 1649977179
transform 1 0 36524 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_391
timestamp 1649977179
transform 1 0 37076 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_397
timestamp 1649977179
transform 1 0 37628 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_409
timestamp 1649977179
transform 1 0 38732 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_417
timestamp 1649977179
transform 1 0 39468 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1649977179
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1649977179
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1649977179
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1649977179
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1649977179
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1649977179
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1649977179
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1649977179
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1649977179
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1649977179
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1649977179
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1649977179
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1649977179
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1649977179
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1649977179
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_569
timestamp 1649977179
transform 1 0 53452 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_575
timestamp 1649977179
transform 1 0 54004 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1649977179
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1649977179
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1649977179
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1649977179
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1649977179
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1649977179
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1649977179
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1649977179
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1649977179
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1649977179
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1649977179
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1649977179
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1649977179
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1649977179
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1649977179
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1649977179
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1649977179
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1649977179
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1649977179
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1649977179
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1649977179
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_83_205
timestamp 1649977179
transform 1 0 19964 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_208
timestamp 1649977179
transform 1 0 20240 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_214
timestamp 1649977179
transform 1 0 20792 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_220
timestamp 1649977179
transform 1 0 21344 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_83_225
timestamp 1649977179
transform 1 0 21804 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_83_235
timestamp 1649977179
transform 1 0 22724 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_244
timestamp 1649977179
transform 1 0 23552 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_250
timestamp 1649977179
transform 1 0 24104 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_257
timestamp 1649977179
transform 1 0 24748 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_266
timestamp 1649977179
transform 1 0 25576 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_276
timestamp 1649977179
transform 1 0 26496 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_291
timestamp 1649977179
transform 1 0 27876 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_83_299
timestamp 1649977179
transform 1 0 28612 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_311
timestamp 1649977179
transform 1 0 29716 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_319
timestamp 1649977179
transform 1 0 30452 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_328
timestamp 1649977179
transform 1 0 31280 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_83_340
timestamp 1649977179
transform 1 0 32384 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_83_355
timestamp 1649977179
transform 1 0 33764 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_366
timestamp 1649977179
transform 1 0 34776 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_373
timestamp 1649977179
transform 1 0 35420 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_379
timestamp 1649977179
transform 1 0 35972 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1649977179
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1649977179
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_395
timestamp 1649977179
transform 1 0 37444 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_407
timestamp 1649977179
transform 1 0 38548 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_419
timestamp 1649977179
transform 1 0 39652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_431
timestamp 1649977179
transform 1 0 40756 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_443
timestamp 1649977179
transform 1 0 41860 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1649977179
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1649977179
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1649977179
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1649977179
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1649977179
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1649977179
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1649977179
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1649977179
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1649977179
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1649977179
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1649977179
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1649977179
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1649977179
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1649977179
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_83_573
timestamp 1649977179
transform 1 0 53820 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_7
timestamp 1649977179
transform 1 0 1748 0 1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_13
timestamp 1649977179
transform 1 0 2300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_25
timestamp 1649977179
transform 1 0 3404 0 1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1649977179
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1649977179
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1649977179
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1649977179
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1649977179
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1649977179
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1649977179
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1649977179
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1649977179
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1649977179
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1649977179
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1649977179
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1649977179
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1649977179
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1649977179
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1649977179
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1649977179
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1649977179
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1649977179
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_209
timestamp 1649977179
transform 1 0 20332 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_214
timestamp 1649977179
transform 1 0 20792 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_220
timestamp 1649977179
transform 1 0 21344 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_226
timestamp 1649977179
transform 1 0 21896 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_232
timestamp 1649977179
transform 1 0 22448 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_238
timestamp 1649977179
transform 1 0 23000 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_84_248
timestamp 1649977179
transform 1 0 23920 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_253
timestamp 1649977179
transform 1 0 24380 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_260
timestamp 1649977179
transform 1 0 25024 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_267
timestamp 1649977179
transform 1 0 25668 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_271
timestamp 1649977179
transform 1 0 26036 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_279
timestamp 1649977179
transform 1 0 26772 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_291
timestamp 1649977179
transform 1 0 27876 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_304
timestamp 1649977179
transform 1 0 29072 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_309
timestamp 1649977179
transform 1 0 29532 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_318
timestamp 1649977179
transform 1 0 30360 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_328
timestamp 1649977179
transform 1 0 31280 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_334
timestamp 1649977179
transform 1 0 31832 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_344
timestamp 1649977179
transform 1 0 32752 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_355
timestamp 1649977179
transform 1 0 33764 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1649977179
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_369
timestamp 1649977179
transform 1 0 35052 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_376
timestamp 1649977179
transform 1 0 35696 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_382
timestamp 1649977179
transform 1 0 36248 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_388
timestamp 1649977179
transform 1 0 36800 0 1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_394
timestamp 1649977179
transform 1 0 37352 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_406
timestamp 1649977179
transform 1 0 38456 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_84_418
timestamp 1649977179
transform 1 0 39560 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1649977179
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1649977179
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1649977179
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1649977179
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1649977179
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1649977179
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1649977179
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1649977179
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1649977179
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1649977179
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1649977179
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1649977179
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1649977179
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1649977179
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1649977179
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_569
timestamp 1649977179
transform 1 0 53452 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_575
timestamp 1649977179
transform 1 0 54004 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1649977179
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1649977179
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1649977179
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1649977179
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1649977179
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1649977179
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1649977179
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1649977179
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1649977179
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1649977179
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1649977179
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1649977179
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1649977179
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1649977179
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1649977179
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1649977179
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1649977179
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1649977179
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1649977179
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1649977179
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1649977179
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1649977179
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_85_217
timestamp 1649977179
transform 1 0 21068 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_220
timestamp 1649977179
transform 1 0 21344 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_227
timestamp 1649977179
transform 1 0 21988 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_233
timestamp 1649977179
transform 1 0 22540 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_239
timestamp 1649977179
transform 1 0 23092 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_250
timestamp 1649977179
transform 1 0 24104 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_85_264
timestamp 1649977179
transform 1 0 25392 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_272
timestamp 1649977179
transform 1 0 26128 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_276
timestamp 1649977179
transform 1 0 26496 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_288
timestamp 1649977179
transform 1 0 27600 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_85_303
timestamp 1649977179
transform 1 0 28980 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_309
timestamp 1649977179
transform 1 0 29532 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_85_319
timestamp 1649977179
transform 1 0 30452 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_326
timestamp 1649977179
transform 1 0 31096 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_332
timestamp 1649977179
transform 1 0 31648 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_339
timestamp 1649977179
transform 1 0 32292 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_345
timestamp 1649977179
transform 1 0 32844 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_351
timestamp 1649977179
transform 1 0 33396 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_357
timestamp 1649977179
transform 1 0 33948 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_365
timestamp 1649977179
transform 1 0 34684 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_372
timestamp 1649977179
transform 1 0 35328 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_378
timestamp 1649977179
transform 1 0 35880 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_384
timestamp 1649977179
transform 1 0 36432 0 -1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1649977179
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1649977179
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1649977179
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1649977179
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1649977179
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1649977179
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1649977179
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1649977179
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1649977179
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1649977179
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1649977179
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1649977179
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1649977179
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1649977179
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1649977179
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1649977179
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1649977179
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1649977179
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_561
timestamp 1649977179
transform 1 0 52716 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_564
timestamp 1649977179
transform 1 0 52992 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_572
timestamp 1649977179
transform 1 0 53728 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1649977179
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1649977179
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1649977179
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1649977179
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1649977179
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1649977179
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1649977179
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1649977179
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1649977179
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1649977179
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1649977179
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1649977179
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1649977179
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1649977179
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1649977179
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1649977179
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1649977179
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1649977179
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1649977179
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1649977179
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1649977179
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1649977179
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1649977179
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_86_221
timestamp 1649977179
transform 1 0 21436 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_225
timestamp 1649977179
transform 1 0 21804 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_231
timestamp 1649977179
transform 1 0 22356 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_237
timestamp 1649977179
transform 1 0 22908 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_248
timestamp 1649977179
transform 1 0 23920 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_259
timestamp 1649977179
transform 1 0 24932 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_266
timestamp 1649977179
transform 1 0 25576 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_273
timestamp 1649977179
transform 1 0 26220 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_282
timestamp 1649977179
transform 1 0 27048 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_288
timestamp 1649977179
transform 1 0 27600 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_295
timestamp 1649977179
transform 1 0 28244 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_86_304
timestamp 1649977179
transform 1 0 29072 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_315
timestamp 1649977179
transform 1 0 30084 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_324
timestamp 1649977179
transform 1 0 30912 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_331
timestamp 1649977179
transform 1 0 31556 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_86_344
timestamp 1649977179
transform 1 0 32752 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_356
timestamp 1649977179
transform 1 0 33856 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_86_370
timestamp 1649977179
transform 1 0 35144 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_377
timestamp 1649977179
transform 1 0 35788 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_383
timestamp 1649977179
transform 1 0 36340 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_389
timestamp 1649977179
transform 1 0 36892 0 1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_395
timestamp 1649977179
transform 1 0 37444 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_407
timestamp 1649977179
transform 1 0 38548 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1649977179
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1649977179
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1649977179
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1649977179
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1649977179
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1649977179
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1649977179
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1649977179
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1649977179
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1649977179
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1649977179
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1649977179
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1649977179
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1649977179
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1649977179
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1649977179
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_569
timestamp 1649977179
transform 1 0 53452 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_575
timestamp 1649977179
transform 1 0 54004 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1649977179
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1649977179
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1649977179
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1649977179
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1649977179
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1649977179
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1649977179
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1649977179
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1649977179
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1649977179
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1649977179
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1649977179
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1649977179
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1649977179
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1649977179
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1649977179
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1649977179
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1649977179
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1649977179
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1649977179
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1649977179
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1649977179
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_87_217
timestamp 1649977179
transform 1 0 21068 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_220
timestamp 1649977179
transform 1 0 21344 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_87_225
timestamp 1649977179
transform 1 0 21804 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_87_230
timestamp 1649977179
transform 1 0 22264 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_87_237
timestamp 1649977179
transform 1 0 22908 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_87_248
timestamp 1649977179
transform 1 0 23920 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_87_255
timestamp 1649977179
transform 1 0 24564 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_87_266
timestamp 1649977179
transform 1 0 25576 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_270
timestamp 1649977179
transform 1 0 25944 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_276
timestamp 1649977179
transform 1 0 26496 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_87_283
timestamp 1649977179
transform 1 0 27140 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_87_291
timestamp 1649977179
transform 1 0 27876 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_294
timestamp 1649977179
transform 1 0 28152 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_87_315
timestamp 1649977179
transform 1 0 30084 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_87_323
timestamp 1649977179
transform 1 0 30820 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_87_330
timestamp 1649977179
transform 1 0 31464 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_87_356
timestamp 1649977179
transform 1 0 33856 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_365
timestamp 1649977179
transform 1 0 34684 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_371
timestamp 1649977179
transform 1 0 35236 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_377
timestamp 1649977179
transform 1 0 35788 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_87_383
timestamp 1649977179
transform 1 0 36340 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1649977179
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1649977179
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1649977179
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1649977179
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1649977179
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1649977179
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1649977179
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1649977179
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1649977179
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1649977179
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1649977179
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1649977179
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1649977179
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1649977179
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1649977179
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1649977179
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1649977179
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1649977179
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1649977179
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1649977179
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_87_573
timestamp 1649977179
transform 1 0 53820 0 -1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_88_5
timestamp 1649977179
transform 1 0 1564 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_17
timestamp 1649977179
transform 1 0 2668 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_88_25
timestamp 1649977179
transform 1 0 3404 0 1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1649977179
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1649977179
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1649977179
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1649977179
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1649977179
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1649977179
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1649977179
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1649977179
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1649977179
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1649977179
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1649977179
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1649977179
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1649977179
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1649977179
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1649977179
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1649977179
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1649977179
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1649977179
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1649977179
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_209
timestamp 1649977179
transform 1 0 20332 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_213
timestamp 1649977179
transform 1 0 20700 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_216
timestamp 1649977179
transform 1 0 20976 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_222
timestamp 1649977179
transform 1 0 21528 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_228
timestamp 1649977179
transform 1 0 22080 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_237
timestamp 1649977179
transform 1 0 22908 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_248
timestamp 1649977179
transform 1 0 23920 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_253
timestamp 1649977179
transform 1 0 24380 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_257
timestamp 1649977179
transform 1 0 24748 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_263
timestamp 1649977179
transform 1 0 25300 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_274
timestamp 1649977179
transform 1 0 26312 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_88_284
timestamp 1649977179
transform 1 0 27232 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_88_292
timestamp 1649977179
transform 1 0 27968 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_88_295
timestamp 1649977179
transform 1 0 28244 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_88_303
timestamp 1649977179
transform 1 0 28980 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1649977179
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_309
timestamp 1649977179
transform 1 0 29532 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_88_319
timestamp 1649977179
transform 1 0 30452 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_325
timestamp 1649977179
transform 1 0 31004 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_88_333
timestamp 1649977179
transform 1 0 31740 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_88_344
timestamp 1649977179
transform 1 0 32752 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_353
timestamp 1649977179
transform 1 0 33580 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_360
timestamp 1649977179
transform 1 0 34224 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_367
timestamp 1649977179
transform 1 0 34868 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_373
timestamp 1649977179
transform 1 0 35420 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_379
timestamp 1649977179
transform 1 0 35972 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_391
timestamp 1649977179
transform 1 0 37076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_403
timestamp 1649977179
transform 1 0 38180 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_415
timestamp 1649977179
transform 1 0 39284 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1649977179
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1649977179
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1649977179
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1649977179
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1649977179
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1649977179
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1649977179
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1649977179
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1649977179
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1649977179
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1649977179
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1649977179
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1649977179
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1649977179
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1649977179
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1649977179
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_569
timestamp 1649977179
transform 1 0 53452 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_575
timestamp 1649977179
transform 1 0 54004 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_7
timestamp 1649977179
transform 1 0 1748 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_19
timestamp 1649977179
transform 1 0 2852 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_31
timestamp 1649977179
transform 1 0 3956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_43
timestamp 1649977179
transform 1 0 5060 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1649977179
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1649977179
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1649977179
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1649977179
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1649977179
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1649977179
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1649977179
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1649977179
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1649977179
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1649977179
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1649977179
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1649977179
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1649977179
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1649977179
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1649977179
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1649977179
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1649977179
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1649977179
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1649977179
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_225
timestamp 1649977179
transform 1 0 21804 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_229
timestamp 1649977179
transform 1 0 22172 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_236
timestamp 1649977179
transform 1 0 22816 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_248
timestamp 1649977179
transform 1 0 23920 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_254
timestamp 1649977179
transform 1 0 24472 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_265
timestamp 1649977179
transform 1 0 25484 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1649977179
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1649977179
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_89_281
timestamp 1649977179
transform 1 0 26956 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_89_284
timestamp 1649977179
transform 1 0 27232 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_290
timestamp 1649977179
transform 1 0 27784 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_293
timestamp 1649977179
transform 1 0 28060 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_89_299
timestamp 1649977179
transform 1 0 28612 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_89_307
timestamp 1649977179
transform 1 0 29348 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_310
timestamp 1649977179
transform 1 0 29624 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_318
timestamp 1649977179
transform 1 0 30360 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_89_327
timestamp 1649977179
transform 1 0 31188 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1649977179
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_341
timestamp 1649977179
transform 1 0 32476 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_89_347
timestamp 1649977179
transform 1 0 33028 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_89_355
timestamp 1649977179
transform 1 0 33764 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_89_370
timestamp 1649977179
transform 1 0 35144 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_376
timestamp 1649977179
transform 1 0 35696 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_382
timestamp 1649977179
transform 1 0 36248 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_388
timestamp 1649977179
transform 1 0 36800 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1649977179
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1649977179
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1649977179
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1649977179
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1649977179
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1649977179
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1649977179
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1649977179
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1649977179
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1649977179
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1649977179
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1649977179
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1649977179
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1649977179
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1649977179
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1649977179
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1649977179
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1649977179
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_89_561
timestamp 1649977179
transform 1 0 52716 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_564
timestamp 1649977179
transform 1 0 52992 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_572
timestamp 1649977179
transform 1 0 53728 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1649977179
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1649977179
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1649977179
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1649977179
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1649977179
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1649977179
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1649977179
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1649977179
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1649977179
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1649977179
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1649977179
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1649977179
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1649977179
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1649977179
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1649977179
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1649977179
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1649977179
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1649977179
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1649977179
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1649977179
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1649977179
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1649977179
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1649977179
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_221
timestamp 1649977179
transform 1 0 21436 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_227
timestamp 1649977179
transform 1 0 21988 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_230
timestamp 1649977179
transform 1 0 22264 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_236
timestamp 1649977179
transform 1 0 22816 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_90_244
timestamp 1649977179
transform 1 0 23552 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_90_253
timestamp 1649977179
transform 1 0 24380 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_90_259
timestamp 1649977179
transform 1 0 24932 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_90_268
timestamp 1649977179
transform 1 0 25760 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_272
timestamp 1649977179
transform 1 0 26128 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_275
timestamp 1649977179
transform 1 0 26404 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_281
timestamp 1649977179
transform 1 0 26956 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_289
timestamp 1649977179
transform 1 0 27692 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_90_295
timestamp 1649977179
transform 1 0 28244 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_301
timestamp 1649977179
transform 1 0 28796 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_304
timestamp 1649977179
transform 1 0 29072 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_311
timestamp 1649977179
transform 1 0 29716 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_317
timestamp 1649977179
transform 1 0 30268 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_324
timestamp 1649977179
transform 1 0 30912 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_331
timestamp 1649977179
transform 1 0 31556 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_337
timestamp 1649977179
transform 1 0 32108 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_90_343
timestamp 1649977179
transform 1 0 32660 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_90_356
timestamp 1649977179
transform 1 0 33856 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_90_372
timestamp 1649977179
transform 1 0 35328 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_378
timestamp 1649977179
transform 1 0 35880 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_384
timestamp 1649977179
transform 1 0 36432 0 1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_90_390
timestamp 1649977179
transform 1 0 36984 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_402
timestamp 1649977179
transform 1 0 38088 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_414
timestamp 1649977179
transform 1 0 39192 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1649977179
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1649977179
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1649977179
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1649977179
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1649977179
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1649977179
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1649977179
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1649977179
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1649977179
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1649977179
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1649977179
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1649977179
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1649977179
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1649977179
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1649977179
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_569
timestamp 1649977179
transform 1 0 53452 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_575
timestamp 1649977179
transform 1 0 54004 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_5
timestamp 1649977179
transform 1 0 1564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_17
timestamp 1649977179
transform 1 0 2668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_29
timestamp 1649977179
transform 1 0 3772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_41
timestamp 1649977179
transform 1 0 4876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_53
timestamp 1649977179
transform 1 0 5980 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1649977179
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1649977179
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1649977179
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1649977179
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1649977179
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1649977179
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1649977179
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1649977179
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1649977179
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1649977179
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1649977179
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1649977179
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1649977179
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1649977179
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1649977179
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1649977179
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1649977179
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1649977179
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_225
timestamp 1649977179
transform 1 0 21804 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_233
timestamp 1649977179
transform 1 0 22540 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_91_238
timestamp 1649977179
transform 1 0 23000 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_251
timestamp 1649977179
transform 1 0 24196 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_91_262
timestamp 1649977179
transform 1 0 25208 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_270
timestamp 1649977179
transform 1 0 25944 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_276
timestamp 1649977179
transform 1 0 26496 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_281
timestamp 1649977179
transform 1 0 26956 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_304
timestamp 1649977179
transform 1 0 29072 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_313
timestamp 1649977179
transform 1 0 29900 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_91_319
timestamp 1649977179
transform 1 0 30452 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_91_331
timestamp 1649977179
transform 1 0 31556 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1649977179
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_339
timestamp 1649977179
transform 1 0 32292 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_345
timestamp 1649977179
transform 1 0 32844 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_357
timestamp 1649977179
transform 1 0 33948 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_368
timestamp 1649977179
transform 1 0 34960 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_378
timestamp 1649977179
transform 1 0 35880 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_91_384
timestamp 1649977179
transform 1 0 36432 0 -1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_91_395
timestamp 1649977179
transform 1 0 37444 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_407
timestamp 1649977179
transform 1 0 38548 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_419
timestamp 1649977179
transform 1 0 39652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_431
timestamp 1649977179
transform 1 0 40756 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_443
timestamp 1649977179
transform 1 0 41860 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1649977179
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1649977179
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1649977179
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1649977179
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1649977179
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1649977179
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1649977179
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1649977179
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1649977179
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1649977179
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1649977179
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1649977179
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1649977179
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1649977179
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_573
timestamp 1649977179
transform 1 0 53820 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_92_7
timestamp 1649977179
transform 1 0 1748 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_19
timestamp 1649977179
transform 1 0 2852 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1649977179
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1649977179
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1649977179
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1649977179
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1649977179
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1649977179
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1649977179
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1649977179
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1649977179
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1649977179
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1649977179
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1649977179
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1649977179
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1649977179
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1649977179
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1649977179
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1649977179
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1649977179
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1649977179
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1649977179
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1649977179
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1649977179
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1649977179
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_248
timestamp 1649977179
transform 1 0 23920 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_92_258
timestamp 1649977179
transform 1 0 24840 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_264
timestamp 1649977179
transform 1 0 25392 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_272
timestamp 1649977179
transform 1 0 26128 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_283
timestamp 1649977179
transform 1 0 27140 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_92_293
timestamp 1649977179
transform 1 0 28060 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_299
timestamp 1649977179
transform 1 0 28612 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_304
timestamp 1649977179
transform 1 0 29072 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_317
timestamp 1649977179
transform 1 0 30268 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_326
timestamp 1649977179
transform 1 0 31096 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_335
timestamp 1649977179
transform 1 0 31924 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_339
timestamp 1649977179
transform 1 0 32292 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_343
timestamp 1649977179
transform 1 0 32660 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_360
timestamp 1649977179
transform 1 0 34224 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_372
timestamp 1649977179
transform 1 0 35328 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_378
timestamp 1649977179
transform 1 0 35880 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_384
timestamp 1649977179
transform 1 0 36432 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_396
timestamp 1649977179
transform 1 0 37536 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_408
timestamp 1649977179
transform 1 0 38640 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1649977179
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1649977179
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1649977179
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1649977179
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1649977179
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1649977179
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1649977179
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1649977179
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1649977179
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1649977179
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1649977179
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1649977179
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1649977179
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1649977179
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1649977179
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_569
timestamp 1649977179
transform 1 0 53452 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_575
timestamp 1649977179
transform 1 0 54004 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_5
timestamp 1649977179
transform 1 0 1564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_17
timestamp 1649977179
transform 1 0 2668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_29
timestamp 1649977179
transform 1 0 3772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_41
timestamp 1649977179
transform 1 0 4876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_93_53
timestamp 1649977179
transform 1 0 5980 0 -1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1649977179
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1649977179
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1649977179
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1649977179
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1649977179
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1649977179
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1649977179
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1649977179
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1649977179
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1649977179
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1649977179
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1649977179
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1649977179
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1649977179
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1649977179
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1649977179
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1649977179
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1649977179
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1649977179
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_237
timestamp 1649977179
transform 1 0 22908 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_245
timestamp 1649977179
transform 1 0 23644 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_250
timestamp 1649977179
transform 1 0 24104 0 -1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_93_260
timestamp 1649977179
transform 1 0 25024 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_274
timestamp 1649977179
transform 1 0 26312 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_93_283
timestamp 1649977179
transform 1 0 27140 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_93_296
timestamp 1649977179
transform 1 0 28336 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_319
timestamp 1649977179
transform 1 0 30452 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_93_330
timestamp 1649977179
transform 1 0 31464 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_93_343
timestamp 1649977179
transform 1 0 32660 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_93_357
timestamp 1649977179
transform 1 0 33948 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_367
timestamp 1649977179
transform 1 0 34868 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1649977179
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1649977179
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1649977179
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1649977179
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1649977179
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1649977179
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1649977179
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1649977179
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1649977179
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1649977179
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1649977179
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1649977179
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1649977179
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1649977179
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1649977179
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1649977179
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1649977179
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1649977179
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1649977179
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1649977179
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1649977179
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_93_561
timestamp 1649977179
transform 1 0 52716 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_564
timestamp 1649977179
transform 1 0 52992 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_572
timestamp 1649977179
transform 1 0 53728 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_3
timestamp 1649977179
transform 1 0 1380 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_7
timestamp 1649977179
transform 1 0 1748 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_19
timestamp 1649977179
transform 1 0 2852 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1649977179
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1649977179
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1649977179
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1649977179
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1649977179
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1649977179
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1649977179
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1649977179
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1649977179
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1649977179
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1649977179
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1649977179
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1649977179
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1649977179
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1649977179
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1649977179
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1649977179
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1649977179
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1649977179
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1649977179
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1649977179
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1649977179
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1649977179
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1649977179
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1649977179
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_255
timestamp 1649977179
transform 1 0 24564 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_267
timestamp 1649977179
transform 1 0 25668 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_279
timestamp 1649977179
transform 1 0 26772 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_296
timestamp 1649977179
transform 1 0 28336 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_300
timestamp 1649977179
transform 1 0 28704 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_304
timestamp 1649977179
transform 1 0 29072 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_316
timestamp 1649977179
transform 1 0 30176 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_323
timestamp 1649977179
transform 1 0 30820 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_327
timestamp 1649977179
transform 1 0 31188 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_345
timestamp 1649977179
transform 1 0 32844 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_94_356
timestamp 1649977179
transform 1 0 33856 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1649977179
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1649977179
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1649977179
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1649977179
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1649977179
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1649977179
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1649977179
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_433
timestamp 1649977179
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_445
timestamp 1649977179
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_457
timestamp 1649977179
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1649977179
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1649977179
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1649977179
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1649977179
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1649977179
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1649977179
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1649977179
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1649977179
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1649977179
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1649977179
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_557
timestamp 1649977179
transform 1 0 52348 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_561
timestamp 1649977179
transform 1 0 52716 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_564
timestamp 1649977179
transform 1 0 52992 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_572
timestamp 1649977179
transform 1 0 53728 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_3
timestamp 1649977179
transform 1 0 1380 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_11
timestamp 1649977179
transform 1 0 2116 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_17
timestamp 1649977179
transform 1 0 2668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_31
timestamp 1649977179
transform 1 0 3956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_43
timestamp 1649977179
transform 1 0 5060 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1649977179
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_57
timestamp 1649977179
transform 1 0 6348 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_63
timestamp 1649977179
transform 1 0 6900 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_75
timestamp 1649977179
transform 1 0 8004 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_87
timestamp 1649977179
transform 1 0 9108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_99
timestamp 1649977179
transform 1 0 10212 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1649977179
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_115
timestamp 1649977179
transform 1 0 11684 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_127
timestamp 1649977179
transform 1 0 12788 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_139
timestamp 1649977179
transform 1 0 13892 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_151
timestamp 1649977179
transform 1 0 14996 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_163
timestamp 1649977179
transform 1 0 16100 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1649977179
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1649977179
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1649977179
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1649977179
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1649977179
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1649977179
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1649977179
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_225
timestamp 1649977179
transform 1 0 21804 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_229
timestamp 1649977179
transform 1 0 22172 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_237
timestamp 1649977179
transform 1 0 22908 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_241
timestamp 1649977179
transform 1 0 23276 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_253
timestamp 1649977179
transform 1 0 24380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_265
timestamp 1649977179
transform 1 0 25484 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_277
timestamp 1649977179
transform 1 0 26588 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_95_297
timestamp 1649977179
transform 1 0 28428 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_303
timestamp 1649977179
transform 1 0 28980 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_310
timestamp 1649977179
transform 1 0 29624 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_316
timestamp 1649977179
transform 1 0 30176 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_319
timestamp 1649977179
transform 1 0 30452 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_325
timestamp 1649977179
transform 1 0 31004 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_331
timestamp 1649977179
transform 1 0 31556 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1649977179
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_95_337
timestamp 1649977179
transform 1 0 32108 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_95_345
timestamp 1649977179
transform 1 0 32844 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_352
timestamp 1649977179
transform 1 0 33488 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_364
timestamp 1649977179
transform 1 0 34592 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_95_369
timestamp 1649977179
transform 1 0 35052 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_377
timestamp 1649977179
transform 1 0 35788 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_381
timestamp 1649977179
transform 1 0 36156 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_95_389
timestamp 1649977179
transform 1 0 36892 0 -1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1649977179
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_405
timestamp 1649977179
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_417
timestamp 1649977179
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_429
timestamp 1649977179
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1649977179
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1649977179
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1649977179
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1649977179
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_473
timestamp 1649977179
transform 1 0 44620 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_479
timestamp 1649977179
transform 1 0 45172 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_491
timestamp 1649977179
transform 1 0 46276 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1649977179
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1649977179
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1649977179
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1649977179
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1649977179
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1649977179
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1649977179
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_95_561
timestamp 1649977179
transform 1 0 52716 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_564
timestamp 1649977179
transform 1 0 52992 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_572
timestamp 1649977179
transform 1 0 53728 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_13
timestamp 1649977179
transform 1 0 2300 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_96_21
timestamp 1649977179
transform 1 0 3036 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1649977179
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_96_29
timestamp 1649977179
transform 1 0 3772 0 1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1649977179
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_96_53
timestamp 1649977179
transform 1 0 5980 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_96_61
timestamp 1649977179
transform 1 0 6716 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_96_69
timestamp 1649977179
transform 1 0 7452 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1649977179
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1649977179
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1649977179
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_97
timestamp 1649977179
transform 1 0 10028 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_108
timestamp 1649977179
transform 1 0 11040 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_96_113
timestamp 1649977179
transform 1 0 11500 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_96_118
timestamp 1649977179
transform 1 0 11960 0 1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_126
timestamp 1649977179
transform 1 0 12696 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_96_138
timestamp 1649977179
transform 1 0 13800 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_141
timestamp 1649977179
transform 1 0 14076 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_147
timestamp 1649977179
transform 1 0 14628 0 1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1649977179
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_96_165
timestamp 1649977179
transform 1 0 16284 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_96_169
timestamp 1649977179
transform 1 0 16652 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_175
timestamp 1649977179
transform 1 0 17204 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_96_181
timestamp 1649977179
transform 1 0 17756 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_189
timestamp 1649977179
transform 1 0 18492 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_192
timestamp 1649977179
transform 1 0 18768 0 1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_207
timestamp 1649977179
transform 1 0 20148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_219
timestamp 1649977179
transform 1 0 21252 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_223
timestamp 1649977179
transform 1 0 21620 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_225
timestamp 1649977179
transform 1 0 21804 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_96_233
timestamp 1649977179
transform 1 0 22540 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_96_247
timestamp 1649977179
transform 1 0 23828 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1649977179
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_96_253
timestamp 1649977179
transform 1 0 24380 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_96_258
timestamp 1649977179
transform 1 0 24840 0 1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_266
timestamp 1649977179
transform 1 0 25576 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_96_278
timestamp 1649977179
transform 1 0 26680 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_96_281
timestamp 1649977179
transform 1 0 26956 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_96_286
timestamp 1649977179
transform 1 0 27416 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_96_300
timestamp 1649977179
transform 1 0 28704 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_96_309
timestamp 1649977179
transform 1 0 29532 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_315
timestamp 1649977179
transform 1 0 30084 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_321
timestamp 1649977179
transform 1 0 30636 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_96_327
timestamp 1649977179
transform 1 0 31188 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_335
timestamp 1649977179
transform 1 0 31924 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_337
timestamp 1649977179
transform 1 0 32108 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_344
timestamp 1649977179
transform 1 0 32752 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_350
timestamp 1649977179
transform 1 0 33304 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_96_356
timestamp 1649977179
transform 1 0 33856 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_96_365
timestamp 1649977179
transform 1 0 34684 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_96_373
timestamp 1649977179
transform 1 0 35420 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_96_385
timestamp 1649977179
transform 1 0 36524 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_391
timestamp 1649977179
transform 1 0 37076 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_393
timestamp 1649977179
transform 1 0 37260 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_96_401
timestamp 1649977179
transform 1 0 37996 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_405
timestamp 1649977179
transform 1 0 38364 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1649977179
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1649977179
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_96_421
timestamp 1649977179
transform 1 0 39836 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_96_426
timestamp 1649977179
transform 1 0 40296 0 1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_434
timestamp 1649977179
transform 1 0 41032 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_96_446
timestamp 1649977179
transform 1 0 42136 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_449
timestamp 1649977179
transform 1 0 42412 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_454
timestamp 1649977179
transform 1 0 42872 0 1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_460
timestamp 1649977179
transform 1 0 43424 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_472
timestamp 1649977179
transform 1 0 44528 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_477
timestamp 1649977179
transform 1 0 44988 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_96_489
timestamp 1649977179
transform 1 0 46092 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_497
timestamp 1649977179
transform 1 0 46828 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_500
timestamp 1649977179
transform 1 0 47104 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_96_509
timestamp 1649977179
transform 1 0 47932 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_96_517
timestamp 1649977179
transform 1 0 48668 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1649977179
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1649977179
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_533
timestamp 1649977179
transform 1 0 50140 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_96_541
timestamp 1649977179
transform 1 0 50876 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_545
timestamp 1649977179
transform 1 0 51244 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_96_553
timestamp 1649977179
transform 1 0 51980 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_559
timestamp 1649977179
transform 1 0 52532 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_96_561
timestamp 1649977179
transform 1 0 52716 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_564
timestamp 1649977179
transform 1 0 52992 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_572
timestamp 1649977179
transform 1 0 53728 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 54372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 54372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 54372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 54372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 54372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 54372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 54372 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 54372 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 54372 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 54372 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 54372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 54372 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 54372 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 54372 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 54372 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 54372 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 54372 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 54372 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 54372 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 54372 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 54372 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 54372 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 54372 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 54372 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 54372 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 54372 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 54372 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 54372 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 54372 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 54372 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 54372 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 54372 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 54372 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 54372 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 54372 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 54372 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 54372 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 54372 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 54372 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 54372 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 54372 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 54372 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 54372 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 54372 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 54372 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 54372 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 54372 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 54372 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 54372 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 54372 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 54372 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 54372 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 54372 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 54372 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 54372 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 54372 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 54372 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 54372 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 54372 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 54372 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 54372 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 54372 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 54372 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 54372 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 54372 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1649977179
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1649977179
transform -1 0 54372 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1649977179
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1649977179
transform -1 0 54372 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1649977179
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1649977179
transform -1 0 54372 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1649977179
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1649977179
transform -1 0 54372 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1649977179
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1649977179
transform -1 0 54372 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1649977179
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1649977179
transform -1 0 54372 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1649977179
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1649977179
transform -1 0 54372 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1649977179
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1649977179
transform -1 0 54372 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1649977179
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1649977179
transform -1 0 54372 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1649977179
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1649977179
transform -1 0 54372 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1649977179
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1649977179
transform -1 0 54372 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1649977179
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1649977179
transform -1 0 54372 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1649977179
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1649977179
transform -1 0 54372 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1649977179
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1649977179
transform -1 0 54372 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1649977179
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1649977179
transform -1 0 54372 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1649977179
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1649977179
transform -1 0 54372 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1649977179
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1649977179
transform -1 0 54372 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1649977179
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1649977179
transform -1 0 54372 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1649977179
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1649977179
transform -1 0 54372 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1649977179
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1649977179
transform -1 0 54372 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1649977179
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1649977179
transform -1 0 54372 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1649977179
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1649977179
transform -1 0 54372 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1649977179
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1649977179
transform -1 0 54372 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1649977179
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1649977179
transform -1 0 54372 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1649977179
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1649977179
transform -1 0 54372 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1649977179
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1649977179
transform -1 0 54372 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1649977179
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1649977179
transform -1 0 54372 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1649977179
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1649977179
transform -1 0 54372 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1649977179
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1649977179
transform -1 0 54372 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1649977179
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1649977179
transform -1 0 54372 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1649977179
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1649977179
transform -1 0 54372 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1649977179
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1649977179
transform -1 0 54372 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1649977179
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1649977179
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1649977179
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1649977179
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1649977179
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1649977179
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1649977179
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1649977179
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1649977179
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1649977179
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1649977179
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1649977179
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1649977179
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1649977179
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1649977179
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1649977179
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1649977179
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1649977179
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1649977179
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1649977179
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1649977179
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1649977179
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1649977179
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1649977179
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1649977179
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1649977179
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1649977179
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1649977179
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1649977179
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1649977179
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1649977179
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1649977179
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1649977179
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1649977179
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1649977179
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1649977179
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1649977179
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1649977179
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1649977179
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1649977179
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1649977179
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1649977179
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1649977179
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1649977179
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1649977179
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1649977179
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1649977179
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1649977179
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1649977179
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1649977179
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1649977179
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1649977179
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1649977179
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1649977179
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1649977179
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1649977179
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1649977179
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1649977179
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1649977179
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1649977179
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1649977179
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1649977179
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1649977179
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1649977179
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1649977179
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1649977179
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1649977179
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1649977179
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1649977179
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1649977179
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1649977179
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1649977179
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1649977179
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1649977179
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1649977179
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1649977179
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1649977179
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1649977179
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1649977179
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1649977179
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1649977179
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1649977179
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1649977179
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1649977179
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1649977179
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1649977179
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1649977179
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1649977179
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1649977179
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1649977179
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1649977179
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1649977179
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1649977179
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1649977179
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1649977179
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1649977179
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1649977179
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1649977179
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1649977179
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1649977179
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1649977179
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1649977179
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1649977179
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1649977179
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1649977179
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1649977179
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1649977179
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1649977179
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1649977179
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1649977179
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1649977179
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1649977179
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1649977179
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1649977179
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1649977179
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1649977179
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1649977179
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1649977179
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1649977179
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1649977179
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1649977179
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1649977179
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1649977179
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1649977179
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1649977179
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1649977179
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1649977179
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1649977179
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1649977179
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1649977179
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1649977179
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1649977179
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1649977179
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1649977179
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1649977179
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1649977179
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1649977179
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1649977179
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1649977179
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1649977179
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1649977179
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1649977179
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1649977179
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1649977179
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1649977179
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1649977179
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1649977179
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1649977179
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1649977179
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1649977179
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1649977179
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1649977179
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1649977179
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1649977179
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1649977179
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1649977179
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1649977179
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1649977179
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1649977179
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1649977179
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1649977179
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1649977179
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1649977179
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1649977179
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1649977179
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1649977179
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1649977179
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1649977179
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1649977179
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1649977179
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1649977179
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1649977179
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1649977179
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1649977179
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1649977179
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1649977179
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1649977179
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1649977179
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1649977179
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1649977179
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1649977179
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1649977179
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1649977179
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1649977179
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1649977179
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1649977179
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1649977179
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1649977179
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1649977179
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1649977179
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1649977179
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1649977179
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1649977179
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1649977179
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1649977179
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1649977179
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1649977179
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1649977179
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1649977179
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1649977179
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1649977179
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1649977179
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1649977179
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1649977179
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1649977179
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1649977179
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1649977179
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1649977179
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1649977179
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1649977179
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1649977179
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1649977179
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1649977179
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1649977179
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1649977179
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1649977179
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1649977179
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1649977179
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1649977179
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1649977179
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1649977179
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1649977179
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1649977179
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1649977179
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1649977179
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1649977179
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1649977179
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1649977179
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1649977179
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1649977179
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1649977179
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1649977179
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1649977179
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1649977179
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1649977179
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1649977179
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1649977179
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1649977179
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1649977179
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1649977179
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1649977179
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1649977179
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1649977179
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1649977179
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1649977179
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1649977179
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1649977179
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1649977179
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1649977179
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1649977179
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1649977179
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1649977179
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1649977179
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1649977179
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1649977179
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1649977179
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1649977179
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1649977179
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1649977179
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1649977179
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1649977179
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1649977179
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1649977179
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1649977179
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1649977179
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1649977179
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1649977179
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1649977179
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1649977179
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1649977179
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1649977179
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1649977179
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1649977179
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1649977179
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1649977179
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1649977179
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1649977179
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1649977179
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1649977179
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1649977179
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1649977179
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1649977179
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1649977179
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1649977179
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1649977179
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1649977179
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1649977179
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1649977179
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1649977179
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1649977179
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1649977179
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1649977179
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1649977179
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1649977179
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1649977179
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1649977179
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1649977179
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1649977179
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1649977179
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1649977179
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1649977179
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1649977179
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1649977179
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1649977179
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1649977179
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1649977179
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1649977179
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1649977179
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1649977179
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1649977179
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1649977179
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1649977179
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1649977179
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1649977179
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1649977179
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1649977179
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1649977179
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1649977179
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1649977179
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1649977179
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1649977179
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1649977179
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1649977179
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1649977179
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1649977179
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1649977179
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1649977179
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1649977179
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1649977179
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1649977179
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1649977179
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1649977179
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1649977179
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1649977179
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1649977179
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1649977179
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1649977179
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1649977179
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1649977179
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1649977179
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1649977179
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1649977179
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1649977179
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1649977179
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1649977179
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1649977179
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1649977179
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1649977179
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1649977179
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1649977179
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1649977179
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1649977179
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1649977179
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1649977179
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1649977179
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1649977179
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1649977179
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1649977179
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1649977179
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1649977179
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1649977179
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1649977179
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1649977179
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1649977179
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1649977179
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1649977179
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1649977179
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1649977179
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1649977179
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1649977179
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1649977179
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1649977179
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1649977179
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1649977179
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1649977179
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1649977179
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1649977179
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1649977179
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1649977179
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1649977179
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1649977179
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1649977179
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1649977179
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1649977179
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1649977179
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1649977179
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1649977179
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1649977179
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1649977179
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1649977179
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1649977179
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1649977179
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1649977179
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1649977179
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1649977179
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1649977179
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1649977179
transform 1 0 6256 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1649977179
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1649977179
transform 1 0 11408 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1649977179
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1649977179
transform 1 0 16560 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1649977179
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1649977179
transform 1 0 21712 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1649977179
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1649977179
transform 1 0 26864 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1649977179
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1649977179
transform 1 0 32016 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1649977179
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1649977179
transform 1 0 37168 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1649977179
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1649977179
transform 1 0 42320 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1649977179
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1649977179
transform 1 0 47472 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1649977179
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1649977179
transform 1 0 52624 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _0727_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 23920 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0728_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22080 0 -1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0729_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 23276 0 1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0730_
timestamp 1649977179
transform 1 0 25300 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0731_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 27232 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0732_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 23092 0 -1 47872
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0733_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 23460 0 -1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0734_
timestamp 1649977179
transform 1 0 22448 0 1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0735_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22632 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0736_
timestamp 1649977179
transform -1 0 22816 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0737_
timestamp 1649977179
transform 1 0 23276 0 1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0738_
timestamp 1649977179
transform 1 0 24840 0 -1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0739_
timestamp 1649977179
transform 1 0 25668 0 1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__buf_8  _0740_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 35788 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_2  _0741_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 30268 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_8  _0742_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 33580 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_1  _0743_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 25116 0 -1 47872
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0744_
timestamp 1649977179
transform -1 0 24748 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0745_
timestamp 1649977179
transform 1 0 23000 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0746_
timestamp 1649977179
transform -1 0 24564 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0747_
timestamp 1649977179
transform 1 0 23368 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0748_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 24932 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0749_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 27140 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _0750_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 39192 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0751_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 31188 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_8  _0752_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 33396 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__a31o_1  _0753_
timestamp 1649977179
transform 1 0 25484 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  _0754_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 29532 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _0755_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 31648 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_8  _0756_
timestamp 1649977179
transform 1 0 27784 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  _0757_
timestamp 1649977179
transform -1 0 25760 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0758_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 35512 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _0759_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 25668 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0760_
timestamp 1649977179
transform -1 0 27508 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_8  _0761_
timestamp 1649977179
transform 1 0 27600 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_1  _0762_
timestamp 1649977179
transform -1 0 24840 0 1 52224
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0763_
timestamp 1649977179
transform 1 0 23828 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0764_
timestamp 1649977179
transform -1 0 23920 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0765_
timestamp 1649977179
transform 1 0 23184 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0766_
timestamp 1649977179
transform 1 0 24564 0 -1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0767_
timestamp 1649977179
transform 1 0 25484 0 1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0768_
timestamp 1649977179
transform 1 0 25484 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0769_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 25852 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0770_
timestamp 1649977179
transform 1 0 26496 0 1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0771_
timestamp 1649977179
transform 1 0 32200 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _0772_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 32936 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0773_
timestamp 1649977179
transform 1 0 26588 0 1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0774_
timestamp 1649977179
transform 1 0 25944 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0775_
timestamp 1649977179
transform 1 0 26220 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 25576 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0777_
timestamp 1649977179
transform -1 0 26496 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0778_
timestamp 1649977179
transform 1 0 26128 0 1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0779_
timestamp 1649977179
transform 1 0 26956 0 -1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__inv_4  _0780_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 31648 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0781_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 27876 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0782_
timestamp 1649977179
transform -1 0 27692 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0783_
timestamp 1649977179
transform -1 0 32752 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0784_
timestamp 1649977179
transform 1 0 32384 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0785_
timestamp 1649977179
transform -1 0 33488 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0786_
timestamp 1649977179
transform -1 0 23920 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_2  _0787_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 24196 0 -1 52224
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0788_
timestamp 1649977179
transform -1 0 30176 0 1 53312
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0789_
timestamp 1649977179
transform 1 0 29440 0 -1 52224
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0790_
timestamp 1649977179
transform -1 0 29624 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0791_
timestamp 1649977179
transform -1 0 29072 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0792_
timestamp 1649977179
transform 1 0 26036 0 -1 52224
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0793_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 28060 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0794_
timestamp 1649977179
transform 1 0 27692 0 -1 53312
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0795_
timestamp 1649977179
transform -1 0 30912 0 1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0796_
timestamp 1649977179
transform -1 0 31556 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0797_
timestamp 1649977179
transform -1 0 29072 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_2  _0798_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 27876 0 -1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0799_
timestamp 1649977179
transform 1 0 27968 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0800_
timestamp 1649977179
transform 1 0 28336 0 -1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0801_
timestamp 1649977179
transform 1 0 29532 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0802_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 28796 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0803_
timestamp 1649977179
transform -1 0 29072 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0804_
timestamp 1649977179
transform -1 0 29716 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0805_
timestamp 1649977179
transform -1 0 29072 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0806_
timestamp 1649977179
transform 1 0 30544 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0807_
timestamp 1649977179
transform 1 0 30636 0 1 52224
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0808_
timestamp 1649977179
transform -1 0 31924 0 1 52224
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0809_
timestamp 1649977179
transform -1 0 31556 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0810_
timestamp 1649977179
transform -1 0 31464 0 -1 53312
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0811_
timestamp 1649977179
transform -1 0 30912 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0812_
timestamp 1649977179
transform 1 0 30728 0 -1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0813_
timestamp 1649977179
transform 1 0 31280 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0814_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 29532 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0815_
timestamp 1649977179
transform 1 0 29992 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0816_
timestamp 1649977179
transform 1 0 29900 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_2  _0817_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 28244 0 1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0818_
timestamp 1649977179
transform -1 0 32384 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0819_
timestamp 1649977179
transform -1 0 31188 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0820_
timestamp 1649977179
transform 1 0 30820 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0821_
timestamp 1649977179
transform 1 0 30728 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0822_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 30452 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0823_
timestamp 1649977179
transform -1 0 40020 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0824_
timestamp 1649977179
transform -1 0 32568 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _0825_
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _0826_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 29624 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0827_
timestamp 1649977179
transform 1 0 30636 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0828_
timestamp 1649977179
transform -1 0 30360 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0829_
timestamp 1649977179
transform 1 0 29716 0 1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0830_
timestamp 1649977179
transform 1 0 29532 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0831_
timestamp 1649977179
transform -1 0 31464 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _0832_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 33028 0 1 52224
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_1  _0833_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 32108 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0834_
timestamp 1649977179
transform -1 0 34868 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0835_
timestamp 1649977179
transform -1 0 32660 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0836_
timestamp 1649977179
transform -1 0 35328 0 1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0837_
timestamp 1649977179
transform -1 0 34684 0 -1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1649977179
transform -1 0 34224 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0839_
timestamp 1649977179
transform -1 0 33580 0 1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0840_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 32752 0 1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0841_
timestamp 1649977179
transform -1 0 32476 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0842_
timestamp 1649977179
transform -1 0 35696 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0843_
timestamp 1649977179
transform 1 0 33488 0 -1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0844_
timestamp 1649977179
transform 1 0 35144 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0845_
timestamp 1649977179
transform 1 0 30544 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0846_
timestamp 1649977179
transform -1 0 32752 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0847_
timestamp 1649977179
transform -1 0 33764 0 1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0848_
timestamp 1649977179
transform 1 0 32108 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0849_
timestamp 1649977179
transform -1 0 33672 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _0850_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 32292 0 1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0851_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 31740 0 1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0852_
timestamp 1649977179
transform -1 0 35144 0 -1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0853_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 33948 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0854_
timestamp 1649977179
transform 1 0 34316 0 -1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0855_
timestamp 1649977179
transform 1 0 35604 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0856_
timestamp 1649977179
transform 1 0 34592 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0857_
timestamp 1649977179
transform -1 0 35880 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0858_
timestamp 1649977179
transform -1 0 35236 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0859_
timestamp 1649977179
transform 1 0 33856 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0860_
timestamp 1649977179
transform 1 0 33396 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0861_
timestamp 1649977179
transform -1 0 35144 0 1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0862_
timestamp 1649977179
transform -1 0 35788 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0863_
timestamp 1649977179
transform -1 0 35328 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0864_
timestamp 1649977179
transform 1 0 34684 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0865_
timestamp 1649977179
transform -1 0 34776 0 -1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0866_
timestamp 1649977179
transform -1 0 32568 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0867_
timestamp 1649977179
transform 1 0 32108 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0868_
timestamp 1649977179
transform -1 0 33396 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0869_
timestamp 1649977179
transform 1 0 32200 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0870_
timestamp 1649977179
transform 1 0 33120 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0871_
timestamp 1649977179
transform 1 0 33212 0 1 53312
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0872_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 34684 0 1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0873_
timestamp 1649977179
transform 1 0 35328 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _0874_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 33212 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _0875_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 33212 0 1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0876_
timestamp 1649977179
transform -1 0 35604 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0877_
timestamp 1649977179
transform -1 0 36432 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0878_
timestamp 1649977179
transform -1 0 35788 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0879_
timestamp 1649977179
transform 1 0 35788 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0880_
timestamp 1649977179
transform 1 0 36616 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0881_
timestamp 1649977179
transform -1 0 36616 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0882_
timestamp 1649977179
transform -1 0 35788 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0883_
timestamp 1649977179
transform 1 0 34132 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0884_
timestamp 1649977179
transform 1 0 34684 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0885_
timestamp 1649977179
transform -1 0 34960 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0886_
timestamp 1649977179
transform -1 0 33120 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0887_
timestamp 1649977179
transform 1 0 32016 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0888_
timestamp 1649977179
transform -1 0 34684 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _0889_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 33120 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__o41a_1  _0890_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 33764 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0891_
timestamp 1649977179
transform 1 0 32476 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0892_
timestamp 1649977179
transform -1 0 33856 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0893_
timestamp 1649977179
transform 1 0 32568 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0894_
timestamp 1649977179
transform -1 0 32384 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0895_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 32752 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0896_
timestamp 1649977179
transform 1 0 33212 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0897_
timestamp 1649977179
transform 1 0 36800 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0898_
timestamp 1649977179
transform 1 0 38916 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0899_
timestamp 1649977179
transform -1 0 37904 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0900_
timestamp 1649977179
transform -1 0 36524 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0901_
timestamp 1649977179
transform -1 0 36708 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0902_
timestamp 1649977179
transform -1 0 36616 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0903_
timestamp 1649977179
transform -1 0 36432 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0904_
timestamp 1649977179
transform -1 0 35788 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _0905_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 36248 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _0906_
timestamp 1649977179
transform -1 0 35052 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0907_
timestamp 1649977179
transform 1 0 35420 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0908_
timestamp 1649977179
transform -1 0 34684 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0909_
timestamp 1649977179
transform 1 0 34684 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0910_
timestamp 1649977179
transform -1 0 34684 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0911_
timestamp 1649977179
transform 1 0 34684 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0912_
timestamp 1649977179
transform 1 0 34224 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0913_
timestamp 1649977179
transform -1 0 35604 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0914_
timestamp 1649977179
transform -1 0 33856 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0915_
timestamp 1649977179
transform 1 0 32936 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0916_
timestamp 1649977179
transform 1 0 33120 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0917_
timestamp 1649977179
transform -1 0 33764 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0918_
timestamp 1649977179
transform -1 0 32660 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0919_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 32384 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0920_
timestamp 1649977179
transform 1 0 34132 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0921_
timestamp 1649977179
transform -1 0 34960 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0922_
timestamp 1649977179
transform 1 0 34960 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0923_
timestamp 1649977179
transform -1 0 35420 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0924_
timestamp 1649977179
transform -1 0 34132 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0925_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 34592 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0926_
timestamp 1649977179
transform -1 0 34224 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0927_
timestamp 1649977179
transform 1 0 33304 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0928_
timestamp 1649977179
transform 1 0 33948 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0929_
timestamp 1649977179
transform -1 0 33580 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0930_
timestamp 1649977179
transform -1 0 33396 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0931_
timestamp 1649977179
transform 1 0 33028 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0932_
timestamp 1649977179
transform -1 0 35604 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0933_
timestamp 1649977179
transform 1 0 35880 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0934_
timestamp 1649977179
transform -1 0 37812 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0935_
timestamp 1649977179
transform -1 0 39100 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0936_
timestamp 1649977179
transform 1 0 39836 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0937_
timestamp 1649977179
transform -1 0 37720 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0938_
timestamp 1649977179
transform -1 0 38548 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0939_
timestamp 1649977179
transform -1 0 38456 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0940_
timestamp 1649977179
transform 1 0 37260 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0941_
timestamp 1649977179
transform 1 0 36432 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0942_
timestamp 1649977179
transform -1 0 37720 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0943_
timestamp 1649977179
transform 1 0 36064 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0944_
timestamp 1649977179
transform -1 0 35236 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0945_
timestamp 1649977179
transform -1 0 35052 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0946_
timestamp 1649977179
transform -1 0 34500 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _0947_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 32936 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0948_
timestamp 1649977179
transform 1 0 34684 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_2  _0949_
timestamp 1649977179
transform -1 0 39376 0 1 40256
box -38 -48 1234 592
use sky130_fd_sc_hd__a22oi_2  _0950_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 38088 0 -1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_2  _0951_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 38180 0 1 39168
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0952_
timestamp 1649977179
transform -1 0 38824 0 -1 36992
box -38 -48 1234 592
use sky130_fd_sc_hd__o21bai_1  _0953_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 36984 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _0954_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 36064 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0955_
timestamp 1649977179
transform -1 0 36800 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0956_
timestamp 1649977179
transform 1 0 32384 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0957_
timestamp 1649977179
transform -1 0 37904 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0958_
timestamp 1649977179
transform 1 0 37352 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0959_
timestamp 1649977179
transform -1 0 38364 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0960_
timestamp 1649977179
transform 1 0 35420 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0961_
timestamp 1649977179
transform -1 0 34408 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0962_
timestamp 1649977179
transform -1 0 35052 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0963_
timestamp 1649977179
transform -1 0 34224 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0964_
timestamp 1649977179
transform -1 0 36892 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0965_
timestamp 1649977179
transform 1 0 35788 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0966_
timestamp 1649977179
transform -1 0 37720 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0967_
timestamp 1649977179
transform -1 0 37720 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0968_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 37720 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0969_
timestamp 1649977179
transform 1 0 39376 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0970_
timestamp 1649977179
transform 1 0 38824 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0971_
timestamp 1649977179
transform 1 0 36248 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0972_
timestamp 1649977179
transform 1 0 37260 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0973_
timestamp 1649977179
transform 1 0 38732 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0974_
timestamp 1649977179
transform 1 0 38732 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0975_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 37996 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _0976_
timestamp 1649977179
transform 1 0 38088 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0977_
timestamp 1649977179
transform -1 0 38364 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0978_
timestamp 1649977179
transform -1 0 37260 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0979_
timestamp 1649977179
transform -1 0 35696 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0980_
timestamp 1649977179
transform -1 0 35512 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0981_
timestamp 1649977179
transform 1 0 35144 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0982_
timestamp 1649977179
transform -1 0 37720 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0983_
timestamp 1649977179
transform -1 0 36800 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0984_
timestamp 1649977179
transform 1 0 34776 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0985_
timestamp 1649977179
transform -1 0 34776 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0986_
timestamp 1649977179
transform -1 0 33028 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0987_
timestamp 1649977179
transform -1 0 33672 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0988_
timestamp 1649977179
transform -1 0 32936 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0989_
timestamp 1649977179
transform 1 0 32108 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0990_
timestamp 1649977179
transform -1 0 31648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0991_
timestamp 1649977179
transform -1 0 30912 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0992_
timestamp 1649977179
transform -1 0 32844 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0993_
timestamp 1649977179
transform 1 0 35512 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0994_
timestamp 1649977179
transform 1 0 35052 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0995_
timestamp 1649977179
transform -1 0 36432 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0996_
timestamp 1649977179
transform -1 0 37996 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0997_
timestamp 1649977179
transform -1 0 36524 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0998_
timestamp 1649977179
transform -1 0 33396 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0999_
timestamp 1649977179
transform -1 0 33120 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1000_
timestamp 1649977179
transform 1 0 33028 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1001_
timestamp 1649977179
transform 1 0 36340 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1002_
timestamp 1649977179
transform -1 0 35512 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _1003_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 39192 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1004_
timestamp 1649977179
transform 1 0 36984 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _1005_
timestamp 1649977179
transform -1 0 32660 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1006_
timestamp 1649977179
transform -1 0 32660 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1007_
timestamp 1649977179
transform -1 0 32476 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1008_
timestamp 1649977179
transform -1 0 31372 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1009_
timestamp 1649977179
transform 1 0 31280 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1010_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 31188 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1011_
timestamp 1649977179
transform -1 0 36340 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1012_
timestamp 1649977179
transform 1 0 35604 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1013_
timestamp 1649977179
transform 1 0 35788 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1014_
timestamp 1649977179
transform 1 0 33672 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1015_
timestamp 1649977179
transform -1 0 34684 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1016_
timestamp 1649977179
transform 1 0 30176 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1017_
timestamp 1649977179
transform -1 0 29624 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1018_
timestamp 1649977179
transform 1 0 33948 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1019_
timestamp 1649977179
transform 1 0 36248 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1020_
timestamp 1649977179
transform 1 0 37260 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1021_
timestamp 1649977179
transform 1 0 36156 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _1022_
timestamp 1649977179
transform -1 0 35880 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1023_
timestamp 1649977179
transform -1 0 33948 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1024_
timestamp 1649977179
transform 1 0 31924 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1025_
timestamp 1649977179
transform 1 0 31280 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1026_
timestamp 1649977179
transform -1 0 29072 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1027_
timestamp 1649977179
transform 1 0 28520 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1028_
timestamp 1649977179
transform -1 0 31556 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1029_
timestamp 1649977179
transform -1 0 36156 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1030_
timestamp 1649977179
transform -1 0 35420 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1031_
timestamp 1649977179
transform 1 0 34684 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1032_
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1033_
timestamp 1649977179
transform 1 0 30452 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1034_
timestamp 1649977179
transform -1 0 29808 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1035_
timestamp 1649977179
transform 1 0 30084 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1036_
timestamp 1649977179
transform 1 0 30176 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _1037_
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1038_
timestamp 1649977179
transform 1 0 28336 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1039_
timestamp 1649977179
transform 1 0 27600 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1040_
timestamp 1649977179
transform 1 0 29624 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1041_
timestamp 1649977179
transform -1 0 31832 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1042_
timestamp 1649977179
transform 1 0 30820 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1043_
timestamp 1649977179
transform -1 0 35788 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1044_
timestamp 1649977179
transform -1 0 36248 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1045_
timestamp 1649977179
transform 1 0 33580 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1046_
timestamp 1649977179
transform -1 0 36432 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1047_
timestamp 1649977179
transform -1 0 36524 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1048_
timestamp 1649977179
transform -1 0 35420 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _1049_
timestamp 1649977179
transform -1 0 31004 0 -1 38080
box -38 -48 1234 592
use sky130_fd_sc_hd__nor3_1  _1050_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 32844 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1051_
timestamp 1649977179
transform 1 0 33764 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1052_
timestamp 1649977179
transform 1 0 33672 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1053_
timestamp 1649977179
transform 1 0 30820 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1054_
timestamp 1649977179
transform 1 0 29624 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1055_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 29532 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1056_
timestamp 1649977179
transform 1 0 30544 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1057_
timestamp 1649977179
transform -1 0 28612 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1058_
timestamp 1649977179
transform 1 0 34960 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_1  _1059_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 35972 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1060_
timestamp 1649977179
transform 1 0 35420 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_4  _1061_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 37628 0 1 40256
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_1  _1062_
timestamp 1649977179
transform -1 0 34224 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1063_
timestamp 1649977179
transform -1 0 36800 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_2  _1064_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 35420 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1065_
timestamp 1649977179
transform 1 0 16100 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1066_
timestamp 1649977179
transform 1 0 17664 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1067_
timestamp 1649977179
transform -1 0 17756 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1068_
timestamp 1649977179
transform 1 0 17572 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1069_
timestamp 1649977179
transform 1 0 17664 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1070_
timestamp 1649977179
transform 1 0 18400 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1071_
timestamp 1649977179
transform -1 0 31004 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1072_
timestamp 1649977179
transform 1 0 32200 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1073_
timestamp 1649977179
transform -1 0 31188 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1074_
timestamp 1649977179
transform -1 0 32200 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1075_
timestamp 1649977179
transform -1 0 29072 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1076_
timestamp 1649977179
transform 1 0 29900 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1077_
timestamp 1649977179
transform 1 0 29532 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1078_
timestamp 1649977179
transform 1 0 30728 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1079_
timestamp 1649977179
transform 1 0 24380 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1080_
timestamp 1649977179
transform 1 0 24380 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1081_
timestamp 1649977179
transform -1 0 25484 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1082_
timestamp 1649977179
transform 1 0 29348 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1083_
timestamp 1649977179
transform 1 0 29624 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1084_
timestamp 1649977179
transform 1 0 28612 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1085_
timestamp 1649977179
transform 1 0 25024 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1086_
timestamp 1649977179
transform 1 0 24656 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1087_
timestamp 1649977179
transform 1 0 25484 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1088_
timestamp 1649977179
transform 1 0 29532 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1089_
timestamp 1649977179
transform 1 0 22540 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1090_
timestamp 1649977179
transform -1 0 22908 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1091_
timestamp 1649977179
transform 1 0 23276 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1092_
timestamp 1649977179
transform 1 0 25392 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1093_
timestamp 1649977179
transform 1 0 25392 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1094_
timestamp 1649977179
transform -1 0 25576 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1095_
timestamp 1649977179
transform -1 0 18124 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1096_
timestamp 1649977179
transform -1 0 16928 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1097_
timestamp 1649977179
transform 1 0 17296 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _1098_
timestamp 1649977179
transform -1 0 18860 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1099_
timestamp 1649977179
transform -1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1100_
timestamp 1649977179
transform 1 0 19136 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1101_
timestamp 1649977179
transform -1 0 18768 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1102_
timestamp 1649977179
transform 1 0 19320 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1103_
timestamp 1649977179
transform -1 0 31832 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1104_
timestamp 1649977179
transform -1 0 31372 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1105_
timestamp 1649977179
transform -1 0 29992 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1106_
timestamp 1649977179
transform -1 0 29900 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1107_
timestamp 1649977179
transform -1 0 31004 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _1108_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 30360 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1109_
timestamp 1649977179
transform 1 0 20884 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1110_
timestamp 1649977179
transform -1 0 20976 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1111_
timestamp 1649977179
transform 1 0 21804 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1112_
timestamp 1649977179
transform -1 0 31464 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1113_
timestamp 1649977179
transform 1 0 29532 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1114_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 29072 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1115_
timestamp 1649977179
transform -1 0 26588 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1116_
timestamp 1649977179
transform 1 0 27692 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1117_
timestamp 1649977179
transform 1 0 30820 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1118_
timestamp 1649977179
transform 1 0 21896 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1119_
timestamp 1649977179
transform 1 0 22356 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1120_
timestamp 1649977179
transform 1 0 22908 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1121_
timestamp 1649977179
transform 1 0 23552 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1122_
timestamp 1649977179
transform 1 0 25116 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1123_
timestamp 1649977179
transform 1 0 23276 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1124_
timestamp 1649977179
transform 1 0 14720 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1125_
timestamp 1649977179
transform 1 0 14720 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1126_
timestamp 1649977179
transform 1 0 15548 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1127_
timestamp 1649977179
transform -1 0 15732 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1128_
timestamp 1649977179
transform -1 0 17296 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1129_
timestamp 1649977179
transform 1 0 16928 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1130_
timestamp 1649977179
transform 1 0 19780 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1131_
timestamp 1649977179
transform 1 0 20148 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1132_
timestamp 1649977179
transform 1 0 20056 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1133_
timestamp 1649977179
transform 1 0 21160 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1134_
timestamp 1649977179
transform 1 0 20608 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1135_
timestamp 1649977179
transform -1 0 25024 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1136_
timestamp 1649977179
transform -1 0 29072 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1137_
timestamp 1649977179
transform 1 0 21896 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1138_
timestamp 1649977179
transform 1 0 22540 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1139_
timestamp 1649977179
transform 1 0 23184 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1140_
timestamp 1649977179
transform 1 0 23552 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1141_
timestamp 1649977179
transform 1 0 24104 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1142_
timestamp 1649977179
transform 1 0 26036 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1143_
timestamp 1649977179
transform -1 0 28244 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1144_
timestamp 1649977179
transform 1 0 28612 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1145_
timestamp 1649977179
transform 1 0 16652 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1146_
timestamp 1649977179
transform 1 0 14076 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1147_
timestamp 1649977179
transform 1 0 14076 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1148_
timestamp 1649977179
transform 1 0 14720 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1149_
timestamp 1649977179
transform 1 0 15824 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1150_
timestamp 1649977179
transform -1 0 16284 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1151_
timestamp 1649977179
transform -1 0 19964 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1152_
timestamp 1649977179
transform -1 0 19872 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1153_
timestamp 1649977179
transform 1 0 19412 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1154_
timestamp 1649977179
transform -1 0 20332 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1155_
timestamp 1649977179
transform 1 0 20424 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1156_
timestamp 1649977179
transform 1 0 20792 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1157_
timestamp 1649977179
transform -1 0 27784 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1158_
timestamp 1649977179
transform 1 0 26956 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1159_
timestamp 1649977179
transform 1 0 16652 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1160_
timestamp 1649977179
transform 1 0 17664 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1161_
timestamp 1649977179
transform 1 0 17480 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1162_
timestamp 1649977179
transform 1 0 14904 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1163_
timestamp 1649977179
transform -1 0 17296 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1164_
timestamp 1649977179
transform 1 0 16284 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1165_
timestamp 1649977179
transform 1 0 15916 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1166_
timestamp 1649977179
transform 1 0 15916 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1167_
timestamp 1649977179
transform 1 0 17020 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1168_
timestamp 1649977179
transform 1 0 16560 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1169_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17848 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _1170_
timestamp 1649977179
transform 1 0 19596 0 -1 41344
box -38 -48 1234 592
use sky130_fd_sc_hd__a21boi_1  _1171_
timestamp 1649977179
transform 1 0 19872 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1172_
timestamp 1649977179
transform 1 0 21620 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1173_
timestamp 1649977179
transform -1 0 27416 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1174_
timestamp 1649977179
transform 1 0 27232 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1175_
timestamp 1649977179
transform 1 0 27784 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1176_
timestamp 1649977179
transform 1 0 26772 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1177_
timestamp 1649977179
transform -1 0 22816 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1178_
timestamp 1649977179
transform -1 0 23368 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1179_
timestamp 1649977179
transform 1 0 22172 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1180_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 24472 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1181_
timestamp 1649977179
transform -1 0 23184 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1182_
timestamp 1649977179
transform -1 0 23920 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1183_
timestamp 1649977179
transform -1 0 24104 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1184_
timestamp 1649977179
transform -1 0 24656 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1185_
timestamp 1649977179
transform 1 0 24380 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1186_
timestamp 1649977179
transform 1 0 26220 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1187_
timestamp 1649977179
transform -1 0 27416 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1188_
timestamp 1649977179
transform 1 0 26956 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1189_
timestamp 1649977179
transform 1 0 23460 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1190_
timestamp 1649977179
transform -1 0 23092 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1191_
timestamp 1649977179
transform 1 0 22816 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1192_
timestamp 1649977179
transform 1 0 25484 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1193_
timestamp 1649977179
transform 1 0 23736 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1194_
timestamp 1649977179
transform -1 0 19872 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1195_
timestamp 1649977179
transform -1 0 19228 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1196_
timestamp 1649977179
transform -1 0 18676 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1197_
timestamp 1649977179
transform -1 0 18768 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1198_
timestamp 1649977179
transform -1 0 18032 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1199_
timestamp 1649977179
transform 1 0 19780 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1200_
timestamp 1649977179
transform -1 0 20056 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1201_
timestamp 1649977179
transform -1 0 20700 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1202_
timestamp 1649977179
transform 1 0 21804 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1203_
timestamp 1649977179
transform 1 0 20792 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1204_
timestamp 1649977179
transform 1 0 21620 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1205_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20240 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1206_
timestamp 1649977179
transform -1 0 20976 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a311oi_2  _1207_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21252 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__a21bo_1  _1208_
timestamp 1649977179
transform 1 0 20608 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1209_
timestamp 1649977179
transform 1 0 21804 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1210_
timestamp 1649977179
transform -1 0 23920 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1211_
timestamp 1649977179
transform -1 0 26588 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1212_
timestamp 1649977179
transform -1 0 23644 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1213_
timestamp 1649977179
transform 1 0 22816 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1214_
timestamp 1649977179
transform -1 0 24564 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1215_
timestamp 1649977179
transform 1 0 23644 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1216_
timestamp 1649977179
transform -1 0 24288 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1217_
timestamp 1649977179
transform -1 0 25484 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1218_
timestamp 1649977179
transform 1 0 24380 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1219_
timestamp 1649977179
transform 1 0 26680 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1220_
timestamp 1649977179
transform 1 0 26680 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1221_
timestamp 1649977179
transform -1 0 17112 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1222_
timestamp 1649977179
transform -1 0 17756 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1223_
timestamp 1649977179
transform -1 0 18216 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1224_
timestamp 1649977179
transform -1 0 19504 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1225_
timestamp 1649977179
transform -1 0 19688 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1226_
timestamp 1649977179
transform -1 0 18400 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1227_
timestamp 1649977179
transform -1 0 17940 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1228_
timestamp 1649977179
transform -1 0 17756 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1229_
timestamp 1649977179
transform 1 0 18400 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1230_
timestamp 1649977179
transform -1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1231_
timestamp 1649977179
transform -1 0 20332 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1232_
timestamp 1649977179
transform 1 0 19964 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1233_
timestamp 1649977179
transform -1 0 22172 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1234_
timestamp 1649977179
transform -1 0 21436 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _1235_
timestamp 1649977179
transform -1 0 26496 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _1236_
timestamp 1649977179
transform 1 0 25116 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1237_
timestamp 1649977179
transform 1 0 26036 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1238_
timestamp 1649977179
transform -1 0 23920 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1239_
timestamp 1649977179
transform -1 0 23920 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1240_
timestamp 1649977179
transform 1 0 23000 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1241_
timestamp 1649977179
transform 1 0 25484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1242_
timestamp 1649977179
transform -1 0 24932 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1243_
timestamp 1649977179
transform -1 0 24840 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1244_
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1245_
timestamp 1649977179
transform 1 0 26956 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1246_
timestamp 1649977179
transform -1 0 19320 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1247_
timestamp 1649977179
transform 1 0 16836 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1248_
timestamp 1649977179
transform 1 0 17388 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1249_
timestamp 1649977179
transform -1 0 18676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1250_
timestamp 1649977179
transform 1 0 19228 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1251_
timestamp 1649977179
transform 1 0 19780 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1252_
timestamp 1649977179
transform 1 0 19044 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1253_
timestamp 1649977179
transform 1 0 22080 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1254_
timestamp 1649977179
transform -1 0 23092 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _1255_
timestamp 1649977179
transform 1 0 19688 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1256_
timestamp 1649977179
transform 1 0 20608 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1257_
timestamp 1649977179
transform 1 0 21804 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1258_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 26404 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1259_
timestamp 1649977179
transform -1 0 25944 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1260_
timestamp 1649977179
transform -1 0 21712 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1261_
timestamp 1649977179
transform -1 0 18584 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1262_
timestamp 1649977179
transform 1 0 17572 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _1263_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17940 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1264_
timestamp 1649977179
transform -1 0 18492 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1265_
timestamp 1649977179
transform -1 0 18216 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1266_
timestamp 1649977179
transform -1 0 18400 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _1267_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17480 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1268_
timestamp 1649977179
transform 1 0 17204 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1269_
timestamp 1649977179
transform 1 0 18492 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1270_
timestamp 1649977179
transform 1 0 19688 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1271_
timestamp 1649977179
transform 1 0 21712 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1272_
timestamp 1649977179
transform 1 0 20976 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1273_
timestamp 1649977179
transform 1 0 22172 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1274_
timestamp 1649977179
transform 1 0 21988 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1275_
timestamp 1649977179
transform -1 0 22908 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1276_
timestamp 1649977179
transform -1 0 25116 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1277_
timestamp 1649977179
transform -1 0 23920 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1278_
timestamp 1649977179
transform 1 0 24380 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1279_
timestamp 1649977179
transform 1 0 24380 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _1280_
timestamp 1649977179
transform 1 0 24472 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1281_
timestamp 1649977179
transform 1 0 23920 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1282_
timestamp 1649977179
transform 1 0 23276 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1283_
timestamp 1649977179
transform 1 0 25024 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1284_
timestamp 1649977179
transform -1 0 25852 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _1285_
timestamp 1649977179
transform 1 0 22540 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1286_
timestamp 1649977179
transform 1 0 26864 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1287_
timestamp 1649977179
transform -1 0 26496 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1288_
timestamp 1649977179
transform -1 0 27232 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1289_
timestamp 1649977179
transform -1 0 21068 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  _1290_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21804 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1291_
timestamp 1649977179
transform 1 0 20792 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1292_
timestamp 1649977179
transform 1 0 20424 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1293_
timestamp 1649977179
transform -1 0 20148 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1294_
timestamp 1649977179
transform 1 0 19780 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1295_
timestamp 1649977179
transform -1 0 21344 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1296_
timestamp 1649977179
transform -1 0 21344 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1297_
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1298_
timestamp 1649977179
transform -1 0 19688 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1299_
timestamp 1649977179
transform -1 0 17848 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1300_
timestamp 1649977179
transform -1 0 18584 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1301_
timestamp 1649977179
transform 1 0 17388 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1302_
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1303_
timestamp 1649977179
transform 1 0 18952 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1304_
timestamp 1649977179
transform -1 0 20148 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1305_
timestamp 1649977179
transform 1 0 20056 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1306_
timestamp 1649977179
transform 1 0 20608 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1307_
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1308_
timestamp 1649977179
transform 1 0 23092 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1309_
timestamp 1649977179
transform 1 0 21896 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1310_
timestamp 1649977179
transform 1 0 21896 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1311_
timestamp 1649977179
transform 1 0 22448 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1312_
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1313_
timestamp 1649977179
transform 1 0 25484 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1314_
timestamp 1649977179
transform -1 0 26128 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1315_
timestamp 1649977179
transform 1 0 22540 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1316_
timestamp 1649977179
transform -1 0 21804 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1317_
timestamp 1649977179
transform 1 0 21252 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1318_
timestamp 1649977179
transform 1 0 22080 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1319_
timestamp 1649977179
transform -1 0 23552 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1320_
timestamp 1649977179
transform -1 0 22908 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _1321_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 24380 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1322_
timestamp 1649977179
transform -1 0 17664 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1323_
timestamp 1649977179
transform -1 0 16836 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1324_
timestamp 1649977179
transform 1 0 16928 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1325_
timestamp 1649977179
transform 1 0 18032 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1326_
timestamp 1649977179
transform 1 0 18032 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1327_
timestamp 1649977179
transform 1 0 18032 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1328_
timestamp 1649977179
transform 1 0 19320 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1329_
timestamp 1649977179
transform 1 0 20240 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1330_
timestamp 1649977179
transform 1 0 20332 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1331_
timestamp 1649977179
transform -1 0 26128 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1332_
timestamp 1649977179
transform -1 0 26220 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1333_
timestamp 1649977179
transform -1 0 26036 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1334_
timestamp 1649977179
transform 1 0 25576 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1335_
timestamp 1649977179
transform -1 0 23736 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1336_
timestamp 1649977179
transform -1 0 23184 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1337_
timestamp 1649977179
transform 1 0 24472 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1338_
timestamp 1649977179
transform 1 0 23552 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1339_
timestamp 1649977179
transform -1 0 22172 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1340_
timestamp 1649977179
transform -1 0 25024 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1341_
timestamp 1649977179
transform -1 0 24472 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1342_
timestamp 1649977179
transform -1 0 18952 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1343_
timestamp 1649977179
transform -1 0 19412 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1344_
timestamp 1649977179
transform -1 0 20148 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1345_
timestamp 1649977179
transform -1 0 19872 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1346_
timestamp 1649977179
transform 1 0 18400 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1347_
timestamp 1649977179
transform 1 0 19504 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1348_
timestamp 1649977179
transform 1 0 20516 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1349_
timestamp 1649977179
transform -1 0 20976 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1350_
timestamp 1649977179
transform -1 0 20884 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1351_
timestamp 1649977179
transform 1 0 20792 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1352_
timestamp 1649977179
transform 1 0 22080 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1353_
timestamp 1649977179
transform -1 0 20424 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1354_
timestamp 1649977179
transform -1 0 21160 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _1355_
timestamp 1649977179
transform 1 0 21160 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1356_
timestamp 1649977179
transform -1 0 23092 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1357_
timestamp 1649977179
transform 1 0 23000 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1358_
timestamp 1649977179
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1359_
timestamp 1649977179
transform 1 0 25116 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _1360_
timestamp 1649977179
transform 1 0 24840 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1361_
timestamp 1649977179
transform 1 0 20608 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1362_
timestamp 1649977179
transform -1 0 20332 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1363_
timestamp 1649977179
transform 1 0 19964 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1364_
timestamp 1649977179
transform -1 0 20240 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1365_
timestamp 1649977179
transform 1 0 19320 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1366_
timestamp 1649977179
transform 1 0 19872 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1367_
timestamp 1649977179
transform 1 0 21160 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1368_
timestamp 1649977179
transform -1 0 22816 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1369_
timestamp 1649977179
transform 1 0 23184 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1370_
timestamp 1649977179
transform -1 0 23460 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1371_
timestamp 1649977179
transform -1 0 23552 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1372_
timestamp 1649977179
transform 1 0 24196 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1373_
timestamp 1649977179
transform 1 0 22908 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1374_
timestamp 1649977179
transform 1 0 23184 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _1375_
timestamp 1649977179
transform -1 0 24104 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1376_
timestamp 1649977179
transform -1 0 25116 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1377_
timestamp 1649977179
transform 1 0 24012 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1378_
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1379_
timestamp 1649977179
transform -1 0 24472 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1380_
timestamp 1649977179
transform 1 0 25116 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1381_
timestamp 1649977179
transform -1 0 25392 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1382_
timestamp 1649977179
transform 1 0 25760 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1383_
timestamp 1649977179
transform -1 0 25944 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1384_
timestamp 1649977179
transform 1 0 24840 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1385_
timestamp 1649977179
transform -1 0 24196 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1386_
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1387_
timestamp 1649977179
transform -1 0 27232 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1388_
timestamp 1649977179
transform 1 0 26312 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1389_
timestamp 1649977179
transform -1 0 27508 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1390_
timestamp 1649977179
transform 1 0 25944 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1391_
timestamp 1649977179
transform 1 0 25944 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _1392_
timestamp 1649977179
transform 1 0 25944 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1393_
timestamp 1649977179
transform 1 0 20608 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1394_
timestamp 1649977179
transform 1 0 20516 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1395_
timestamp 1649977179
transform -1 0 22080 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1396_
timestamp 1649977179
transform -1 0 20240 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1397_
timestamp 1649977179
transform 1 0 20608 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1398_
timestamp 1649977179
transform 1 0 21620 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1399_
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1400_
timestamp 1649977179
transform 1 0 20976 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1401_
timestamp 1649977179
transform 1 0 21252 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1402_
timestamp 1649977179
transform -1 0 22632 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _1403_
timestamp 1649977179
transform 1 0 22356 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1404_
timestamp 1649977179
transform -1 0 22724 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1405_
timestamp 1649977179
transform 1 0 24564 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1406_
timestamp 1649977179
transform -1 0 26772 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1407_
timestamp 1649977179
transform 1 0 24564 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _1408_
timestamp 1649977179
transform -1 0 25944 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1409_
timestamp 1649977179
transform -1 0 27324 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1410_
timestamp 1649977179
transform 1 0 22632 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1411_
timestamp 1649977179
transform -1 0 28336 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1412_
timestamp 1649977179
transform -1 0 31464 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1413_
timestamp 1649977179
transform -1 0 31280 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1414_
timestamp 1649977179
transform -1 0 31556 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1415_
timestamp 1649977179
transform 1 0 21344 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1416_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20700 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1417_
timestamp 1649977179
transform -1 0 30268 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1418_
timestamp 1649977179
transform 1 0 29808 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1419_
timestamp 1649977179
transform -1 0 29072 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1420_
timestamp 1649977179
transform 1 0 30820 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1421_
timestamp 1649977179
transform -1 0 28152 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1422_
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1423_
timestamp 1649977179
transform -1 0 28980 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1424_
timestamp 1649977179
transform 1 0 28796 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1425_
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1426_
timestamp 1649977179
transform -1 0 29992 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1427_
timestamp 1649977179
transform -1 0 28980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _1428_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 27692 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1429_
timestamp 1649977179
transform -1 0 27600 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1430_
timestamp 1649977179
transform -1 0 28244 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1431_
timestamp 1649977179
transform -1 0 29072 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1432_
timestamp 1649977179
transform 1 0 28244 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1433_
timestamp 1649977179
transform -1 0 34316 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1434_
timestamp 1649977179
transform 1 0 29164 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1435_
timestamp 1649977179
transform 1 0 30084 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1436_
timestamp 1649977179
transform 1 0 29900 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1437_
timestamp 1649977179
transform 1 0 30912 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1438_
timestamp 1649977179
transform -1 0 29072 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1439_
timestamp 1649977179
transform -1 0 30912 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1440_
timestamp 1649977179
transform 1 0 29992 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1441_
timestamp 1649977179
transform -1 0 31280 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1442_
timestamp 1649977179
transform 1 0 30360 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1443_
timestamp 1649977179
transform 1 0 30084 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1444_
timestamp 1649977179
transform 1 0 31096 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1445_
timestamp 1649977179
transform 1 0 31648 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1446_
timestamp 1649977179
transform 1 0 24840 0 1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1447_
timestamp 1649977179
transform 1 0 26036 0 -1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1448_
timestamp 1649977179
transform 1 0 24012 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1449_
timestamp 1649977179
transform 1 0 25392 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1450_
timestamp 1649977179
transform -1 0 26772 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1451_
timestamp 1649977179
transform -1 0 27232 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1452_
timestamp 1649977179
transform -1 0 25024 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1453_
timestamp 1649977179
transform -1 0 25392 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1454_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 28060 0 1 45696
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1455_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 27324 0 -1 52224
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1456_
timestamp 1649977179
transform 1 0 28704 0 -1 53312
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1457_
timestamp 1649977179
transform -1 0 30084 0 -1 50048
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1458_
timestamp 1649977179
transform 1 0 32108 0 -1 50048
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1459_
timestamp 1649977179
transform -1 0 32844 0 1 53312
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1460_
timestamp 1649977179
transform 1 0 31464 0 1 43520
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1461_
timestamp 1649977179
transform 1 0 32108 0 1 41344
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1462_
timestamp 1649977179
transform 1 0 32108 0 -1 39168
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1463_
timestamp 1649977179
transform -1 0 32016 0 1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1464_
timestamp 1649977179
transform 1 0 32384 0 1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1465_
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1466_
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1467_
timestamp 1649977179
transform -1 0 29072 0 1 35904
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1468_
timestamp 1649977179
transform -1 0 31004 0 -1 42432
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1469_
timestamp 1649977179
transform 1 0 26956 0 1 43520
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1470_
timestamp 1649977179
transform 1 0 29532 0 1 44608
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1471_
timestamp 1649977179
transform 1 0 29532 0 1 43520
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1472_
timestamp 1649977179
transform 1 0 26956 0 -1 41344
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1473_
timestamp 1649977179
transform 1 0 26956 0 1 39168
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1474_
timestamp 1649977179
transform 1 0 26956 0 -1 38080
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1475_
timestamp 1649977179
transform -1 0 26956 0 1 35904
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1476_
timestamp 1649977179
transform 1 0 26588 0 1 34816
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1477_
timestamp 1649977179
transform -1 0 28060 0 1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1478_
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1479_
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1480_
timestamp 1649977179
transform -1 0 27876 0 1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1481_
timestamp 1649977179
transform 1 0 26588 0 1 29376
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1482_
timestamp 1649977179
transform 1 0 28428 0 -1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1483_
timestamp 1649977179
transform -1 0 32568 0 1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1484_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 26864 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1485_
timestamp 1649977179
transform -1 0 28428 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 31740 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1649977179
transform -1 0 30452 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1649977179
transform -1 0 30452 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1649977179
transform -1 0 30452 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1649977179
transform 1 0 28612 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  input1 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 53728 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1649977179
transform -1 0 53728 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1649977179
transform -1 0 53728 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input4 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1748 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input5
timestamp 1649977179
transform 1 0 50508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 1649977179
transform 1 0 1380 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1649977179
transform 1 0 53360 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input8
timestamp 1649977179
transform 1 0 41308 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input9
timestamp 1649977179
transform 1 0 1748 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1649977179
transform 1 0 1748 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1649977179
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1649977179
transform 1 0 2668 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input13
timestamp 1649977179
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input14
timestamp 1649977179
transform 1 0 1380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1649977179
transform 1 0 1748 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1649977179
transform -1 0 53728 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1649977179
transform -1 0 25576 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input18
timestamp 1649977179
transform 1 0 47932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1649977179
transform 1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1649977179
transform 1 0 1748 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1649977179
transform 1 0 1748 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1649977179
transform 1 0 32292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1649977179
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input24
timestamp 1649977179
transform -1 0 53728 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input25
timestamp 1649977179
transform 1 0 1748 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1649977179
transform -1 0 53728 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1649977179
transform -1 0 35420 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19228 0 1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1649977179
transform -1 0 53728 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input30
timestamp 1649977179
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input31
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1649977179
transform -1 0 53728 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1649977179
transform 1 0 22172 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1649977179
transform -1 0 53728 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1649977179
transform -1 0 53728 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input36
timestamp 1649977179
transform 1 0 23276 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input37
timestamp 1649977179
transform 1 0 45172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1649977179
transform -1 0 53728 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1649977179
transform 1 0 7820 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1649977179
transform 1 0 1748 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1649977179
transform 1 0 27784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input42
timestamp 1649977179
transform 1 0 1748 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1649977179
transform 1 0 35052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1649977179
transform -1 0 11040 0 1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1649977179
transform 1 0 27784 0 1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1649977179
transform 1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp 1649977179
transform 1 0 1380 0 1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1649977179
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1649977179
transform -1 0 49404 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1649977179
transform -1 0 39100 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1649977179
transform -1 0 26220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input53
timestamp 1649977179
transform -1 0 53728 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input54
timestamp 1649977179
transform -1 0 53728 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1649977179
transform 1 0 1748 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1649977179
transform -1 0 53728 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1649977179
transform -1 0 11040 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1649977179
transform 1 0 19412 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input59
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1649977179
transform -1 0 53728 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1649977179
transform 1 0 30360 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1649977179
transform 1 0 45172 0 1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1649977179
transform 1 0 42596 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input64
timestamp 1649977179
transform 1 0 3956 0 1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1649977179
transform 1 0 12328 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input66
timestamp 1649977179
transform 1 0 38732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input67
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input68
timestamp 1649977179
transform 1 0 1380 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input69
timestamp 1649977179
transform -1 0 53728 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform -1 0 14628 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform -1 0 37628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform -1 0 13340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform 1 0 53360 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform 1 0 53360 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform 1 0 53360 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform 1 0 40664 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform -1 0 17204 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform 1 0 53360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform 1 0 53360 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform 1 0 51612 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform 1 0 29716 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform -1 0 1748 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform 1 0 53360 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform -1 0 1748 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform -1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform 1 0 36156 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform -1 0 1748 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform 1 0 43240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform 1 0 47564 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform -1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform -1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform -1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform 1 0 51612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform 1 0 53360 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform 1 0 53360 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform -1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform -1 0 1748 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform 1 0 53360 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform -1 0 6716 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform 1 0 53360 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform 1 0 53360 0 1 36992
box -38 -48 406 592
<< labels >>
flabel metal3 s 54697 9528 55497 9648 0 FreeSans 480 0 0 0 alu_branch
port 0 nsew signal input
flabel metal3 s 54697 48288 55497 48408 0 FreeSans 480 0 0 0 branch
port 1 nsew signal input
flabel metal2 s 31574 56841 31630 57641 0 FreeSans 224 90 0 0 clk
port 2 nsew signal input
flabel metal3 s 54697 55088 55497 55208 0 FreeSans 480 0 0 0 immediate[0]
port 3 nsew signal input
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 immediate[10]
port 4 nsew signal input
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 immediate[11]
port 5 nsew signal input
flabel metal3 s 0 52368 800 52488 0 FreeSans 480 0 0 0 immediate[12]
port 6 nsew signal input
flabel metal2 s 53470 56841 53526 57641 0 FreeSans 224 90 0 0 immediate[13]
port 7 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 immediate[14]
port 8 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 immediate[15]
port 9 nsew signal input
flabel metal3 s 0 43528 800 43648 0 FreeSans 480 0 0 0 immediate[16]
port 10 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 immediate[17]
port 11 nsew signal input
flabel metal3 s 0 54408 800 54528 0 FreeSans 480 0 0 0 immediate[18]
port 12 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 immediate[19]
port 13 nsew signal input
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 immediate[1]
port 14 nsew signal input
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 immediate[20]
port 15 nsew signal input
flabel metal3 s 54697 41488 55497 41608 0 FreeSans 480 0 0 0 immediate[21]
port 16 nsew signal input
flabel metal2 s 25134 56841 25190 57641 0 FreeSans 224 90 0 0 immediate[22]
port 17 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 immediate[23]
port 18 nsew signal input
flabel metal3 s 0 36048 800 36168 0 FreeSans 480 0 0 0 immediate[24]
port 19 nsew signal input
flabel metal3 s 0 45568 800 45688 0 FreeSans 480 0 0 0 immediate[25]
port 20 nsew signal input
flabel metal3 s 0 38768 800 38888 0 FreeSans 480 0 0 0 immediate[26]
port 21 nsew signal input
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 immediate[27]
port 22 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 immediate[28]
port 23 nsew signal input
flabel metal3 s 54697 8 55497 128 0 FreeSans 480 0 0 0 immediate[29]
port 24 nsew signal input
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 immediate[2]
port 25 nsew signal input
flabel metal3 s 54697 29928 55497 30048 0 FreeSans 480 0 0 0 immediate[30]
port 26 nsew signal input
flabel metal2 s 34150 56841 34206 57641 0 FreeSans 224 90 0 0 immediate[31]
port 27 nsew signal input
flabel metal2 s 18694 56841 18750 57641 0 FreeSans 224 90 0 0 immediate[3]
port 28 nsew signal input
flabel metal3 s 54697 53048 55497 53168 0 FreeSans 480 0 0 0 immediate[4]
port 29 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 immediate[5]
port 30 nsew signal input
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 immediate[6]
port 31 nsew signal input
flabel metal3 s 54697 50328 55497 50448 0 FreeSans 480 0 0 0 immediate[7]
port 32 nsew signal input
flabel metal2 s 21270 56841 21326 57641 0 FreeSans 224 90 0 0 immediate[8]
port 33 nsew signal input
flabel metal3 s 54697 13608 55497 13728 0 FreeSans 480 0 0 0 immediate[9]
port 34 nsew signal input
flabel metal3 s 54697 18368 55497 18488 0 FreeSans 480 0 0 0 jump_jal
port 35 nsew signal input
flabel metal2 s 23202 56841 23258 57641 0 FreeSans 224 90 0 0 jump_jalr
port 36 nsew signal input
flabel metal2 s 14186 56841 14242 57641 0 FreeSans 224 90 0 0 pc_out[0]
port 37 nsew signal tristate
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 pc_out[10]
port 38 nsew signal tristate
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 pc_out[11]
port 39 nsew signal tristate
flabel metal3 s 54697 43528 55497 43648 0 FreeSans 480 0 0 0 pc_out[12]
port 40 nsew signal tristate
flabel metal2 s 54114 0 54170 800 0 FreeSans 224 90 0 0 pc_out[13]
port 41 nsew signal tristate
flabel metal3 s 54697 23128 55497 23248 0 FreeSans 480 0 0 0 pc_out[14]
port 42 nsew signal tristate
flabel metal2 s 40590 56841 40646 57641 0 FreeSans 224 90 0 0 pc_out[15]
port 43 nsew signal tristate
flabel metal2 s 16762 56841 16818 57641 0 FreeSans 224 90 0 0 pc_out[16]
port 44 nsew signal tristate
flabel metal3 s 54697 2728 55497 2848 0 FreeSans 480 0 0 0 pc_out[17]
port 45 nsew signal tristate
flabel metal3 s 54697 46248 55497 46368 0 FreeSans 480 0 0 0 pc_out[18]
port 46 nsew signal tristate
flabel metal2 s 51538 56841 51594 57641 0 FreeSans 224 90 0 0 pc_out[19]
port 47 nsew signal tristate
flabel metal2 s 29642 56841 29698 57641 0 FreeSans 224 90 0 0 pc_out[1]
port 48 nsew signal tristate
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 pc_out[20]
port 49 nsew signal tristate
flabel metal3 s 54697 11568 55497 11688 0 FreeSans 480 0 0 0 pc_out[21]
port 50 nsew signal tristate
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 pc_out[22]
port 51 nsew signal tristate
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 pc_out[23]
port 52 nsew signal tristate
flabel metal2 s 36082 56841 36138 57641 0 FreeSans 224 90 0 0 pc_out[24]
port 53 nsew signal tristate
flabel metal3 s 0 40808 800 40928 0 FreeSans 480 0 0 0 pc_out[25]
port 54 nsew signal tristate
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 pc_out[26]
port 55 nsew signal tristate
flabel metal2 s 47030 56841 47086 57641 0 FreeSans 224 90 0 0 pc_out[27]
port 56 nsew signal tristate
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 pc_out[28]
port 57 nsew signal tristate
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 pc_out[29]
port 58 nsew signal tristate
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 pc_out[2]
port 59 nsew signal tristate
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 pc_out[30]
port 60 nsew signal tristate
flabel metal3 s 54697 25168 55497 25288 0 FreeSans 480 0 0 0 pc_out[31]
port 61 nsew signal tristate
flabel metal3 s 54697 16328 55497 16448 0 FreeSans 480 0 0 0 pc_out[3]
port 62 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 pc_out[4]
port 63 nsew signal tristate
flabel metal3 s 0 47608 800 47728 0 FreeSans 480 0 0 0 pc_out[5]
port 64 nsew signal tristate
flabel metal3 s 54697 4768 55497 4888 0 FreeSans 480 0 0 0 pc_out[6]
port 65 nsew signal tristate
flabel metal2 s 5814 56841 5870 57641 0 FreeSans 224 90 0 0 pc_out[7]
port 66 nsew signal tristate
flabel metal3 s 54697 21088 55497 21208 0 FreeSans 480 0 0 0 pc_out[8]
port 67 nsew signal tristate
flabel metal3 s 54697 36728 55497 36848 0 FreeSans 480 0 0 0 pc_out[9]
port 68 nsew signal tristate
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 rs1_data[0]
port 69 nsew signal input
flabel metal3 s 54697 39448 55497 39568 0 FreeSans 480 0 0 0 rs1_data[10]
port 70 nsew signal input
flabel metal2 s 7746 56841 7802 57641 0 FreeSans 224 90 0 0 rs1_data[11]
port 71 nsew signal input
flabel metal3 s 0 34008 800 34128 0 FreeSans 480 0 0 0 rs1_data[12]
port 72 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 rs1_data[13]
port 73 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 rs1_data[14]
port 74 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 rs1_data[15]
port 75 nsew signal input
flabel metal2 s 10322 56841 10378 57641 0 FreeSans 224 90 0 0 rs1_data[16]
port 76 nsew signal input
flabel metal2 s 27710 56841 27766 57641 0 FreeSans 224 90 0 0 rs1_data[17]
port 77 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 rs1_data[18]
port 78 nsew signal input
flabel metal3 s 0 57128 800 57248 0 FreeSans 480 0 0 0 rs1_data[19]
port 79 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 rs1_data[1]
port 80 nsew signal input
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 rs1_data[20]
port 81 nsew signal input
flabel metal2 s 48962 56841 49018 57641 0 FreeSans 224 90 0 0 rs1_data[21]
port 82 nsew signal input
flabel metal2 s 38658 56841 38714 57641 0 FreeSans 224 90 0 0 rs1_data[22]
port 83 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 rs1_data[23]
port 84 nsew signal input
flabel metal2 s 55402 56841 55458 57641 0 FreeSans 224 90 0 0 rs1_data[24]
port 85 nsew signal input
flabel metal3 s 54697 6808 55497 6928 0 FreeSans 480 0 0 0 rs1_data[25]
port 86 nsew signal input
flabel metal2 s 1306 56841 1362 57641 0 FreeSans 224 90 0 0 rs1_data[26]
port 87 nsew signal input
flabel metal3 s 54697 31968 55497 32088 0 FreeSans 480 0 0 0 rs1_data[27]
port 88 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 rs1_data[28]
port 89 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 rs1_data[29]
port 90 nsew signal input
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 rs1_data[2]
port 91 nsew signal input
flabel metal3 s 54697 34688 55497 34808 0 FreeSans 480 0 0 0 rs1_data[30]
port 92 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 rs1_data[31]
port 93 nsew signal input
flabel metal2 s 45098 56841 45154 57641 0 FreeSans 224 90 0 0 rs1_data[3]
port 94 nsew signal input
flabel metal2 s 42522 56841 42578 57641 0 FreeSans 224 90 0 0 rs1_data[4]
port 95 nsew signal input
flabel metal2 s 3882 56841 3938 57641 0 FreeSans 224 90 0 0 rs1_data[5]
port 96 nsew signal input
flabel metal2 s 12254 56841 12310 57641 0 FreeSans 224 90 0 0 rs1_data[6]
port 97 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 rs1_data[7]
port 98 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 rs1_data[8]
port 99 nsew signal input
flabel metal3 s 0 50328 800 50448 0 FreeSans 480 0 0 0 rs1_data[9]
port 100 nsew signal input
flabel metal3 s 54697 27888 55497 28008 0 FreeSans 480 0 0 0 rst_n
port 101 nsew signal input
flabel metal4 s 4208 2128 4528 54992 0 FreeSans 1920 90 0 0 vccd1
port 102 nsew power bidirectional
flabel metal4 s 34928 2128 35248 54992 0 FreeSans 1920 90 0 0 vccd1
port 102 nsew power bidirectional
flabel metal4 s 19568 2128 19888 54992 0 FreeSans 1920 90 0 0 vssd1
port 103 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 54992 0 FreeSans 1920 90 0 0 vssd1
port 103 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 55497 57641
<< end >>
