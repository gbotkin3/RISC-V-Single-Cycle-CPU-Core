VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RISC_V
  CLASS BLOCK ;
  FOREIGN RISC_V ;
  ORIGIN 0.000 0.000 ;
  SIZE 2820.000 BY 3420.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1329.440 4.000 1330.040 ;
    END
  END clk
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2614.730 3416.000 2615.010 3420.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2266.970 3416.000 2267.250 3420.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1927.840 4.000 1928.440 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1761.240 4.000 1761.840 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 809.240 2820.000 809.840 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2791.440 4.000 2792.040 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 3416.000 1008.230 3420.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 3416.000 821.470 3420.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.030 3416.000 1858.310 3420.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 941.840 2820.000 942.440 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2489.150 3416.000 2489.430 3420.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2060.440 4.000 2061.040 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.650 0.000 1603.930 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1241.040 2820.000 1241.640 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2708.110 3416.000 2708.390 3420.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2556.840 4.000 2557.440 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 3236.840 2820.000 3237.440 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2138.640 2820.000 2139.240 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2737.090 0.000 2737.370 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2141.390 3416.000 2141.670 3420.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1919.210 0.000 1919.490 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3124.640 4.000 3125.240 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 3416.000 947.050 3420.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2937.640 2820.000 2938.240 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1373.640 2820.000 1374.240 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3056.640 4.000 3057.240 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.010 3416.000 2048.290 3420.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2536.440 2820.000 2537.040 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 0.000 692.670 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1907.440 2820.000 1908.040 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 146.240 2820.000 146.840 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.810 0.000 1855.090 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.240 4.000 996.840 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1030.240 4.000 1030.840 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 975.840 2820.000 976.440 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 3202.840 2820.000 3203.440 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2675.910 0.000 2676.190 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2373.240 2820.000 2373.840 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 3403.440 2820.000 3404.040 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1980.390 0.000 1980.670 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 3416.000 538.110 3420.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 3416.000 473.710 3420.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.510 3416.000 1323.790 3420.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2390.240 4.000 2390.840 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2771.040 2820.000 2771.640 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1774.840 2820.000 1775.440 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3321.840 4.000 3322.440 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 10.240 2820.000 10.840 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 642.640 2820.000 643.240 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2206.640 2820.000 2207.240 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 3369.440 2820.000 3370.040 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1638.840 2820.000 1639.440 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 3070.240 2820.000 3070.840 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2325.640 4.000 2326.240 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.450 3416.000 1732.730 3420.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2492.240 4.000 2492.840 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 0.000 721.650 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2611.510 0.000 2611.790 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.330 3416.000 1262.610 3420.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2138.170 0.000 2138.450 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2205.790 3416.000 2206.070 3420.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 112.240 2820.000 112.840 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.030 0.000 1697.310 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.690 3416.000 1545.970 3420.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.470 0.000 1542.750 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2805.040 2820.000 2805.640 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 3416.000 1072.630 3420.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1873.440 2820.000 1874.040 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2360.350 0.000 2360.630 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2638.440 2820.000 2639.040 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2604.440 2820.000 2605.040 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.290 0.000 1320.570 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2091.040 4.000 2091.640 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 843.240 2820.000 843.840 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 3416.000 380.330 3420.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2421.530 0.000 2421.810 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 278.840 2820.000 279.440 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3257.240 4.000 3257.840 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1193.440 4.000 1194.040 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 3270.840 2820.000 3271.440 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.310 0.000 1130.590 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.670 0.000 1413.950 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 3416.000 283.730 3420.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 3002.240 2820.000 3002.840 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 3416.000 567.090 3420.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3389.840 4.000 3390.440 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2424.240 4.000 2424.840 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 3416.000 222.550 3420.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1009.840 2820.000 1010.440 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 0.000 911.630 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.730 3416.000 1166.010 3420.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 3416.000 1291.590 3420.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 544.040 2820.000 544.640 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 0.000 786.050 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.670 3416.000 1574.950 3420.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2403.840 2820.000 2404.440 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 442.040 2820.000 442.640 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2804.710 3416.000 2804.990 3420.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1825.840 4.000 1826.440 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1606.870 3416.000 1607.150 3420.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2424.750 3416.000 2425.030 3420.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2869.640 2820.000 2870.240 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2835.640 2820.000 2836.240 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1394.040 4.000 1394.640 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 0.000 596.070 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 3416.000 96.970 3420.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2227.040 4.000 2227.640 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1259.110 0.000 1259.390 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.730 0.000 1005.010 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2643.710 0.000 2643.990 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 0.000 847.230 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3189.240 4.000 3189.840 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2257.640 4.000 2258.240 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 3416.000 695.890 3420.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 962.240 4.000 962.840 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 3416.000 1198.210 3420.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1441.640 2820.000 1442.240 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.910 0.000 1227.190 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 741.240 2820.000 741.840 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3223.240 4.000 3223.840 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 608.640 2820.000 609.240 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.240 4.000 928.840 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2769.290 0.000 2769.570 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 0.000 976.030 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2331.370 3416.000 2331.650 3420.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1958.440 4.000 1959.040 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 3416.000 32.570 3420.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1384.690 0.000 1384.970 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3022.640 4.000 3023.240 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.290 3416.000 1481.570 3420.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.070 3416.000 1639.350 3420.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 907.840 2820.000 908.440 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 3104.240 2820.000 3104.840 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.930 0.000 2486.210 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1339.640 2820.000 1340.240 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1407.640 2820.000 1408.240 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1951.410 0.000 1951.690 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.930 0.000 1037.210 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1074.440 2820.000 1075.040 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2737.040 2820.000 2737.640 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2291.640 4.000 2292.240 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2305.240 2820.000 2305.840 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1992.440 4.000 1993.040 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1275.040 2820.000 1275.640 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3355.840 4.000 3356.440 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1972.040 2820.000 1972.640 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.270 3416.000 1671.550 3420.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 775.240 2820.000 775.840 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.890 3416.000 1417.170 3420.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 3416.000 441.510 3420.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2271.240 2820.000 2271.840 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.710 0.000 1194.990 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.130 0.000 1069.410 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1309.040 2820.000 1309.640 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 3416.000 757.070 3420.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 3416.000 254.750 3420.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 510.040 2820.000 510.640 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.490 0.000 1352.770 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2456.950 3416.000 2457.230 3420.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2339.240 2820.000 2339.840 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3090.640 4.000 3091.240 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1295.440 4.000 1296.040 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1761.430 0.000 1761.710 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 3416.000 505.910 3420.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2363.570 3416.000 2363.850 3420.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2471.840 2820.000 2472.440 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2689.440 4.000 2690.040 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 3416.000 0.370 3420.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.250 3416.000 1700.530 3420.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2458.240 4.000 2458.840 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2547.110 0.000 2547.390 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1540.240 2820.000 1540.840 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 343.440 2820.000 344.040 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.530 3416.000 1133.810 3420.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.450 0.000 1571.730 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3155.240 4.000 3155.840 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.870 0.000 1446.150 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 710.640 2820.000 711.240 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2521.350 3416.000 2521.630 3420.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.040 4.000 629.640 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.490 3416.000 1513.770 3420.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1128.840 4.000 1129.440 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2646.930 3416.000 2647.210 3420.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 3416.000 315.930 3420.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 863.640 4.000 864.240 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 244.840 2820.000 245.440 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2924.040 4.000 2924.640 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2723.440 4.000 2724.040 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.630 0.000 1793.910 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1475.640 2820.000 1476.240 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1176.440 2820.000 1177.040 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 3416.000 850.450 3420.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1740.840 2820.000 1741.440 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2170.370 0.000 2170.650 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2109.190 0.000 2109.470 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2518.130 0.000 2518.410 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2159.040 4.000 2159.640 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.950 0.000 2296.230 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1492.640 4.000 1493.240 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2359.640 4.000 2360.240 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 3335.440 2820.000 3336.040 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1727.240 4.000 1727.840 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 0.000 818.250 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1938.040 2820.000 1938.640 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.310 0.000 2579.590 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2173.590 3416.000 2173.870 3420.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 3416.000 412.530 3420.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2971.640 2820.000 2972.240 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.840 4.000 1163.440 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2703.040 2820.000 2703.640 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.090 3416.000 1449.370 3420.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1428.040 4.000 1428.640 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1893.840 4.000 1894.440 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.550 3416.000 1104.830 3420.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 3416.000 631.490 3420.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1510.270 0.000 1510.550 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 210.840 2820.000 211.440 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 3301.440 2820.000 3302.040 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 476.040 2820.000 476.640 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.130 3416.000 1230.410 3420.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1288.090 0.000 1288.370 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2550.330 3416.000 2550.610 3420.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2590.840 4.000 2591.440 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.330 0.000 1101.610 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1608.240 2820.000 1608.840 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2890.040 4.000 2890.640 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2263.750 0.000 2264.030 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 78.240 2820.000 78.840 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2074.040 2820.000 2074.640 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2080.210 3416.000 2080.490 3420.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1706.840 2820.000 1707.440 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2526.240 4.000 2526.840 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1859.840 4.000 1860.440 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 411.440 2820.000 412.040 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1829.050 3416.000 1829.330 3420.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2704.890 0.000 2705.170 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 3416.000 158.150 3420.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1672.840 2820.000 1673.440 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3287.840 4.000 3288.440 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2172.640 2820.000 2173.240 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2801.490 0.000 2801.770 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 3416.000 914.850 3420.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2582.530 3416.000 2582.810 3420.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2505.840 2820.000 2506.440 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 3416.000 789.270 3420.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 3416.000 1040.430 3420.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 676.640 2820.000 677.240 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1693.240 4.000 1693.840 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1526.640 4.000 1527.240 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1983.610 3416.000 1983.890 3420.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.710 3416.000 1355.990 3420.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 3416.000 190.350 3420.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1261.440 4.000 1262.040 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2988.640 4.000 2989.240 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2437.840 2820.000 2438.440 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2237.240 2820.000 2237.840 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.010 0.000 1887.290 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2040.040 2820.000 2040.640 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1560.640 4.000 1561.240 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 44.240 2820.000 44.840 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1890.230 3416.000 1890.510 3420.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2740.310 3416.000 2740.590 3420.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.050 0.000 1668.330 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.240 4.000 894.840 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 877.240 2820.000 877.840 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 3416.000 348.130 3420.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 3416.000 979.250 3420.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1227.440 4.000 1228.040 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 3168.840 2820.000 3169.440 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2299.170 3416.000 2299.450 3420.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1506.240 2820.000 1506.840 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2328.150 0.000 2328.430 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1360.040 4.000 1360.640 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2234.770 0.000 2235.050 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1659.240 4.000 1659.840 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2193.040 4.000 2193.640 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 176.840 2820.000 177.440 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1040.440 2820.000 1041.040 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 3416.000 882.650 3420.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2903.640 2820.000 2904.240 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2624.840 4.000 2625.440 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2856.040 4.000 2856.640 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2757.440 4.000 2758.040 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1839.440 2820.000 1840.040 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.230 0.000 1729.510 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1954.630 3416.000 1954.910 3420.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2679.130 3416.000 2679.410 3420.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 3416.000 64.770 3420.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1462.040 4.000 1462.640 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1628.640 4.000 1629.240 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2772.510 3416.000 2772.790 3420.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2026.440 4.000 2027.040 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1207.040 2820.000 1207.640 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2076.990 0.000 2077.270 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2395.770 3416.000 2396.050 3420.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 3416.000 599.290 3420.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 0.000 943.830 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2104.640 2820.000 2105.240 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2453.730 0.000 2454.010 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1142.440 2820.000 1143.040 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1791.840 4.000 1792.440 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 309.440 2820.000 310.040 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.070 0.000 1478.350 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1574.240 2820.000 1574.840 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2237.990 3416.000 2238.270 3420.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 3036.240 2820.000 3036.840 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 377.440 2820.000 378.040 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2006.040 2820.000 2006.640 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 3134.840 2820.000 3135.440 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.410 3416.000 2112.690 3420.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 578.040 2820.000 578.640 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2015.810 3416.000 2016.090 3420.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2044.790 0.000 2045.070 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1060.840 4.000 1061.440 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.590 0.000 2012.870 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.550 0.000 2392.830 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1594.640 4.000 1595.240 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2825.440 4.000 2826.040 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 3416.000 663.690 3420.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1094.840 4.000 1095.440 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 0.000 628.270 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.910 3416.000 1388.190 3420.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 3416.000 724.870 3420.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1635.850 0.000 1636.130 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.430 3416.000 1922.710 3420.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1108.440 2820.000 1109.040 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2125.040 4.000 2125.640 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2672.440 2820.000 2673.040 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 0.000 1162.790 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 2570.440 2820.000 2571.040 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1825.830 0.000 1826.110 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1796.850 3416.000 1797.130 3420.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.650 3416.000 1764.930 3420.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2958.040 4.000 2958.640 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 3416.000 129.170 3420.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2202.570 0.000 2202.850 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2658.840 4.000 2659.440 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2816.000 1805.440 2820.000 1806.040 ;
    END
  END la_oenb[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2632.240 10.640 2633.840 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2785.840 10.640 2787.440 3408.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 3408.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2709.040 10.640 2710.640 3408.400 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2814.280 3408.245 ;
      LAYER met1 ;
        RECT 0.070 10.640 2814.280 3408.400 ;
      LAYER met2 ;
        RECT 0.650 3415.720 32.010 3416.730 ;
        RECT 32.850 3415.720 64.210 3416.730 ;
        RECT 65.050 3415.720 96.410 3416.730 ;
        RECT 97.250 3415.720 128.610 3416.730 ;
        RECT 129.450 3415.720 157.590 3416.730 ;
        RECT 158.430 3415.720 189.790 3416.730 ;
        RECT 190.630 3415.720 221.990 3416.730 ;
        RECT 222.830 3415.720 254.190 3416.730 ;
        RECT 255.030 3415.720 283.170 3416.730 ;
        RECT 284.010 3415.720 315.370 3416.730 ;
        RECT 316.210 3415.720 347.570 3416.730 ;
        RECT 348.410 3415.720 379.770 3416.730 ;
        RECT 380.610 3415.720 411.970 3416.730 ;
        RECT 412.810 3415.720 440.950 3416.730 ;
        RECT 441.790 3415.720 473.150 3416.730 ;
        RECT 473.990 3415.720 505.350 3416.730 ;
        RECT 506.190 3415.720 537.550 3416.730 ;
        RECT 538.390 3415.720 566.530 3416.730 ;
        RECT 567.370 3415.720 598.730 3416.730 ;
        RECT 599.570 3415.720 630.930 3416.730 ;
        RECT 631.770 3415.720 663.130 3416.730 ;
        RECT 663.970 3415.720 695.330 3416.730 ;
        RECT 696.170 3415.720 724.310 3416.730 ;
        RECT 725.150 3415.720 756.510 3416.730 ;
        RECT 757.350 3415.720 788.710 3416.730 ;
        RECT 789.550 3415.720 820.910 3416.730 ;
        RECT 821.750 3415.720 849.890 3416.730 ;
        RECT 850.730 3415.720 882.090 3416.730 ;
        RECT 882.930 3415.720 914.290 3416.730 ;
        RECT 915.130 3415.720 946.490 3416.730 ;
        RECT 947.330 3415.720 978.690 3416.730 ;
        RECT 979.530 3415.720 1007.670 3416.730 ;
        RECT 1008.510 3415.720 1039.870 3416.730 ;
        RECT 1040.710 3415.720 1072.070 3416.730 ;
        RECT 1072.910 3415.720 1104.270 3416.730 ;
        RECT 1105.110 3415.720 1133.250 3416.730 ;
        RECT 1134.090 3415.720 1165.450 3416.730 ;
        RECT 1166.290 3415.720 1197.650 3416.730 ;
        RECT 1198.490 3415.720 1229.850 3416.730 ;
        RECT 1230.690 3415.720 1262.050 3416.730 ;
        RECT 1262.890 3415.720 1291.030 3416.730 ;
        RECT 1291.870 3415.720 1323.230 3416.730 ;
        RECT 1324.070 3415.720 1355.430 3416.730 ;
        RECT 1356.270 3415.720 1387.630 3416.730 ;
        RECT 1388.470 3415.720 1416.610 3416.730 ;
        RECT 1417.450 3415.720 1448.810 3416.730 ;
        RECT 1449.650 3415.720 1481.010 3416.730 ;
        RECT 1481.850 3415.720 1513.210 3416.730 ;
        RECT 1514.050 3415.720 1545.410 3416.730 ;
        RECT 1546.250 3415.720 1574.390 3416.730 ;
        RECT 1575.230 3415.720 1606.590 3416.730 ;
        RECT 1607.430 3415.720 1638.790 3416.730 ;
        RECT 1639.630 3415.720 1670.990 3416.730 ;
        RECT 1671.830 3415.720 1699.970 3416.730 ;
        RECT 1700.810 3415.720 1732.170 3416.730 ;
        RECT 1733.010 3415.720 1764.370 3416.730 ;
        RECT 1765.210 3415.720 1796.570 3416.730 ;
        RECT 1797.410 3415.720 1828.770 3416.730 ;
        RECT 1829.610 3415.720 1857.750 3416.730 ;
        RECT 1858.590 3415.720 1889.950 3416.730 ;
        RECT 1890.790 3415.720 1922.150 3416.730 ;
        RECT 1922.990 3415.720 1954.350 3416.730 ;
        RECT 1955.190 3415.720 1983.330 3416.730 ;
        RECT 1984.170 3415.720 2015.530 3416.730 ;
        RECT 2016.370 3415.720 2047.730 3416.730 ;
        RECT 2048.570 3415.720 2079.930 3416.730 ;
        RECT 2080.770 3415.720 2112.130 3416.730 ;
        RECT 2112.970 3415.720 2141.110 3416.730 ;
        RECT 2141.950 3415.720 2173.310 3416.730 ;
        RECT 2174.150 3415.720 2205.510 3416.730 ;
        RECT 2206.350 3415.720 2237.710 3416.730 ;
        RECT 2238.550 3415.720 2266.690 3416.730 ;
        RECT 2267.530 3415.720 2298.890 3416.730 ;
        RECT 2299.730 3415.720 2331.090 3416.730 ;
        RECT 2331.930 3415.720 2363.290 3416.730 ;
        RECT 2364.130 3415.720 2395.490 3416.730 ;
        RECT 2396.330 3415.720 2424.470 3416.730 ;
        RECT 2425.310 3415.720 2456.670 3416.730 ;
        RECT 2457.510 3415.720 2488.870 3416.730 ;
        RECT 2489.710 3415.720 2521.070 3416.730 ;
        RECT 2521.910 3415.720 2550.050 3416.730 ;
        RECT 2550.890 3415.720 2582.250 3416.730 ;
        RECT 2583.090 3415.720 2614.450 3416.730 ;
        RECT 2615.290 3415.720 2646.650 3416.730 ;
        RECT 2647.490 3415.720 2678.850 3416.730 ;
        RECT 2679.690 3415.720 2707.830 3416.730 ;
        RECT 2708.670 3415.720 2740.030 3416.730 ;
        RECT 2740.870 3415.720 2772.230 3416.730 ;
        RECT 2773.070 3415.720 2804.430 3416.730 ;
        RECT 2805.270 3415.720 2810.970 3416.730 ;
        RECT 0.100 4.280 2810.970 3415.720 ;
        RECT 0.650 4.000 28.790 4.280 ;
        RECT 29.630 4.000 60.990 4.280 ;
        RECT 61.830 4.000 93.190 4.280 ;
        RECT 94.030 4.000 125.390 4.280 ;
        RECT 126.230 4.000 154.370 4.280 ;
        RECT 155.210 4.000 186.570 4.280 ;
        RECT 187.410 4.000 218.770 4.280 ;
        RECT 219.610 4.000 250.970 4.280 ;
        RECT 251.810 4.000 279.950 4.280 ;
        RECT 280.790 4.000 312.150 4.280 ;
        RECT 312.990 4.000 344.350 4.280 ;
        RECT 345.190 4.000 376.550 4.280 ;
        RECT 377.390 4.000 408.750 4.280 ;
        RECT 409.590 4.000 437.730 4.280 ;
        RECT 438.570 4.000 469.930 4.280 ;
        RECT 470.770 4.000 502.130 4.280 ;
        RECT 502.970 4.000 534.330 4.280 ;
        RECT 535.170 4.000 563.310 4.280 ;
        RECT 564.150 4.000 595.510 4.280 ;
        RECT 596.350 4.000 627.710 4.280 ;
        RECT 628.550 4.000 659.910 4.280 ;
        RECT 660.750 4.000 692.110 4.280 ;
        RECT 692.950 4.000 721.090 4.280 ;
        RECT 721.930 4.000 753.290 4.280 ;
        RECT 754.130 4.000 785.490 4.280 ;
        RECT 786.330 4.000 817.690 4.280 ;
        RECT 818.530 4.000 846.670 4.280 ;
        RECT 847.510 4.000 878.870 4.280 ;
        RECT 879.710 4.000 911.070 4.280 ;
        RECT 911.910 4.000 943.270 4.280 ;
        RECT 944.110 4.000 975.470 4.280 ;
        RECT 976.310 4.000 1004.450 4.280 ;
        RECT 1005.290 4.000 1036.650 4.280 ;
        RECT 1037.490 4.000 1068.850 4.280 ;
        RECT 1069.690 4.000 1101.050 4.280 ;
        RECT 1101.890 4.000 1130.030 4.280 ;
        RECT 1130.870 4.000 1162.230 4.280 ;
        RECT 1163.070 4.000 1194.430 4.280 ;
        RECT 1195.270 4.000 1226.630 4.280 ;
        RECT 1227.470 4.000 1258.830 4.280 ;
        RECT 1259.670 4.000 1287.810 4.280 ;
        RECT 1288.650 4.000 1320.010 4.280 ;
        RECT 1320.850 4.000 1352.210 4.280 ;
        RECT 1353.050 4.000 1384.410 4.280 ;
        RECT 1385.250 4.000 1413.390 4.280 ;
        RECT 1414.230 4.000 1445.590 4.280 ;
        RECT 1446.430 4.000 1477.790 4.280 ;
        RECT 1478.630 4.000 1509.990 4.280 ;
        RECT 1510.830 4.000 1542.190 4.280 ;
        RECT 1543.030 4.000 1571.170 4.280 ;
        RECT 1572.010 4.000 1603.370 4.280 ;
        RECT 1604.210 4.000 1635.570 4.280 ;
        RECT 1636.410 4.000 1667.770 4.280 ;
        RECT 1668.610 4.000 1696.750 4.280 ;
        RECT 1697.590 4.000 1728.950 4.280 ;
        RECT 1729.790 4.000 1761.150 4.280 ;
        RECT 1761.990 4.000 1793.350 4.280 ;
        RECT 1794.190 4.000 1825.550 4.280 ;
        RECT 1826.390 4.000 1854.530 4.280 ;
        RECT 1855.370 4.000 1886.730 4.280 ;
        RECT 1887.570 4.000 1918.930 4.280 ;
        RECT 1919.770 4.000 1951.130 4.280 ;
        RECT 1951.970 4.000 1980.110 4.280 ;
        RECT 1980.950 4.000 2012.310 4.280 ;
        RECT 2013.150 4.000 2044.510 4.280 ;
        RECT 2045.350 4.000 2076.710 4.280 ;
        RECT 2077.550 4.000 2108.910 4.280 ;
        RECT 2109.750 4.000 2137.890 4.280 ;
        RECT 2138.730 4.000 2170.090 4.280 ;
        RECT 2170.930 4.000 2202.290 4.280 ;
        RECT 2203.130 4.000 2234.490 4.280 ;
        RECT 2235.330 4.000 2263.470 4.280 ;
        RECT 2264.310 4.000 2295.670 4.280 ;
        RECT 2296.510 4.000 2327.870 4.280 ;
        RECT 2328.710 4.000 2360.070 4.280 ;
        RECT 2360.910 4.000 2392.270 4.280 ;
        RECT 2393.110 4.000 2421.250 4.280 ;
        RECT 2422.090 4.000 2453.450 4.280 ;
        RECT 2454.290 4.000 2485.650 4.280 ;
        RECT 2486.490 4.000 2517.850 4.280 ;
        RECT 2518.690 4.000 2546.830 4.280 ;
        RECT 2547.670 4.000 2579.030 4.280 ;
        RECT 2579.870 4.000 2611.230 4.280 ;
        RECT 2612.070 4.000 2643.430 4.280 ;
        RECT 2644.270 4.000 2675.630 4.280 ;
        RECT 2676.470 4.000 2704.610 4.280 ;
        RECT 2705.450 4.000 2736.810 4.280 ;
        RECT 2737.650 4.000 2769.010 4.280 ;
        RECT 2769.850 4.000 2801.210 4.280 ;
        RECT 2802.050 4.000 2810.970 4.280 ;
      LAYER met3 ;
        RECT 4.000 3404.440 2816.000 3408.325 ;
        RECT 4.000 3403.040 2815.600 3404.440 ;
        RECT 4.000 3390.840 2816.000 3403.040 ;
        RECT 4.400 3389.440 2816.000 3390.840 ;
        RECT 4.000 3370.440 2816.000 3389.440 ;
        RECT 4.000 3369.040 2815.600 3370.440 ;
        RECT 4.000 3356.840 2816.000 3369.040 ;
        RECT 4.400 3355.440 2816.000 3356.840 ;
        RECT 4.000 3336.440 2816.000 3355.440 ;
        RECT 4.000 3335.040 2815.600 3336.440 ;
        RECT 4.000 3322.840 2816.000 3335.040 ;
        RECT 4.400 3321.440 2816.000 3322.840 ;
        RECT 4.000 3302.440 2816.000 3321.440 ;
        RECT 4.000 3301.040 2815.600 3302.440 ;
        RECT 4.000 3288.840 2816.000 3301.040 ;
        RECT 4.400 3287.440 2816.000 3288.840 ;
        RECT 4.000 3271.840 2816.000 3287.440 ;
        RECT 4.000 3270.440 2815.600 3271.840 ;
        RECT 4.000 3258.240 2816.000 3270.440 ;
        RECT 4.400 3256.840 2816.000 3258.240 ;
        RECT 4.000 3237.840 2816.000 3256.840 ;
        RECT 4.000 3236.440 2815.600 3237.840 ;
        RECT 4.000 3224.240 2816.000 3236.440 ;
        RECT 4.400 3222.840 2816.000 3224.240 ;
        RECT 4.000 3203.840 2816.000 3222.840 ;
        RECT 4.000 3202.440 2815.600 3203.840 ;
        RECT 4.000 3190.240 2816.000 3202.440 ;
        RECT 4.400 3188.840 2816.000 3190.240 ;
        RECT 4.000 3169.840 2816.000 3188.840 ;
        RECT 4.000 3168.440 2815.600 3169.840 ;
        RECT 4.000 3156.240 2816.000 3168.440 ;
        RECT 4.400 3154.840 2816.000 3156.240 ;
        RECT 4.000 3135.840 2816.000 3154.840 ;
        RECT 4.000 3134.440 2815.600 3135.840 ;
        RECT 4.000 3125.640 2816.000 3134.440 ;
        RECT 4.400 3124.240 2816.000 3125.640 ;
        RECT 4.000 3105.240 2816.000 3124.240 ;
        RECT 4.000 3103.840 2815.600 3105.240 ;
        RECT 4.000 3091.640 2816.000 3103.840 ;
        RECT 4.400 3090.240 2816.000 3091.640 ;
        RECT 4.000 3071.240 2816.000 3090.240 ;
        RECT 4.000 3069.840 2815.600 3071.240 ;
        RECT 4.000 3057.640 2816.000 3069.840 ;
        RECT 4.400 3056.240 2816.000 3057.640 ;
        RECT 4.000 3037.240 2816.000 3056.240 ;
        RECT 4.000 3035.840 2815.600 3037.240 ;
        RECT 4.000 3023.640 2816.000 3035.840 ;
        RECT 4.400 3022.240 2816.000 3023.640 ;
        RECT 4.000 3003.240 2816.000 3022.240 ;
        RECT 4.000 3001.840 2815.600 3003.240 ;
        RECT 4.000 2989.640 2816.000 3001.840 ;
        RECT 4.400 2988.240 2816.000 2989.640 ;
        RECT 4.000 2972.640 2816.000 2988.240 ;
        RECT 4.000 2971.240 2815.600 2972.640 ;
        RECT 4.000 2959.040 2816.000 2971.240 ;
        RECT 4.400 2957.640 2816.000 2959.040 ;
        RECT 4.000 2938.640 2816.000 2957.640 ;
        RECT 4.000 2937.240 2815.600 2938.640 ;
        RECT 4.000 2925.040 2816.000 2937.240 ;
        RECT 4.400 2923.640 2816.000 2925.040 ;
        RECT 4.000 2904.640 2816.000 2923.640 ;
        RECT 4.000 2903.240 2815.600 2904.640 ;
        RECT 4.000 2891.040 2816.000 2903.240 ;
        RECT 4.400 2889.640 2816.000 2891.040 ;
        RECT 4.000 2870.640 2816.000 2889.640 ;
        RECT 4.000 2869.240 2815.600 2870.640 ;
        RECT 4.000 2857.040 2816.000 2869.240 ;
        RECT 4.400 2855.640 2816.000 2857.040 ;
        RECT 4.000 2836.640 2816.000 2855.640 ;
        RECT 4.000 2835.240 2815.600 2836.640 ;
        RECT 4.000 2826.440 2816.000 2835.240 ;
        RECT 4.400 2825.040 2816.000 2826.440 ;
        RECT 4.000 2806.040 2816.000 2825.040 ;
        RECT 4.000 2804.640 2815.600 2806.040 ;
        RECT 4.000 2792.440 2816.000 2804.640 ;
        RECT 4.400 2791.040 2816.000 2792.440 ;
        RECT 4.000 2772.040 2816.000 2791.040 ;
        RECT 4.000 2770.640 2815.600 2772.040 ;
        RECT 4.000 2758.440 2816.000 2770.640 ;
        RECT 4.400 2757.040 2816.000 2758.440 ;
        RECT 4.000 2738.040 2816.000 2757.040 ;
        RECT 4.000 2736.640 2815.600 2738.040 ;
        RECT 4.000 2724.440 2816.000 2736.640 ;
        RECT 4.400 2723.040 2816.000 2724.440 ;
        RECT 4.000 2704.040 2816.000 2723.040 ;
        RECT 4.000 2702.640 2815.600 2704.040 ;
        RECT 4.000 2690.440 2816.000 2702.640 ;
        RECT 4.400 2689.040 2816.000 2690.440 ;
        RECT 4.000 2673.440 2816.000 2689.040 ;
        RECT 4.000 2672.040 2815.600 2673.440 ;
        RECT 4.000 2659.840 2816.000 2672.040 ;
        RECT 4.400 2658.440 2816.000 2659.840 ;
        RECT 4.000 2639.440 2816.000 2658.440 ;
        RECT 4.000 2638.040 2815.600 2639.440 ;
        RECT 4.000 2625.840 2816.000 2638.040 ;
        RECT 4.400 2624.440 2816.000 2625.840 ;
        RECT 4.000 2605.440 2816.000 2624.440 ;
        RECT 4.000 2604.040 2815.600 2605.440 ;
        RECT 4.000 2591.840 2816.000 2604.040 ;
        RECT 4.400 2590.440 2816.000 2591.840 ;
        RECT 4.000 2571.440 2816.000 2590.440 ;
        RECT 4.000 2570.040 2815.600 2571.440 ;
        RECT 4.000 2557.840 2816.000 2570.040 ;
        RECT 4.400 2556.440 2816.000 2557.840 ;
        RECT 4.000 2537.440 2816.000 2556.440 ;
        RECT 4.000 2536.040 2815.600 2537.440 ;
        RECT 4.000 2527.240 2816.000 2536.040 ;
        RECT 4.400 2525.840 2816.000 2527.240 ;
        RECT 4.000 2506.840 2816.000 2525.840 ;
        RECT 4.000 2505.440 2815.600 2506.840 ;
        RECT 4.000 2493.240 2816.000 2505.440 ;
        RECT 4.400 2491.840 2816.000 2493.240 ;
        RECT 4.000 2472.840 2816.000 2491.840 ;
        RECT 4.000 2471.440 2815.600 2472.840 ;
        RECT 4.000 2459.240 2816.000 2471.440 ;
        RECT 4.400 2457.840 2816.000 2459.240 ;
        RECT 4.000 2438.840 2816.000 2457.840 ;
        RECT 4.000 2437.440 2815.600 2438.840 ;
        RECT 4.000 2425.240 2816.000 2437.440 ;
        RECT 4.400 2423.840 2816.000 2425.240 ;
        RECT 4.000 2404.840 2816.000 2423.840 ;
        RECT 4.000 2403.440 2815.600 2404.840 ;
        RECT 4.000 2391.240 2816.000 2403.440 ;
        RECT 4.400 2389.840 2816.000 2391.240 ;
        RECT 4.000 2374.240 2816.000 2389.840 ;
        RECT 4.000 2372.840 2815.600 2374.240 ;
        RECT 4.000 2360.640 2816.000 2372.840 ;
        RECT 4.400 2359.240 2816.000 2360.640 ;
        RECT 4.000 2340.240 2816.000 2359.240 ;
        RECT 4.000 2338.840 2815.600 2340.240 ;
        RECT 4.000 2326.640 2816.000 2338.840 ;
        RECT 4.400 2325.240 2816.000 2326.640 ;
        RECT 4.000 2306.240 2816.000 2325.240 ;
        RECT 4.000 2304.840 2815.600 2306.240 ;
        RECT 4.000 2292.640 2816.000 2304.840 ;
        RECT 4.400 2291.240 2816.000 2292.640 ;
        RECT 4.000 2272.240 2816.000 2291.240 ;
        RECT 4.000 2270.840 2815.600 2272.240 ;
        RECT 4.000 2258.640 2816.000 2270.840 ;
        RECT 4.400 2257.240 2816.000 2258.640 ;
        RECT 4.000 2238.240 2816.000 2257.240 ;
        RECT 4.000 2236.840 2815.600 2238.240 ;
        RECT 4.000 2228.040 2816.000 2236.840 ;
        RECT 4.400 2226.640 2816.000 2228.040 ;
        RECT 4.000 2207.640 2816.000 2226.640 ;
        RECT 4.000 2206.240 2815.600 2207.640 ;
        RECT 4.000 2194.040 2816.000 2206.240 ;
        RECT 4.400 2192.640 2816.000 2194.040 ;
        RECT 4.000 2173.640 2816.000 2192.640 ;
        RECT 4.000 2172.240 2815.600 2173.640 ;
        RECT 4.000 2160.040 2816.000 2172.240 ;
        RECT 4.400 2158.640 2816.000 2160.040 ;
        RECT 4.000 2139.640 2816.000 2158.640 ;
        RECT 4.000 2138.240 2815.600 2139.640 ;
        RECT 4.000 2126.040 2816.000 2138.240 ;
        RECT 4.400 2124.640 2816.000 2126.040 ;
        RECT 4.000 2105.640 2816.000 2124.640 ;
        RECT 4.000 2104.240 2815.600 2105.640 ;
        RECT 4.000 2092.040 2816.000 2104.240 ;
        RECT 4.400 2090.640 2816.000 2092.040 ;
        RECT 4.000 2075.040 2816.000 2090.640 ;
        RECT 4.000 2073.640 2815.600 2075.040 ;
        RECT 4.000 2061.440 2816.000 2073.640 ;
        RECT 4.400 2060.040 2816.000 2061.440 ;
        RECT 4.000 2041.040 2816.000 2060.040 ;
        RECT 4.000 2039.640 2815.600 2041.040 ;
        RECT 4.000 2027.440 2816.000 2039.640 ;
        RECT 4.400 2026.040 2816.000 2027.440 ;
        RECT 4.000 2007.040 2816.000 2026.040 ;
        RECT 4.000 2005.640 2815.600 2007.040 ;
        RECT 4.000 1993.440 2816.000 2005.640 ;
        RECT 4.400 1992.040 2816.000 1993.440 ;
        RECT 4.000 1973.040 2816.000 1992.040 ;
        RECT 4.000 1971.640 2815.600 1973.040 ;
        RECT 4.000 1959.440 2816.000 1971.640 ;
        RECT 4.400 1958.040 2816.000 1959.440 ;
        RECT 4.000 1939.040 2816.000 1958.040 ;
        RECT 4.000 1937.640 2815.600 1939.040 ;
        RECT 4.000 1928.840 2816.000 1937.640 ;
        RECT 4.400 1927.440 2816.000 1928.840 ;
        RECT 4.000 1908.440 2816.000 1927.440 ;
        RECT 4.000 1907.040 2815.600 1908.440 ;
        RECT 4.000 1894.840 2816.000 1907.040 ;
        RECT 4.400 1893.440 2816.000 1894.840 ;
        RECT 4.000 1874.440 2816.000 1893.440 ;
        RECT 4.000 1873.040 2815.600 1874.440 ;
        RECT 4.000 1860.840 2816.000 1873.040 ;
        RECT 4.400 1859.440 2816.000 1860.840 ;
        RECT 4.000 1840.440 2816.000 1859.440 ;
        RECT 4.000 1839.040 2815.600 1840.440 ;
        RECT 4.000 1826.840 2816.000 1839.040 ;
        RECT 4.400 1825.440 2816.000 1826.840 ;
        RECT 4.000 1806.440 2816.000 1825.440 ;
        RECT 4.000 1805.040 2815.600 1806.440 ;
        RECT 4.000 1792.840 2816.000 1805.040 ;
        RECT 4.400 1791.440 2816.000 1792.840 ;
        RECT 4.000 1775.840 2816.000 1791.440 ;
        RECT 4.000 1774.440 2815.600 1775.840 ;
        RECT 4.000 1762.240 2816.000 1774.440 ;
        RECT 4.400 1760.840 2816.000 1762.240 ;
        RECT 4.000 1741.840 2816.000 1760.840 ;
        RECT 4.000 1740.440 2815.600 1741.840 ;
        RECT 4.000 1728.240 2816.000 1740.440 ;
        RECT 4.400 1726.840 2816.000 1728.240 ;
        RECT 4.000 1707.840 2816.000 1726.840 ;
        RECT 4.000 1706.440 2815.600 1707.840 ;
        RECT 4.000 1694.240 2816.000 1706.440 ;
        RECT 4.400 1692.840 2816.000 1694.240 ;
        RECT 4.000 1673.840 2816.000 1692.840 ;
        RECT 4.000 1672.440 2815.600 1673.840 ;
        RECT 4.000 1660.240 2816.000 1672.440 ;
        RECT 4.400 1658.840 2816.000 1660.240 ;
        RECT 4.000 1639.840 2816.000 1658.840 ;
        RECT 4.000 1638.440 2815.600 1639.840 ;
        RECT 4.000 1629.640 2816.000 1638.440 ;
        RECT 4.400 1628.240 2816.000 1629.640 ;
        RECT 4.000 1609.240 2816.000 1628.240 ;
        RECT 4.000 1607.840 2815.600 1609.240 ;
        RECT 4.000 1595.640 2816.000 1607.840 ;
        RECT 4.400 1594.240 2816.000 1595.640 ;
        RECT 4.000 1575.240 2816.000 1594.240 ;
        RECT 4.000 1573.840 2815.600 1575.240 ;
        RECT 4.000 1561.640 2816.000 1573.840 ;
        RECT 4.400 1560.240 2816.000 1561.640 ;
        RECT 4.000 1541.240 2816.000 1560.240 ;
        RECT 4.000 1539.840 2815.600 1541.240 ;
        RECT 4.000 1527.640 2816.000 1539.840 ;
        RECT 4.400 1526.240 2816.000 1527.640 ;
        RECT 4.000 1507.240 2816.000 1526.240 ;
        RECT 4.000 1505.840 2815.600 1507.240 ;
        RECT 4.000 1493.640 2816.000 1505.840 ;
        RECT 4.400 1492.240 2816.000 1493.640 ;
        RECT 4.000 1476.640 2816.000 1492.240 ;
        RECT 4.000 1475.240 2815.600 1476.640 ;
        RECT 4.000 1463.040 2816.000 1475.240 ;
        RECT 4.400 1461.640 2816.000 1463.040 ;
        RECT 4.000 1442.640 2816.000 1461.640 ;
        RECT 4.000 1441.240 2815.600 1442.640 ;
        RECT 4.000 1429.040 2816.000 1441.240 ;
        RECT 4.400 1427.640 2816.000 1429.040 ;
        RECT 4.000 1408.640 2816.000 1427.640 ;
        RECT 4.000 1407.240 2815.600 1408.640 ;
        RECT 4.000 1395.040 2816.000 1407.240 ;
        RECT 4.400 1393.640 2816.000 1395.040 ;
        RECT 4.000 1374.640 2816.000 1393.640 ;
        RECT 4.000 1373.240 2815.600 1374.640 ;
        RECT 4.000 1361.040 2816.000 1373.240 ;
        RECT 4.400 1359.640 2816.000 1361.040 ;
        RECT 4.000 1340.640 2816.000 1359.640 ;
        RECT 4.000 1339.240 2815.600 1340.640 ;
        RECT 4.000 1330.440 2816.000 1339.240 ;
        RECT 4.400 1329.040 2816.000 1330.440 ;
        RECT 4.000 1310.040 2816.000 1329.040 ;
        RECT 4.000 1308.640 2815.600 1310.040 ;
        RECT 4.000 1296.440 2816.000 1308.640 ;
        RECT 4.400 1295.040 2816.000 1296.440 ;
        RECT 4.000 1276.040 2816.000 1295.040 ;
        RECT 4.000 1274.640 2815.600 1276.040 ;
        RECT 4.000 1262.440 2816.000 1274.640 ;
        RECT 4.400 1261.040 2816.000 1262.440 ;
        RECT 4.000 1242.040 2816.000 1261.040 ;
        RECT 4.000 1240.640 2815.600 1242.040 ;
        RECT 4.000 1228.440 2816.000 1240.640 ;
        RECT 4.400 1227.040 2816.000 1228.440 ;
        RECT 4.000 1208.040 2816.000 1227.040 ;
        RECT 4.000 1206.640 2815.600 1208.040 ;
        RECT 4.000 1194.440 2816.000 1206.640 ;
        RECT 4.400 1193.040 2816.000 1194.440 ;
        RECT 4.000 1177.440 2816.000 1193.040 ;
        RECT 4.000 1176.040 2815.600 1177.440 ;
        RECT 4.000 1163.840 2816.000 1176.040 ;
        RECT 4.400 1162.440 2816.000 1163.840 ;
        RECT 4.000 1143.440 2816.000 1162.440 ;
        RECT 4.000 1142.040 2815.600 1143.440 ;
        RECT 4.000 1129.840 2816.000 1142.040 ;
        RECT 4.400 1128.440 2816.000 1129.840 ;
        RECT 4.000 1109.440 2816.000 1128.440 ;
        RECT 4.000 1108.040 2815.600 1109.440 ;
        RECT 4.000 1095.840 2816.000 1108.040 ;
        RECT 4.400 1094.440 2816.000 1095.840 ;
        RECT 4.000 1075.440 2816.000 1094.440 ;
        RECT 4.000 1074.040 2815.600 1075.440 ;
        RECT 4.000 1061.840 2816.000 1074.040 ;
        RECT 4.400 1060.440 2816.000 1061.840 ;
        RECT 4.000 1041.440 2816.000 1060.440 ;
        RECT 4.000 1040.040 2815.600 1041.440 ;
        RECT 4.000 1031.240 2816.000 1040.040 ;
        RECT 4.400 1029.840 2816.000 1031.240 ;
        RECT 4.000 1010.840 2816.000 1029.840 ;
        RECT 4.000 1009.440 2815.600 1010.840 ;
        RECT 4.000 997.240 2816.000 1009.440 ;
        RECT 4.400 995.840 2816.000 997.240 ;
        RECT 4.000 976.840 2816.000 995.840 ;
        RECT 4.000 975.440 2815.600 976.840 ;
        RECT 4.000 963.240 2816.000 975.440 ;
        RECT 4.400 961.840 2816.000 963.240 ;
        RECT 4.000 942.840 2816.000 961.840 ;
        RECT 4.000 941.440 2815.600 942.840 ;
        RECT 4.000 929.240 2816.000 941.440 ;
        RECT 4.400 927.840 2816.000 929.240 ;
        RECT 4.000 908.840 2816.000 927.840 ;
        RECT 4.000 907.440 2815.600 908.840 ;
        RECT 4.000 895.240 2816.000 907.440 ;
        RECT 4.400 893.840 2816.000 895.240 ;
        RECT 4.000 878.240 2816.000 893.840 ;
        RECT 4.000 876.840 2815.600 878.240 ;
        RECT 4.000 864.640 2816.000 876.840 ;
        RECT 4.400 863.240 2816.000 864.640 ;
        RECT 4.000 844.240 2816.000 863.240 ;
        RECT 4.000 842.840 2815.600 844.240 ;
        RECT 4.000 830.640 2816.000 842.840 ;
        RECT 4.400 829.240 2816.000 830.640 ;
        RECT 4.000 810.240 2816.000 829.240 ;
        RECT 4.000 808.840 2815.600 810.240 ;
        RECT 4.000 796.640 2816.000 808.840 ;
        RECT 4.400 795.240 2816.000 796.640 ;
        RECT 4.000 776.240 2816.000 795.240 ;
        RECT 4.000 774.840 2815.600 776.240 ;
        RECT 4.000 762.640 2816.000 774.840 ;
        RECT 4.400 761.240 2816.000 762.640 ;
        RECT 4.000 742.240 2816.000 761.240 ;
        RECT 4.000 740.840 2815.600 742.240 ;
        RECT 4.000 732.040 2816.000 740.840 ;
        RECT 4.400 730.640 2816.000 732.040 ;
        RECT 4.000 711.640 2816.000 730.640 ;
        RECT 4.000 710.240 2815.600 711.640 ;
        RECT 4.000 698.040 2816.000 710.240 ;
        RECT 4.400 696.640 2816.000 698.040 ;
        RECT 4.000 677.640 2816.000 696.640 ;
        RECT 4.000 676.240 2815.600 677.640 ;
        RECT 4.000 664.040 2816.000 676.240 ;
        RECT 4.400 662.640 2816.000 664.040 ;
        RECT 4.000 643.640 2816.000 662.640 ;
        RECT 4.000 642.240 2815.600 643.640 ;
        RECT 4.000 630.040 2816.000 642.240 ;
        RECT 4.400 628.640 2816.000 630.040 ;
        RECT 4.000 609.640 2816.000 628.640 ;
        RECT 4.000 608.240 2815.600 609.640 ;
        RECT 4.000 596.040 2816.000 608.240 ;
        RECT 4.400 594.640 2816.000 596.040 ;
        RECT 4.000 579.040 2816.000 594.640 ;
        RECT 4.000 577.640 2815.600 579.040 ;
        RECT 4.000 565.440 2816.000 577.640 ;
        RECT 4.400 564.040 2816.000 565.440 ;
        RECT 4.000 545.040 2816.000 564.040 ;
        RECT 4.000 543.640 2815.600 545.040 ;
        RECT 4.000 531.440 2816.000 543.640 ;
        RECT 4.400 530.040 2816.000 531.440 ;
        RECT 4.000 511.040 2816.000 530.040 ;
        RECT 4.000 509.640 2815.600 511.040 ;
        RECT 4.000 497.440 2816.000 509.640 ;
        RECT 4.400 496.040 2816.000 497.440 ;
        RECT 4.000 477.040 2816.000 496.040 ;
        RECT 4.000 475.640 2815.600 477.040 ;
        RECT 4.000 463.440 2816.000 475.640 ;
        RECT 4.400 462.040 2816.000 463.440 ;
        RECT 4.000 443.040 2816.000 462.040 ;
        RECT 4.000 441.640 2815.600 443.040 ;
        RECT 4.000 432.840 2816.000 441.640 ;
        RECT 4.400 431.440 2816.000 432.840 ;
        RECT 4.000 412.440 2816.000 431.440 ;
        RECT 4.000 411.040 2815.600 412.440 ;
        RECT 4.000 398.840 2816.000 411.040 ;
        RECT 4.400 397.440 2816.000 398.840 ;
        RECT 4.000 378.440 2816.000 397.440 ;
        RECT 4.000 377.040 2815.600 378.440 ;
        RECT 4.000 364.840 2816.000 377.040 ;
        RECT 4.400 363.440 2816.000 364.840 ;
        RECT 4.000 344.440 2816.000 363.440 ;
        RECT 4.000 343.040 2815.600 344.440 ;
        RECT 4.000 330.840 2816.000 343.040 ;
        RECT 4.400 329.440 2816.000 330.840 ;
        RECT 4.000 310.440 2816.000 329.440 ;
        RECT 4.000 309.040 2815.600 310.440 ;
        RECT 4.000 296.840 2816.000 309.040 ;
        RECT 4.400 295.440 2816.000 296.840 ;
        RECT 4.000 279.840 2816.000 295.440 ;
        RECT 4.000 278.440 2815.600 279.840 ;
        RECT 4.000 266.240 2816.000 278.440 ;
        RECT 4.400 264.840 2816.000 266.240 ;
        RECT 4.000 245.840 2816.000 264.840 ;
        RECT 4.000 244.440 2815.600 245.840 ;
        RECT 4.000 232.240 2816.000 244.440 ;
        RECT 4.400 230.840 2816.000 232.240 ;
        RECT 4.000 211.840 2816.000 230.840 ;
        RECT 4.000 210.440 2815.600 211.840 ;
        RECT 4.000 198.240 2816.000 210.440 ;
        RECT 4.400 196.840 2816.000 198.240 ;
        RECT 4.000 177.840 2816.000 196.840 ;
        RECT 4.000 176.440 2815.600 177.840 ;
        RECT 4.000 164.240 2816.000 176.440 ;
        RECT 4.400 162.840 2816.000 164.240 ;
        RECT 4.000 147.240 2816.000 162.840 ;
        RECT 4.000 145.840 2815.600 147.240 ;
        RECT 4.000 133.640 2816.000 145.840 ;
        RECT 4.400 132.240 2816.000 133.640 ;
        RECT 4.000 113.240 2816.000 132.240 ;
        RECT 4.000 111.840 2815.600 113.240 ;
        RECT 4.000 99.640 2816.000 111.840 ;
        RECT 4.400 98.240 2816.000 99.640 ;
        RECT 4.000 79.240 2816.000 98.240 ;
        RECT 4.000 77.840 2815.600 79.240 ;
        RECT 4.000 65.640 2816.000 77.840 ;
        RECT 4.400 64.240 2816.000 65.640 ;
        RECT 4.000 45.240 2816.000 64.240 ;
        RECT 4.000 43.840 2815.600 45.240 ;
        RECT 4.000 31.640 2816.000 43.840 ;
        RECT 4.400 30.240 2816.000 31.640 ;
        RECT 4.000 11.240 2816.000 30.240 ;
        RECT 4.000 10.375 2815.600 11.240 ;
      LAYER met4 ;
        RECT 872.455 11.735 942.240 3406.625 ;
        RECT 944.640 11.735 1019.040 3406.625 ;
        RECT 1021.440 11.735 1095.840 3406.625 ;
        RECT 1098.240 11.735 1172.640 3406.625 ;
        RECT 1175.040 11.735 1249.440 3406.625 ;
        RECT 1251.840 11.735 1326.240 3406.625 ;
        RECT 1328.640 11.735 1403.040 3406.625 ;
        RECT 1405.440 11.735 1479.840 3406.625 ;
        RECT 1482.240 11.735 1556.640 3406.625 ;
        RECT 1559.040 11.735 1633.440 3406.625 ;
        RECT 1635.840 11.735 1710.240 3406.625 ;
        RECT 1712.640 11.735 1787.040 3406.625 ;
        RECT 1789.440 11.735 1863.840 3406.625 ;
        RECT 1866.240 11.735 1892.145 3406.625 ;
  END
END RISC_V
END LIBRARY

