magic
tech sky130B
magscale 1 2
timestamp 1663700488
<< obsli1 >>
rect 1104 2159 98808 97393
<< obsm1 >>
rect 14 960 99254 97776
<< metal2 >>
rect 18 99200 74 100000
rect 1950 99200 2006 100000
rect 4526 99200 4582 100000
rect 6458 99200 6514 100000
rect 9034 99200 9090 100000
rect 10966 99200 11022 100000
rect 13542 99200 13598 100000
rect 15474 99200 15530 100000
rect 18050 99200 18106 100000
rect 19982 99200 20038 100000
rect 22558 99200 22614 100000
rect 24490 99200 24546 100000
rect 27066 99200 27122 100000
rect 28998 99200 29054 100000
rect 31574 99200 31630 100000
rect 33506 99200 33562 100000
rect 36082 99200 36138 100000
rect 38014 99200 38070 100000
rect 40590 99200 40646 100000
rect 42522 99200 42578 100000
rect 45098 99200 45154 100000
rect 47030 99200 47086 100000
rect 49606 99200 49662 100000
rect 51538 99200 51594 100000
rect 54114 99200 54170 100000
rect 56046 99200 56102 100000
rect 58622 99200 58678 100000
rect 60554 99200 60610 100000
rect 63130 99200 63186 100000
rect 65062 99200 65118 100000
rect 67638 99200 67694 100000
rect 69570 99200 69626 100000
rect 72146 99200 72202 100000
rect 74078 99200 74134 100000
rect 76654 99200 76710 100000
rect 78586 99200 78642 100000
rect 81162 99200 81218 100000
rect 83094 99200 83150 100000
rect 85670 99200 85726 100000
rect 87602 99200 87658 100000
rect 90178 99200 90234 100000
rect 92110 99200 92166 100000
rect 94686 99200 94742 100000
rect 96618 99200 96674 100000
rect 99194 99200 99250 100000
rect 18 0 74 800
rect 1950 0 2006 800
rect 4526 0 4582 800
rect 6458 0 6514 800
rect 9034 0 9090 800
rect 10966 0 11022 800
rect 13542 0 13598 800
rect 15474 0 15530 800
rect 18050 0 18106 800
rect 19982 0 20038 800
rect 22558 0 22614 800
rect 24490 0 24546 800
rect 27066 0 27122 800
rect 28998 0 29054 800
rect 31574 0 31630 800
rect 33506 0 33562 800
rect 36082 0 36138 800
rect 38014 0 38070 800
rect 40590 0 40646 800
rect 42522 0 42578 800
rect 45098 0 45154 800
rect 47030 0 47086 800
rect 49606 0 49662 800
rect 51538 0 51594 800
rect 54114 0 54170 800
rect 56046 0 56102 800
rect 58622 0 58678 800
rect 60554 0 60610 800
rect 63130 0 63186 800
rect 65062 0 65118 800
rect 67638 0 67694 800
rect 69570 0 69626 800
rect 72146 0 72202 800
rect 74078 0 74134 800
rect 76654 0 76710 800
rect 78586 0 78642 800
rect 81162 0 81218 800
rect 83094 0 83150 800
rect 85670 0 85726 800
rect 87602 0 87658 800
rect 90178 0 90234 800
rect 92110 0 92166 800
rect 94686 0 94742 800
rect 96618 0 96674 800
rect 99194 0 99250 800
<< obsm2 >>
rect 130 99144 1894 99362
rect 2062 99144 4470 99362
rect 4638 99144 6402 99362
rect 6570 99144 8978 99362
rect 9146 99144 10910 99362
rect 11078 99144 13486 99362
rect 13654 99144 15418 99362
rect 15586 99144 17994 99362
rect 18162 99144 19926 99362
rect 20094 99144 22502 99362
rect 22670 99144 24434 99362
rect 24602 99144 27010 99362
rect 27178 99144 28942 99362
rect 29110 99144 31518 99362
rect 31686 99144 33450 99362
rect 33618 99144 36026 99362
rect 36194 99144 37958 99362
rect 38126 99144 40534 99362
rect 40702 99144 42466 99362
rect 42634 99144 45042 99362
rect 45210 99144 46974 99362
rect 47142 99144 49550 99362
rect 49718 99144 51482 99362
rect 51650 99144 54058 99362
rect 54226 99144 55990 99362
rect 56158 99144 58566 99362
rect 58734 99144 60498 99362
rect 60666 99144 63074 99362
rect 63242 99144 65006 99362
rect 65174 99144 67582 99362
rect 67750 99144 69514 99362
rect 69682 99144 72090 99362
rect 72258 99144 74022 99362
rect 74190 99144 76598 99362
rect 76766 99144 78530 99362
rect 78698 99144 81106 99362
rect 81274 99144 83038 99362
rect 83206 99144 85614 99362
rect 85782 99144 87546 99362
rect 87714 99144 90122 99362
rect 90290 99144 92054 99362
rect 92222 99144 94630 99362
rect 94798 99144 96562 99362
rect 96730 99144 99138 99362
rect 20 856 99248 99144
rect 130 711 1894 856
rect 2062 711 4470 856
rect 4638 711 6402 856
rect 6570 711 8978 856
rect 9146 711 10910 856
rect 11078 711 13486 856
rect 13654 711 15418 856
rect 15586 711 17994 856
rect 18162 711 19926 856
rect 20094 711 22502 856
rect 22670 711 24434 856
rect 24602 711 27010 856
rect 27178 711 28942 856
rect 29110 711 31518 856
rect 31686 711 33450 856
rect 33618 711 36026 856
rect 36194 711 37958 856
rect 38126 711 40534 856
rect 40702 711 42466 856
rect 42634 711 45042 856
rect 45210 711 46974 856
rect 47142 711 49550 856
rect 49718 711 51482 856
rect 51650 711 54058 856
rect 54226 711 55990 856
rect 56158 711 58566 856
rect 58734 711 60498 856
rect 60666 711 63074 856
rect 63242 711 65006 856
rect 65174 711 67582 856
rect 67750 711 69514 856
rect 69682 711 72090 856
rect 72258 711 74022 856
rect 74190 711 76598 856
rect 76766 711 78530 856
rect 78698 711 81106 856
rect 81274 711 83038 856
rect 83206 711 85614 856
rect 85782 711 87546 856
rect 87714 711 90122 856
rect 90290 711 92054 856
rect 92222 711 94630 856
rect 94798 711 96562 856
rect 96730 711 99138 856
<< metal3 >>
rect 99200 98608 100000 98728
rect 0 97248 800 97368
rect 99200 95888 100000 96008
rect 0 95208 800 95328
rect 99200 93848 100000 93968
rect 0 92488 800 92608
rect 99200 91128 100000 91248
rect 0 90448 800 90568
rect 99200 89088 100000 89208
rect 0 87728 800 87848
rect 99200 86368 100000 86488
rect 0 85688 800 85808
rect 99200 84328 100000 84448
rect 0 82968 800 83088
rect 99200 81608 100000 81728
rect 0 80928 800 81048
rect 99200 79568 100000 79688
rect 0 78208 800 78328
rect 99200 76848 100000 76968
rect 0 76168 800 76288
rect 99200 74808 100000 74928
rect 0 73448 800 73568
rect 99200 72088 100000 72208
rect 0 71408 800 71528
rect 99200 70048 100000 70168
rect 0 68688 800 68808
rect 99200 67328 100000 67448
rect 0 66648 800 66768
rect 99200 65288 100000 65408
rect 0 63928 800 64048
rect 99200 62568 100000 62688
rect 0 61888 800 62008
rect 99200 60528 100000 60648
rect 0 59168 800 59288
rect 99200 57808 100000 57928
rect 0 57128 800 57248
rect 99200 55768 100000 55888
rect 0 54408 800 54528
rect 99200 53048 100000 53168
rect 0 52368 800 52488
rect 99200 51008 100000 51128
rect 0 49648 800 49768
rect 99200 48288 100000 48408
rect 0 47608 800 47728
rect 99200 46248 100000 46368
rect 0 44888 800 45008
rect 99200 43528 100000 43648
rect 0 42848 800 42968
rect 99200 41488 100000 41608
rect 0 40128 800 40248
rect 99200 38768 100000 38888
rect 0 38088 800 38208
rect 99200 36728 100000 36848
rect 0 35368 800 35488
rect 99200 34008 100000 34128
rect 0 33328 800 33448
rect 99200 31968 100000 32088
rect 0 30608 800 30728
rect 99200 29248 100000 29368
rect 0 28568 800 28688
rect 99200 27208 100000 27328
rect 0 25848 800 25968
rect 99200 24488 100000 24608
rect 0 23808 800 23928
rect 99200 22448 100000 22568
rect 0 21088 800 21208
rect 99200 19728 100000 19848
rect 0 19048 800 19168
rect 99200 17688 100000 17808
rect 0 16328 800 16448
rect 99200 14968 100000 15088
rect 0 14288 800 14408
rect 99200 12928 100000 13048
rect 0 11568 800 11688
rect 99200 10208 100000 10328
rect 0 9528 800 9648
rect 99200 8168 100000 8288
rect 0 6808 800 6928
rect 99200 5448 100000 5568
rect 0 4768 800 4888
rect 99200 3408 100000 3528
rect 0 2048 800 2168
rect 99200 688 100000 808
<< obsm3 >>
rect 790 98528 99120 98701
rect 790 97448 99200 98528
rect 880 97168 99200 97448
rect 790 96088 99200 97168
rect 790 95808 99120 96088
rect 790 95408 99200 95808
rect 880 95128 99200 95408
rect 790 94048 99200 95128
rect 790 93768 99120 94048
rect 790 92688 99200 93768
rect 880 92408 99200 92688
rect 790 91328 99200 92408
rect 790 91048 99120 91328
rect 790 90648 99200 91048
rect 880 90368 99200 90648
rect 790 89288 99200 90368
rect 790 89008 99120 89288
rect 790 87928 99200 89008
rect 880 87648 99200 87928
rect 790 86568 99200 87648
rect 790 86288 99120 86568
rect 790 85888 99200 86288
rect 880 85608 99200 85888
rect 790 84528 99200 85608
rect 790 84248 99120 84528
rect 790 83168 99200 84248
rect 880 82888 99200 83168
rect 790 81808 99200 82888
rect 790 81528 99120 81808
rect 790 81128 99200 81528
rect 880 80848 99200 81128
rect 790 79768 99200 80848
rect 790 79488 99120 79768
rect 790 78408 99200 79488
rect 880 78128 99200 78408
rect 790 77048 99200 78128
rect 790 76768 99120 77048
rect 790 76368 99200 76768
rect 880 76088 99200 76368
rect 790 75008 99200 76088
rect 790 74728 99120 75008
rect 790 73648 99200 74728
rect 880 73368 99200 73648
rect 790 72288 99200 73368
rect 790 72008 99120 72288
rect 790 71608 99200 72008
rect 880 71328 99200 71608
rect 790 70248 99200 71328
rect 790 69968 99120 70248
rect 790 68888 99200 69968
rect 880 68608 99200 68888
rect 790 67528 99200 68608
rect 790 67248 99120 67528
rect 790 66848 99200 67248
rect 880 66568 99200 66848
rect 790 65488 99200 66568
rect 790 65208 99120 65488
rect 790 64128 99200 65208
rect 880 63848 99200 64128
rect 790 62768 99200 63848
rect 790 62488 99120 62768
rect 790 62088 99200 62488
rect 880 61808 99200 62088
rect 790 60728 99200 61808
rect 790 60448 99120 60728
rect 790 59368 99200 60448
rect 880 59088 99200 59368
rect 790 58008 99200 59088
rect 790 57728 99120 58008
rect 790 57328 99200 57728
rect 880 57048 99200 57328
rect 790 55968 99200 57048
rect 790 55688 99120 55968
rect 790 54608 99200 55688
rect 880 54328 99200 54608
rect 790 53248 99200 54328
rect 790 52968 99120 53248
rect 790 52568 99200 52968
rect 880 52288 99200 52568
rect 790 51208 99200 52288
rect 790 50928 99120 51208
rect 790 49848 99200 50928
rect 880 49568 99200 49848
rect 790 48488 99200 49568
rect 790 48208 99120 48488
rect 790 47808 99200 48208
rect 880 47528 99200 47808
rect 790 46448 99200 47528
rect 790 46168 99120 46448
rect 790 45088 99200 46168
rect 880 44808 99200 45088
rect 790 43728 99200 44808
rect 790 43448 99120 43728
rect 790 43048 99200 43448
rect 880 42768 99200 43048
rect 790 41688 99200 42768
rect 790 41408 99120 41688
rect 790 40328 99200 41408
rect 880 40048 99200 40328
rect 790 38968 99200 40048
rect 790 38688 99120 38968
rect 790 38288 99200 38688
rect 880 38008 99200 38288
rect 790 36928 99200 38008
rect 790 36648 99120 36928
rect 790 35568 99200 36648
rect 880 35288 99200 35568
rect 790 34208 99200 35288
rect 790 33928 99120 34208
rect 790 33528 99200 33928
rect 880 33248 99200 33528
rect 790 32168 99200 33248
rect 790 31888 99120 32168
rect 790 30808 99200 31888
rect 880 30528 99200 30808
rect 790 29448 99200 30528
rect 790 29168 99120 29448
rect 790 28768 99200 29168
rect 880 28488 99200 28768
rect 790 27408 99200 28488
rect 790 27128 99120 27408
rect 790 26048 99200 27128
rect 880 25768 99200 26048
rect 790 24688 99200 25768
rect 790 24408 99120 24688
rect 790 24008 99200 24408
rect 880 23728 99200 24008
rect 790 22648 99200 23728
rect 790 22368 99120 22648
rect 790 21288 99200 22368
rect 880 21008 99200 21288
rect 790 19928 99200 21008
rect 790 19648 99120 19928
rect 790 19248 99200 19648
rect 880 18968 99200 19248
rect 790 17888 99200 18968
rect 790 17608 99120 17888
rect 790 16528 99200 17608
rect 880 16248 99200 16528
rect 790 15168 99200 16248
rect 790 14888 99120 15168
rect 790 14488 99200 14888
rect 880 14208 99200 14488
rect 790 13128 99200 14208
rect 790 12848 99120 13128
rect 790 11768 99200 12848
rect 880 11488 99200 11768
rect 790 10408 99200 11488
rect 790 10128 99120 10408
rect 790 9728 99200 10128
rect 880 9448 99200 9728
rect 790 8368 99200 9448
rect 790 8088 99120 8368
rect 790 7008 99200 8088
rect 880 6728 99200 7008
rect 790 5648 99200 6728
rect 790 5368 99120 5648
rect 790 4968 99200 5368
rect 880 4688 99200 4968
rect 790 3608 99200 4688
rect 790 3328 99120 3608
rect 790 2248 99200 3328
rect 880 1968 99200 2248
rect 790 888 99200 1968
rect 790 715 99120 888
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
<< obsm4 >>
rect 795 97504 92309 97613
rect 795 2048 4128 97504
rect 4608 2048 19488 97504
rect 19968 2048 34848 97504
rect 35328 2048 50208 97504
rect 50688 2048 65568 97504
rect 66048 2048 80928 97504
rect 81408 2048 92309 97504
rect 795 987 92309 2048
<< labels >>
rlabel metal2 s 96618 99200 96674 100000 6 clk
port 1 nsew signal input
rlabel metal2 s 40590 99200 40646 100000 6 funct3[0]
port 2 nsew signal output
rlabel metal3 s 99200 12928 100000 13048 6 funct3[1]
port 3 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 funct3[2]
port 4 nsew signal output
rlabel metal3 s 0 80928 800 81048 6 funct7[0]
port 5 nsew signal output
rlabel metal2 s 13542 99200 13598 100000 6 funct7[1]
port 6 nsew signal output
rlabel metal3 s 0 57128 800 57248 6 funct7[2]
port 7 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 funct7[3]
port 8 nsew signal output
rlabel metal2 s 81162 0 81218 800 6 funct7[4]
port 9 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 funct7[5]
port 10 nsew signal output
rlabel metal3 s 99200 93848 100000 93968 6 funct7[6]
port 11 nsew signal output
rlabel metal2 s 65062 99200 65118 100000 6 immediate[0]
port 12 nsew signal output
rlabel metal2 s 60554 99200 60610 100000 6 immediate[10]
port 13 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 immediate[11]
port 14 nsew signal output
rlabel metal2 s 47030 99200 47086 100000 6 immediate[12]
port 15 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 immediate[13]
port 16 nsew signal output
rlabel metal2 s 9034 99200 9090 100000 6 immediate[14]
port 17 nsew signal output
rlabel metal2 s 18 99200 74 100000 6 immediate[15]
port 18 nsew signal output
rlabel metal2 s 58622 99200 58678 100000 6 immediate[16]
port 19 nsew signal output
rlabel metal3 s 99200 14968 100000 15088 6 immediate[17]
port 20 nsew signal output
rlabel metal2 s 22558 99200 22614 100000 6 immediate[18]
port 21 nsew signal output
rlabel metal2 s 45098 99200 45154 100000 6 immediate[19]
port 22 nsew signal output
rlabel metal3 s 99200 43528 100000 43648 6 immediate[1]
port 23 nsew signal output
rlabel metal2 s 24490 99200 24546 100000 6 immediate[20]
port 24 nsew signal output
rlabel metal3 s 99200 89088 100000 89208 6 immediate[21]
port 25 nsew signal output
rlabel metal3 s 99200 8168 100000 8288 6 immediate[22]
port 26 nsew signal output
rlabel metal2 s 76654 99200 76710 100000 6 immediate[23]
port 27 nsew signal output
rlabel metal3 s 99200 5448 100000 5568 6 immediate[24]
port 28 nsew signal output
rlabel metal2 s 78586 0 78642 800 6 immediate[25]
port 29 nsew signal output
rlabel metal3 s 0 52368 800 52488 6 immediate[26]
port 30 nsew signal output
rlabel metal2 s 6458 99200 6514 100000 6 immediate[27]
port 31 nsew signal output
rlabel metal3 s 0 61888 800 62008 6 immediate[28]
port 32 nsew signal output
rlabel metal3 s 99200 84328 100000 84448 6 immediate[29]
port 33 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 immediate[2]
port 34 nsew signal output
rlabel metal2 s 19982 99200 20038 100000 6 immediate[30]
port 35 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 immediate[31]
port 36 nsew signal output
rlabel metal2 s 90178 99200 90234 100000 6 immediate[3]
port 37 nsew signal output
rlabel metal2 s 4526 99200 4582 100000 6 immediate[4]
port 38 nsew signal output
rlabel metal2 s 31574 99200 31630 100000 6 immediate[5]
port 39 nsew signal output
rlabel metal3 s 99200 79568 100000 79688 6 immediate[6]
port 40 nsew signal output
rlabel metal3 s 99200 62568 100000 62688 6 immediate[7]
port 41 nsew signal output
rlabel metal3 s 99200 41488 100000 41608 6 immediate[8]
port 42 nsew signal output
rlabel metal2 s 81162 99200 81218 100000 6 immediate[9]
port 43 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 instruction_type_output[0]
port 44 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 instruction_type_output[1]
port 45 nsew signal output
rlabel metal2 s 99194 0 99250 800 6 instruction_type_output[2]
port 46 nsew signal output
rlabel metal3 s 99200 76848 100000 76968 6 instruction_type_output[3]
port 47 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 instruction_type_output[4]
port 48 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 instruction_type_output[5]
port 49 nsew signal output
rlabel metal3 s 99200 53048 100000 53168 6 la_instruction_input[0]
port 50 nsew signal input
rlabel metal2 s 94686 99200 94742 100000 6 la_instruction_input[10]
port 51 nsew signal input
rlabel metal2 s 42522 99200 42578 100000 6 la_instruction_input[11]
port 52 nsew signal input
rlabel metal3 s 99200 48288 100000 48408 6 la_instruction_input[12]
port 53 nsew signal input
rlabel metal2 s 92110 99200 92166 100000 6 la_instruction_input[13]
port 54 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 la_instruction_input[14]
port 55 nsew signal input
rlabel metal3 s 99200 19728 100000 19848 6 la_instruction_input[15]
port 56 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 la_instruction_input[16]
port 57 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 la_instruction_input[17]
port 58 nsew signal input
rlabel metal2 s 87602 99200 87658 100000 6 la_instruction_input[18]
port 59 nsew signal input
rlabel metal3 s 99200 98608 100000 98728 6 la_instruction_input[19]
port 60 nsew signal input
rlabel metal2 s 38014 99200 38070 100000 6 la_instruction_input[1]
port 61 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 la_instruction_input[20]
port 62 nsew signal input
rlabel metal2 s 63130 99200 63186 100000 6 la_instruction_input[21]
port 63 nsew signal input
rlabel metal2 s 10966 99200 11022 100000 6 la_instruction_input[22]
port 64 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 la_instruction_input[23]
port 65 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 la_instruction_input[24]
port 66 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 la_instruction_input[25]
port 67 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 la_instruction_input[26]
port 68 nsew signal input
rlabel metal2 s 85670 99200 85726 100000 6 la_instruction_input[27]
port 69 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 la_instruction_input[28]
port 70 nsew signal input
rlabel metal3 s 99200 24488 100000 24608 6 la_instruction_input[29]
port 71 nsew signal input
rlabel metal3 s 99200 36728 100000 36848 6 la_instruction_input[2]
port 72 nsew signal input
rlabel metal3 s 0 95208 800 95328 6 la_instruction_input[30]
port 73 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 la_instruction_input[31]
port 74 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 la_instruction_input[3]
port 75 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_instruction_input[4]
port 76 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 la_instruction_input[5]
port 77 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 la_instruction_input[6]
port 78 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 la_instruction_input[7]
port 79 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 la_instruction_input[8]
port 80 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 la_instruction_input[9]
port 81 nsew signal input
rlabel metal2 s 28998 99200 29054 100000 6 la_instruction_read[0]
port 82 nsew signal output
rlabel metal2 s 36082 99200 36138 100000 6 la_instruction_read[10]
port 83 nsew signal output
rlabel metal3 s 0 76168 800 76288 6 la_instruction_read[11]
port 84 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 la_instruction_read[12]
port 85 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 la_instruction_read[13]
port 86 nsew signal output
rlabel metal3 s 99200 81608 100000 81728 6 la_instruction_read[14]
port 87 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 la_instruction_read[15]
port 88 nsew signal output
rlabel metal3 s 0 90448 800 90568 6 la_instruction_read[16]
port 89 nsew signal output
rlabel metal3 s 99200 70048 100000 70168 6 la_instruction_read[17]
port 90 nsew signal output
rlabel metal2 s 27066 99200 27122 100000 6 la_instruction_read[18]
port 91 nsew signal output
rlabel metal3 s 99200 27208 100000 27328 6 la_instruction_read[19]
port 92 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 la_instruction_read[1]
port 93 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 la_instruction_read[20]
port 94 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 la_instruction_read[21]
port 95 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 la_instruction_read[22]
port 96 nsew signal output
rlabel metal3 s 99200 51008 100000 51128 6 la_instruction_read[23]
port 97 nsew signal output
rlabel metal3 s 0 42848 800 42968 6 la_instruction_read[24]
port 98 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 la_instruction_read[25]
port 99 nsew signal output
rlabel metal2 s 54114 99200 54170 100000 6 la_instruction_read[26]
port 100 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 la_instruction_read[27]
port 101 nsew signal output
rlabel metal3 s 0 92488 800 92608 6 la_instruction_read[28]
port 102 nsew signal output
rlabel metal3 s 99200 91128 100000 91248 6 la_instruction_read[29]
port 103 nsew signal output
rlabel metal3 s 99200 31968 100000 32088 6 la_instruction_read[2]
port 104 nsew signal output
rlabel metal2 s 56046 99200 56102 100000 6 la_instruction_read[30]
port 105 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 la_instruction_read[31]
port 106 nsew signal output
rlabel metal2 s 67638 99200 67694 100000 6 la_instruction_read[3]
port 107 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 la_instruction_read[4]
port 108 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 la_instruction_read[5]
port 109 nsew signal output
rlabel metal3 s 99200 10208 100000 10328 6 la_instruction_read[6]
port 110 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 la_instruction_read[7]
port 111 nsew signal output
rlabel metal3 s 99200 74808 100000 74928 6 la_instruction_read[8]
port 112 nsew signal output
rlabel metal3 s 99200 55768 100000 55888 6 la_instruction_read[9]
port 113 nsew signal output
rlabel metal2 s 74078 99200 74134 100000 6 la_instruction_select[0]
port 114 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 la_instruction_select[1]
port 115 nsew signal input
rlabel metal3 s 99200 22448 100000 22568 6 la_instruction_select[2]
port 116 nsew signal input
rlabel metal3 s 99200 57808 100000 57928 6 la_instruction_select[3]
port 117 nsew signal input
rlabel metal2 s 33506 99200 33562 100000 6 la_instruction_write
port 118 nsew signal input
rlabel metal3 s 99200 38768 100000 38888 6 opcode[0]
port 119 nsew signal output
rlabel metal3 s 99200 688 100000 808 6 opcode[1]
port 120 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 opcode[2]
port 121 nsew signal output
rlabel metal3 s 99200 72088 100000 72208 6 opcode[3]
port 122 nsew signal output
rlabel metal2 s 78586 99200 78642 100000 6 opcode[4]
port 123 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 opcode[5]
port 124 nsew signal output
rlabel metal3 s 99200 29248 100000 29368 6 opcode[6]
port 125 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 pc[0]
port 126 nsew signal input
rlabel metal3 s 99200 3408 100000 3528 6 pc[10]
port 127 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 pc[11]
port 128 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 pc[12]
port 129 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 pc[13]
port 130 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 pc[14]
port 131 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 pc[15]
port 132 nsew signal input
rlabel metal3 s 99200 86368 100000 86488 6 pc[16]
port 133 nsew signal input
rlabel metal3 s 99200 60528 100000 60648 6 pc[17]
port 134 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 pc[18]
port 135 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 pc[19]
port 136 nsew signal input
rlabel metal3 s 99200 34008 100000 34128 6 pc[1]
port 137 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 pc[20]
port 138 nsew signal input
rlabel metal3 s 99200 65288 100000 65408 6 pc[21]
port 139 nsew signal input
rlabel metal3 s 99200 95888 100000 96008 6 pc[22]
port 140 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 pc[23]
port 141 nsew signal input
rlabel metal2 s 99194 99200 99250 100000 6 pc[24]
port 142 nsew signal input
rlabel metal3 s 0 68688 800 68808 6 pc[25]
port 143 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 pc[26]
port 144 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 pc[27]
port 145 nsew signal input
rlabel metal2 s 18 0 74 800 6 pc[28]
port 146 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 pc[29]
port 147 nsew signal input
rlabel metal3 s 0 82968 800 83088 6 pc[2]
port 148 nsew signal input
rlabel metal2 s 15474 99200 15530 100000 6 pc[30]
port 149 nsew signal input
rlabel metal2 s 51538 99200 51594 100000 6 pc[31]
port 150 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 pc[3]
port 151 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 pc[4]
port 152 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 pc[5]
port 153 nsew signal input
rlabel metal2 s 69570 99200 69626 100000 6 pc[6]
port 154 nsew signal input
rlabel metal2 s 49606 99200 49662 100000 6 pc[7]
port 155 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 pc[8]
port 156 nsew signal input
rlabel metal2 s 83094 99200 83150 100000 6 pc[9]
port 157 nsew signal input
rlabel metal3 s 99200 17688 100000 17808 6 rd[0]
port 158 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 rd[1]
port 159 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 rd[2]
port 160 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 rd[3]
port 161 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 rd[4]
port 162 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 rs1[0]
port 163 nsew signal output
rlabel metal3 s 99200 67328 100000 67448 6 rs1[1]
port 164 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 rs1[2]
port 165 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 rs1[3]
port 166 nsew signal output
rlabel metal2 s 72146 99200 72202 100000 6 rs1[4]
port 167 nsew signal output
rlabel metal2 s 1950 99200 2006 100000 6 rs2[0]
port 168 nsew signal output
rlabel metal2 s 18050 99200 18106 100000 6 rs2[1]
port 169 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 rs2[2]
port 170 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 rs2[3]
port 171 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 rs2[4]
port 172 nsew signal output
rlabel metal3 s 99200 46248 100000 46368 6 rst_n
port 173 nsew signal input
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 174 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 174 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 174 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 174 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 175 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 175 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 175 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 15633532
string GDS_FILE /home/drewarosa/RISC-V-Single-Cycle-CPU-Core/openlane/IMemory/runs/22_09_20_14_56/results/signoff/IMemory.magic.gds
string GDS_START 601638
<< end >>

