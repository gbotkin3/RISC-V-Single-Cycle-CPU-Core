magic
tech sky130B
magscale 1 2
timestamp 1663853063
<< nwell >>
rect 1066 148229 147790 148550
rect 1066 147141 147790 147707
rect 1066 146053 147790 146619
rect 1066 144965 147790 145531
rect 1066 143877 147790 144443
rect 1066 142789 147790 143355
rect 1066 141701 147790 142267
rect 1066 140613 147790 141179
rect 1066 139525 147790 140091
rect 1066 138437 147790 139003
rect 1066 137349 147790 137915
rect 1066 136261 147790 136827
rect 1066 135173 147790 135739
rect 1066 134085 147790 134651
rect 1066 132997 147790 133563
rect 1066 131909 147790 132475
rect 1066 130821 147790 131387
rect 1066 129733 147790 130299
rect 1066 128645 147790 129211
rect 1066 127557 147790 128123
rect 1066 126469 147790 127035
rect 1066 125381 147790 125947
rect 1066 124293 147790 124859
rect 1066 123205 147790 123771
rect 1066 122117 147790 122683
rect 1066 121029 147790 121595
rect 1066 119941 147790 120507
rect 1066 118853 147790 119419
rect 1066 117765 147790 118331
rect 1066 116677 147790 117243
rect 1066 115589 147790 116155
rect 1066 114501 147790 115067
rect 1066 113413 147790 113979
rect 1066 112325 147790 112891
rect 1066 111237 147790 111803
rect 1066 110149 147790 110715
rect 1066 109061 147790 109627
rect 1066 107973 147790 108539
rect 1066 106885 147790 107451
rect 1066 105797 147790 106363
rect 1066 104709 147790 105275
rect 1066 103621 147790 104187
rect 1066 102533 147790 103099
rect 1066 101445 147790 102011
rect 1066 100357 147790 100923
rect 1066 99269 147790 99835
rect 1066 98181 147790 98747
rect 1066 97093 147790 97659
rect 1066 96005 147790 96571
rect 1066 94917 147790 95483
rect 1066 93829 147790 94395
rect 1066 92741 147790 93307
rect 1066 91653 147790 92219
rect 1066 90565 147790 91131
rect 1066 89477 147790 90043
rect 1066 88389 147790 88955
rect 1066 87301 147790 87867
rect 1066 86213 147790 86779
rect 1066 85125 147790 85691
rect 1066 84037 147790 84603
rect 1066 82949 147790 83515
rect 1066 81861 147790 82427
rect 1066 80773 147790 81339
rect 1066 79685 147790 80251
rect 1066 78597 147790 79163
rect 1066 77509 147790 78075
rect 1066 76421 147790 76987
rect 1066 75333 147790 75899
rect 1066 74245 147790 74811
rect 1066 73157 147790 73723
rect 1066 72069 147790 72635
rect 1066 70981 147790 71547
rect 1066 69893 147790 70459
rect 1066 68805 147790 69371
rect 1066 67717 147790 68283
rect 1066 66629 147790 67195
rect 1066 65541 147790 66107
rect 1066 64453 147790 65019
rect 1066 63365 147790 63931
rect 1066 62277 147790 62843
rect 1066 61189 147790 61755
rect 1066 60101 147790 60667
rect 1066 59013 147790 59579
rect 1066 57925 147790 58491
rect 1066 56837 147790 57403
rect 1066 55749 147790 56315
rect 1066 54661 147790 55227
rect 1066 53573 147790 54139
rect 1066 52485 147790 53051
rect 1066 51397 147790 51963
rect 1066 50309 147790 50875
rect 1066 49221 147790 49787
rect 1066 48133 147790 48699
rect 1066 47045 147790 47611
rect 1066 45957 147790 46523
rect 1066 44869 147790 45435
rect 1066 43781 147790 44347
rect 1066 42693 147790 43259
rect 1066 41605 147790 42171
rect 1066 40517 147790 41083
rect 1066 39429 147790 39995
rect 1066 38341 147790 38907
rect 1066 37253 147790 37819
rect 1066 36165 147790 36731
rect 1066 35077 147790 35643
rect 1066 33989 147790 34555
rect 1066 32901 147790 33467
rect 1066 31813 147790 32379
rect 1066 30725 147790 31291
rect 1066 29637 147790 30203
rect 1066 28549 147790 29115
rect 1066 27461 147790 28027
rect 1066 26373 147790 26939
rect 1066 25285 147790 25851
rect 1066 24197 147790 24763
rect 1066 23109 147790 23675
rect 1066 22021 147790 22587
rect 1066 20933 147790 21499
rect 1066 19845 147790 20411
rect 1066 18757 147790 19323
rect 1066 17669 147790 18235
rect 1066 16581 147790 17147
rect 1066 15493 147790 16059
rect 1066 14405 147790 14971
rect 1066 13317 147790 13883
rect 1066 12229 147790 12795
rect 1066 11141 147790 11707
rect 1066 10053 147790 10619
rect 1066 8965 147790 9531
rect 1066 7877 147790 8443
rect 1066 6789 147790 7355
rect 1066 5701 147790 6267
rect 1066 4613 147790 5179
rect 1066 3525 147790 4091
rect 1066 2437 147790 3003
<< obsli1 >>
rect 1104 2159 147752 148529
<< obsm1 >>
rect 1104 348 148566 150272
<< metal2 >>
rect 3790 0 3846 800
rect 4158 0 4214 800
rect 4526 0 4582 800
rect 4894 0 4950 800
rect 5262 0 5318 800
rect 5630 0 5686 800
rect 5998 0 6054 800
rect 6366 0 6422 800
rect 6734 0 6790 800
rect 7102 0 7158 800
rect 7470 0 7526 800
rect 7838 0 7894 800
rect 8206 0 8262 800
rect 8574 0 8630 800
rect 8942 0 8998 800
rect 9310 0 9366 800
rect 9678 0 9734 800
rect 10046 0 10102 800
rect 10414 0 10470 800
rect 10782 0 10838 800
rect 11150 0 11206 800
rect 11518 0 11574 800
rect 11886 0 11942 800
rect 12254 0 12310 800
rect 12622 0 12678 800
rect 12990 0 13046 800
rect 13358 0 13414 800
rect 13726 0 13782 800
rect 14094 0 14150 800
rect 14462 0 14518 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15566 0 15622 800
rect 15934 0 15990 800
rect 16302 0 16358 800
rect 16670 0 16726 800
rect 17038 0 17094 800
rect 17406 0 17462 800
rect 17774 0 17830 800
rect 18142 0 18198 800
rect 18510 0 18566 800
rect 18878 0 18934 800
rect 19246 0 19302 800
rect 19614 0 19670 800
rect 19982 0 20038 800
rect 20350 0 20406 800
rect 20718 0 20774 800
rect 21086 0 21142 800
rect 21454 0 21510 800
rect 21822 0 21878 800
rect 22190 0 22246 800
rect 22558 0 22614 800
rect 22926 0 22982 800
rect 23294 0 23350 800
rect 23662 0 23718 800
rect 24030 0 24086 800
rect 24398 0 24454 800
rect 24766 0 24822 800
rect 25134 0 25190 800
rect 25502 0 25558 800
rect 25870 0 25926 800
rect 26238 0 26294 800
rect 26606 0 26662 800
rect 26974 0 27030 800
rect 27342 0 27398 800
rect 27710 0 27766 800
rect 28078 0 28134 800
rect 28446 0 28502 800
rect 28814 0 28870 800
rect 29182 0 29238 800
rect 29550 0 29606 800
rect 29918 0 29974 800
rect 30286 0 30342 800
rect 30654 0 30710 800
rect 31022 0 31078 800
rect 31390 0 31446 800
rect 31758 0 31814 800
rect 32126 0 32182 800
rect 32494 0 32550 800
rect 32862 0 32918 800
rect 33230 0 33286 800
rect 33598 0 33654 800
rect 33966 0 34022 800
rect 34334 0 34390 800
rect 34702 0 34758 800
rect 35070 0 35126 800
rect 35438 0 35494 800
rect 35806 0 35862 800
rect 36174 0 36230 800
rect 36542 0 36598 800
rect 36910 0 36966 800
rect 37278 0 37334 800
rect 37646 0 37702 800
rect 38014 0 38070 800
rect 38382 0 38438 800
rect 38750 0 38806 800
rect 39118 0 39174 800
rect 39486 0 39542 800
rect 39854 0 39910 800
rect 40222 0 40278 800
rect 40590 0 40646 800
rect 40958 0 41014 800
rect 41326 0 41382 800
rect 41694 0 41750 800
rect 42062 0 42118 800
rect 42430 0 42486 800
rect 42798 0 42854 800
rect 43166 0 43222 800
rect 43534 0 43590 800
rect 43902 0 43958 800
rect 44270 0 44326 800
rect 44638 0 44694 800
rect 45006 0 45062 800
rect 45374 0 45430 800
rect 45742 0 45798 800
rect 46110 0 46166 800
rect 46478 0 46534 800
rect 46846 0 46902 800
rect 47214 0 47270 800
rect 47582 0 47638 800
rect 47950 0 48006 800
rect 48318 0 48374 800
rect 48686 0 48742 800
rect 49054 0 49110 800
rect 49422 0 49478 800
rect 49790 0 49846 800
rect 50158 0 50214 800
rect 50526 0 50582 800
rect 50894 0 50950 800
rect 51262 0 51318 800
rect 51630 0 51686 800
rect 51998 0 52054 800
rect 52366 0 52422 800
rect 52734 0 52790 800
rect 53102 0 53158 800
rect 53470 0 53526 800
rect 53838 0 53894 800
rect 54206 0 54262 800
rect 54574 0 54630 800
rect 54942 0 54998 800
rect 55310 0 55366 800
rect 55678 0 55734 800
rect 56046 0 56102 800
rect 56414 0 56470 800
rect 56782 0 56838 800
rect 57150 0 57206 800
rect 57518 0 57574 800
rect 57886 0 57942 800
rect 58254 0 58310 800
rect 58622 0 58678 800
rect 58990 0 59046 800
rect 59358 0 59414 800
rect 59726 0 59782 800
rect 60094 0 60150 800
rect 60462 0 60518 800
rect 60830 0 60886 800
rect 61198 0 61254 800
rect 61566 0 61622 800
rect 61934 0 61990 800
rect 62302 0 62358 800
rect 62670 0 62726 800
rect 63038 0 63094 800
rect 63406 0 63462 800
rect 63774 0 63830 800
rect 64142 0 64198 800
rect 64510 0 64566 800
rect 64878 0 64934 800
rect 65246 0 65302 800
rect 65614 0 65670 800
rect 65982 0 66038 800
rect 66350 0 66406 800
rect 66718 0 66774 800
rect 67086 0 67142 800
rect 67454 0 67510 800
rect 67822 0 67878 800
rect 68190 0 68246 800
rect 68558 0 68614 800
rect 68926 0 68982 800
rect 69294 0 69350 800
rect 69662 0 69718 800
rect 70030 0 70086 800
rect 70398 0 70454 800
rect 70766 0 70822 800
rect 71134 0 71190 800
rect 71502 0 71558 800
rect 71870 0 71926 800
rect 72238 0 72294 800
rect 72606 0 72662 800
rect 72974 0 73030 800
rect 73342 0 73398 800
rect 73710 0 73766 800
rect 74078 0 74134 800
rect 74446 0 74502 800
rect 74814 0 74870 800
rect 75182 0 75238 800
rect 75550 0 75606 800
rect 75918 0 75974 800
rect 76286 0 76342 800
rect 76654 0 76710 800
rect 77022 0 77078 800
rect 77390 0 77446 800
rect 77758 0 77814 800
rect 78126 0 78182 800
rect 78494 0 78550 800
rect 78862 0 78918 800
rect 79230 0 79286 800
rect 79598 0 79654 800
rect 79966 0 80022 800
rect 80334 0 80390 800
rect 80702 0 80758 800
rect 81070 0 81126 800
rect 81438 0 81494 800
rect 81806 0 81862 800
rect 82174 0 82230 800
rect 82542 0 82598 800
rect 82910 0 82966 800
rect 83278 0 83334 800
rect 83646 0 83702 800
rect 84014 0 84070 800
rect 84382 0 84438 800
rect 84750 0 84806 800
rect 85118 0 85174 800
rect 85486 0 85542 800
rect 85854 0 85910 800
rect 86222 0 86278 800
rect 86590 0 86646 800
rect 86958 0 87014 800
rect 87326 0 87382 800
rect 87694 0 87750 800
rect 88062 0 88118 800
rect 88430 0 88486 800
rect 88798 0 88854 800
rect 89166 0 89222 800
rect 89534 0 89590 800
rect 89902 0 89958 800
rect 90270 0 90326 800
rect 90638 0 90694 800
rect 91006 0 91062 800
rect 91374 0 91430 800
rect 91742 0 91798 800
rect 92110 0 92166 800
rect 92478 0 92534 800
rect 92846 0 92902 800
rect 93214 0 93270 800
rect 93582 0 93638 800
rect 93950 0 94006 800
rect 94318 0 94374 800
rect 94686 0 94742 800
rect 95054 0 95110 800
rect 95422 0 95478 800
rect 95790 0 95846 800
rect 96158 0 96214 800
rect 96526 0 96582 800
rect 96894 0 96950 800
rect 97262 0 97318 800
rect 97630 0 97686 800
rect 97998 0 98054 800
rect 98366 0 98422 800
rect 98734 0 98790 800
rect 99102 0 99158 800
rect 99470 0 99526 800
rect 99838 0 99894 800
rect 100206 0 100262 800
rect 100574 0 100630 800
rect 100942 0 100998 800
rect 101310 0 101366 800
rect 101678 0 101734 800
rect 102046 0 102102 800
rect 102414 0 102470 800
rect 102782 0 102838 800
rect 103150 0 103206 800
rect 103518 0 103574 800
rect 103886 0 103942 800
rect 104254 0 104310 800
rect 104622 0 104678 800
rect 104990 0 105046 800
rect 105358 0 105414 800
rect 105726 0 105782 800
rect 106094 0 106150 800
rect 106462 0 106518 800
rect 106830 0 106886 800
rect 107198 0 107254 800
rect 107566 0 107622 800
rect 107934 0 107990 800
rect 108302 0 108358 800
rect 108670 0 108726 800
rect 109038 0 109094 800
rect 109406 0 109462 800
rect 109774 0 109830 800
rect 110142 0 110198 800
rect 110510 0 110566 800
rect 110878 0 110934 800
rect 111246 0 111302 800
rect 111614 0 111670 800
rect 111982 0 112038 800
rect 112350 0 112406 800
rect 112718 0 112774 800
rect 113086 0 113142 800
rect 113454 0 113510 800
rect 113822 0 113878 800
rect 114190 0 114246 800
rect 114558 0 114614 800
rect 114926 0 114982 800
rect 115294 0 115350 800
rect 115662 0 115718 800
rect 116030 0 116086 800
rect 116398 0 116454 800
rect 116766 0 116822 800
rect 117134 0 117190 800
rect 117502 0 117558 800
rect 117870 0 117926 800
rect 118238 0 118294 800
rect 118606 0 118662 800
rect 118974 0 119030 800
rect 119342 0 119398 800
rect 119710 0 119766 800
rect 120078 0 120134 800
rect 120446 0 120502 800
rect 120814 0 120870 800
rect 121182 0 121238 800
rect 121550 0 121606 800
rect 121918 0 121974 800
rect 122286 0 122342 800
rect 122654 0 122710 800
rect 123022 0 123078 800
rect 123390 0 123446 800
rect 123758 0 123814 800
rect 124126 0 124182 800
rect 124494 0 124550 800
rect 124862 0 124918 800
rect 125230 0 125286 800
rect 125598 0 125654 800
rect 125966 0 126022 800
rect 126334 0 126390 800
rect 126702 0 126758 800
rect 127070 0 127126 800
rect 127438 0 127494 800
rect 127806 0 127862 800
rect 128174 0 128230 800
rect 128542 0 128598 800
rect 128910 0 128966 800
rect 129278 0 129334 800
rect 129646 0 129702 800
rect 130014 0 130070 800
rect 130382 0 130438 800
rect 130750 0 130806 800
rect 131118 0 131174 800
rect 131486 0 131542 800
rect 131854 0 131910 800
rect 132222 0 132278 800
rect 132590 0 132646 800
rect 132958 0 133014 800
rect 133326 0 133382 800
rect 133694 0 133750 800
rect 134062 0 134118 800
rect 134430 0 134486 800
rect 134798 0 134854 800
rect 135166 0 135222 800
rect 135534 0 135590 800
rect 135902 0 135958 800
rect 136270 0 136326 800
rect 136638 0 136694 800
rect 137006 0 137062 800
rect 137374 0 137430 800
rect 137742 0 137798 800
rect 138110 0 138166 800
rect 138478 0 138534 800
rect 138846 0 138902 800
rect 139214 0 139270 800
rect 139582 0 139638 800
rect 139950 0 140006 800
rect 140318 0 140374 800
rect 140686 0 140742 800
rect 141054 0 141110 800
rect 141422 0 141478 800
rect 141790 0 141846 800
rect 142158 0 142214 800
rect 142526 0 142582 800
rect 142894 0 142950 800
rect 143262 0 143318 800
rect 143630 0 143686 800
rect 143998 0 144054 800
rect 144366 0 144422 800
rect 144734 0 144790 800
rect 145102 0 145158 800
<< obsm2 >>
rect 1400 856 148560 150657
rect 1400 342 3734 856
rect 3902 342 4102 856
rect 4270 342 4470 856
rect 4638 342 4838 856
rect 5006 342 5206 856
rect 5374 342 5574 856
rect 5742 342 5942 856
rect 6110 342 6310 856
rect 6478 342 6678 856
rect 6846 342 7046 856
rect 7214 342 7414 856
rect 7582 342 7782 856
rect 7950 342 8150 856
rect 8318 342 8518 856
rect 8686 342 8886 856
rect 9054 342 9254 856
rect 9422 342 9622 856
rect 9790 342 9990 856
rect 10158 342 10358 856
rect 10526 342 10726 856
rect 10894 342 11094 856
rect 11262 342 11462 856
rect 11630 342 11830 856
rect 11998 342 12198 856
rect 12366 342 12566 856
rect 12734 342 12934 856
rect 13102 342 13302 856
rect 13470 342 13670 856
rect 13838 342 14038 856
rect 14206 342 14406 856
rect 14574 342 14774 856
rect 14942 342 15142 856
rect 15310 342 15510 856
rect 15678 342 15878 856
rect 16046 342 16246 856
rect 16414 342 16614 856
rect 16782 342 16982 856
rect 17150 342 17350 856
rect 17518 342 17718 856
rect 17886 342 18086 856
rect 18254 342 18454 856
rect 18622 342 18822 856
rect 18990 342 19190 856
rect 19358 342 19558 856
rect 19726 342 19926 856
rect 20094 342 20294 856
rect 20462 342 20662 856
rect 20830 342 21030 856
rect 21198 342 21398 856
rect 21566 342 21766 856
rect 21934 342 22134 856
rect 22302 342 22502 856
rect 22670 342 22870 856
rect 23038 342 23238 856
rect 23406 342 23606 856
rect 23774 342 23974 856
rect 24142 342 24342 856
rect 24510 342 24710 856
rect 24878 342 25078 856
rect 25246 342 25446 856
rect 25614 342 25814 856
rect 25982 342 26182 856
rect 26350 342 26550 856
rect 26718 342 26918 856
rect 27086 342 27286 856
rect 27454 342 27654 856
rect 27822 342 28022 856
rect 28190 342 28390 856
rect 28558 342 28758 856
rect 28926 342 29126 856
rect 29294 342 29494 856
rect 29662 342 29862 856
rect 30030 342 30230 856
rect 30398 342 30598 856
rect 30766 342 30966 856
rect 31134 342 31334 856
rect 31502 342 31702 856
rect 31870 342 32070 856
rect 32238 342 32438 856
rect 32606 342 32806 856
rect 32974 342 33174 856
rect 33342 342 33542 856
rect 33710 342 33910 856
rect 34078 342 34278 856
rect 34446 342 34646 856
rect 34814 342 35014 856
rect 35182 342 35382 856
rect 35550 342 35750 856
rect 35918 342 36118 856
rect 36286 342 36486 856
rect 36654 342 36854 856
rect 37022 342 37222 856
rect 37390 342 37590 856
rect 37758 342 37958 856
rect 38126 342 38326 856
rect 38494 342 38694 856
rect 38862 342 39062 856
rect 39230 342 39430 856
rect 39598 342 39798 856
rect 39966 342 40166 856
rect 40334 342 40534 856
rect 40702 342 40902 856
rect 41070 342 41270 856
rect 41438 342 41638 856
rect 41806 342 42006 856
rect 42174 342 42374 856
rect 42542 342 42742 856
rect 42910 342 43110 856
rect 43278 342 43478 856
rect 43646 342 43846 856
rect 44014 342 44214 856
rect 44382 342 44582 856
rect 44750 342 44950 856
rect 45118 342 45318 856
rect 45486 342 45686 856
rect 45854 342 46054 856
rect 46222 342 46422 856
rect 46590 342 46790 856
rect 46958 342 47158 856
rect 47326 342 47526 856
rect 47694 342 47894 856
rect 48062 342 48262 856
rect 48430 342 48630 856
rect 48798 342 48998 856
rect 49166 342 49366 856
rect 49534 342 49734 856
rect 49902 342 50102 856
rect 50270 342 50470 856
rect 50638 342 50838 856
rect 51006 342 51206 856
rect 51374 342 51574 856
rect 51742 342 51942 856
rect 52110 342 52310 856
rect 52478 342 52678 856
rect 52846 342 53046 856
rect 53214 342 53414 856
rect 53582 342 53782 856
rect 53950 342 54150 856
rect 54318 342 54518 856
rect 54686 342 54886 856
rect 55054 342 55254 856
rect 55422 342 55622 856
rect 55790 342 55990 856
rect 56158 342 56358 856
rect 56526 342 56726 856
rect 56894 342 57094 856
rect 57262 342 57462 856
rect 57630 342 57830 856
rect 57998 342 58198 856
rect 58366 342 58566 856
rect 58734 342 58934 856
rect 59102 342 59302 856
rect 59470 342 59670 856
rect 59838 342 60038 856
rect 60206 342 60406 856
rect 60574 342 60774 856
rect 60942 342 61142 856
rect 61310 342 61510 856
rect 61678 342 61878 856
rect 62046 342 62246 856
rect 62414 342 62614 856
rect 62782 342 62982 856
rect 63150 342 63350 856
rect 63518 342 63718 856
rect 63886 342 64086 856
rect 64254 342 64454 856
rect 64622 342 64822 856
rect 64990 342 65190 856
rect 65358 342 65558 856
rect 65726 342 65926 856
rect 66094 342 66294 856
rect 66462 342 66662 856
rect 66830 342 67030 856
rect 67198 342 67398 856
rect 67566 342 67766 856
rect 67934 342 68134 856
rect 68302 342 68502 856
rect 68670 342 68870 856
rect 69038 342 69238 856
rect 69406 342 69606 856
rect 69774 342 69974 856
rect 70142 342 70342 856
rect 70510 342 70710 856
rect 70878 342 71078 856
rect 71246 342 71446 856
rect 71614 342 71814 856
rect 71982 342 72182 856
rect 72350 342 72550 856
rect 72718 342 72918 856
rect 73086 342 73286 856
rect 73454 342 73654 856
rect 73822 342 74022 856
rect 74190 342 74390 856
rect 74558 342 74758 856
rect 74926 342 75126 856
rect 75294 342 75494 856
rect 75662 342 75862 856
rect 76030 342 76230 856
rect 76398 342 76598 856
rect 76766 342 76966 856
rect 77134 342 77334 856
rect 77502 342 77702 856
rect 77870 342 78070 856
rect 78238 342 78438 856
rect 78606 342 78806 856
rect 78974 342 79174 856
rect 79342 342 79542 856
rect 79710 342 79910 856
rect 80078 342 80278 856
rect 80446 342 80646 856
rect 80814 342 81014 856
rect 81182 342 81382 856
rect 81550 342 81750 856
rect 81918 342 82118 856
rect 82286 342 82486 856
rect 82654 342 82854 856
rect 83022 342 83222 856
rect 83390 342 83590 856
rect 83758 342 83958 856
rect 84126 342 84326 856
rect 84494 342 84694 856
rect 84862 342 85062 856
rect 85230 342 85430 856
rect 85598 342 85798 856
rect 85966 342 86166 856
rect 86334 342 86534 856
rect 86702 342 86902 856
rect 87070 342 87270 856
rect 87438 342 87638 856
rect 87806 342 88006 856
rect 88174 342 88374 856
rect 88542 342 88742 856
rect 88910 342 89110 856
rect 89278 342 89478 856
rect 89646 342 89846 856
rect 90014 342 90214 856
rect 90382 342 90582 856
rect 90750 342 90950 856
rect 91118 342 91318 856
rect 91486 342 91686 856
rect 91854 342 92054 856
rect 92222 342 92422 856
rect 92590 342 92790 856
rect 92958 342 93158 856
rect 93326 342 93526 856
rect 93694 342 93894 856
rect 94062 342 94262 856
rect 94430 342 94630 856
rect 94798 342 94998 856
rect 95166 342 95366 856
rect 95534 342 95734 856
rect 95902 342 96102 856
rect 96270 342 96470 856
rect 96638 342 96838 856
rect 97006 342 97206 856
rect 97374 342 97574 856
rect 97742 342 97942 856
rect 98110 342 98310 856
rect 98478 342 98678 856
rect 98846 342 99046 856
rect 99214 342 99414 856
rect 99582 342 99782 856
rect 99950 342 100150 856
rect 100318 342 100518 856
rect 100686 342 100886 856
rect 101054 342 101254 856
rect 101422 342 101622 856
rect 101790 342 101990 856
rect 102158 342 102358 856
rect 102526 342 102726 856
rect 102894 342 103094 856
rect 103262 342 103462 856
rect 103630 342 103830 856
rect 103998 342 104198 856
rect 104366 342 104566 856
rect 104734 342 104934 856
rect 105102 342 105302 856
rect 105470 342 105670 856
rect 105838 342 106038 856
rect 106206 342 106406 856
rect 106574 342 106774 856
rect 106942 342 107142 856
rect 107310 342 107510 856
rect 107678 342 107878 856
rect 108046 342 108246 856
rect 108414 342 108614 856
rect 108782 342 108982 856
rect 109150 342 109350 856
rect 109518 342 109718 856
rect 109886 342 110086 856
rect 110254 342 110454 856
rect 110622 342 110822 856
rect 110990 342 111190 856
rect 111358 342 111558 856
rect 111726 342 111926 856
rect 112094 342 112294 856
rect 112462 342 112662 856
rect 112830 342 113030 856
rect 113198 342 113398 856
rect 113566 342 113766 856
rect 113934 342 114134 856
rect 114302 342 114502 856
rect 114670 342 114870 856
rect 115038 342 115238 856
rect 115406 342 115606 856
rect 115774 342 115974 856
rect 116142 342 116342 856
rect 116510 342 116710 856
rect 116878 342 117078 856
rect 117246 342 117446 856
rect 117614 342 117814 856
rect 117982 342 118182 856
rect 118350 342 118550 856
rect 118718 342 118918 856
rect 119086 342 119286 856
rect 119454 342 119654 856
rect 119822 342 120022 856
rect 120190 342 120390 856
rect 120558 342 120758 856
rect 120926 342 121126 856
rect 121294 342 121494 856
rect 121662 342 121862 856
rect 122030 342 122230 856
rect 122398 342 122598 856
rect 122766 342 122966 856
rect 123134 342 123334 856
rect 123502 342 123702 856
rect 123870 342 124070 856
rect 124238 342 124438 856
rect 124606 342 124806 856
rect 124974 342 125174 856
rect 125342 342 125542 856
rect 125710 342 125910 856
rect 126078 342 126278 856
rect 126446 342 126646 856
rect 126814 342 127014 856
rect 127182 342 127382 856
rect 127550 342 127750 856
rect 127918 342 128118 856
rect 128286 342 128486 856
rect 128654 342 128854 856
rect 129022 342 129222 856
rect 129390 342 129590 856
rect 129758 342 129958 856
rect 130126 342 130326 856
rect 130494 342 130694 856
rect 130862 342 131062 856
rect 131230 342 131430 856
rect 131598 342 131798 856
rect 131966 342 132166 856
rect 132334 342 132534 856
rect 132702 342 132902 856
rect 133070 342 133270 856
rect 133438 342 133638 856
rect 133806 342 134006 856
rect 134174 342 134374 856
rect 134542 342 134742 856
rect 134910 342 135110 856
rect 135278 342 135478 856
rect 135646 342 135846 856
rect 136014 342 136214 856
rect 136382 342 136582 856
rect 136750 342 136950 856
rect 137118 342 137318 856
rect 137486 342 137686 856
rect 137854 342 138054 856
rect 138222 342 138422 856
rect 138590 342 138790 856
rect 138958 342 139158 856
rect 139326 342 139526 856
rect 139694 342 139894 856
rect 140062 342 140262 856
rect 140430 342 140630 856
rect 140798 342 140998 856
rect 141166 342 141366 856
rect 141534 342 141734 856
rect 141902 342 142102 856
rect 142270 342 142470 856
rect 142638 342 142838 856
rect 143006 342 143206 856
rect 143374 342 143574 856
rect 143742 342 143942 856
rect 144110 342 144310 856
rect 144478 342 144678 856
rect 144846 342 145046 856
rect 145214 342 148560 856
<< obsm3 >>
rect 1669 851 147831 150788
<< metal4 >>
rect 4208 2128 4528 148560
rect 19568 2128 19888 148560
rect 34928 2128 35248 148560
rect 50288 2128 50608 148560
rect 65648 2128 65968 148560
rect 81008 2128 81328 148560
rect 96368 2128 96688 148560
rect 111728 2128 112048 148560
rect 127088 2128 127408 148560
rect 142448 2128 142768 148560
<< obsm4 >>
rect 2451 148640 146221 150789
rect 2451 2048 4128 148640
rect 4608 2048 19488 148640
rect 19968 2048 34848 148640
rect 35328 2048 50208 148640
rect 50688 2048 65568 148640
rect 66048 2048 80928 148640
rect 81408 2048 96288 148640
rect 96768 2048 111648 148640
rect 112128 2048 127008 148640
rect 127488 2048 142368 148640
rect 142848 2048 146221 148640
rect 2451 1531 146221 2048
<< labels >>
rlabel metal2 s 145102 0 145158 800 6 clk
port 1 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 la_data_in[0]
port 2 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 la_data_in[100]
port 3 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 la_data_in[101]
port 4 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_data_in[102]
port 5 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 la_data_in[103]
port 6 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 la_data_in[104]
port 7 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 la_data_in[105]
port 8 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 la_data_in[106]
port 9 nsew signal input
rlabel metal2 s 121918 0 121974 800 6 la_data_in[107]
port 10 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_data_in[108]
port 11 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 la_data_in[109]
port 12 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 la_data_in[10]
port 13 nsew signal input
rlabel metal2 s 125230 0 125286 800 6 la_data_in[110]
port 14 nsew signal input
rlabel metal2 s 126334 0 126390 800 6 la_data_in[111]
port 15 nsew signal input
rlabel metal2 s 127438 0 127494 800 6 la_data_in[112]
port 16 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 la_data_in[113]
port 17 nsew signal input
rlabel metal2 s 129646 0 129702 800 6 la_data_in[114]
port 18 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 la_data_in[115]
port 19 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 la_data_in[116]
port 20 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 la_data_in[117]
port 21 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 la_data_in[118]
port 22 nsew signal input
rlabel metal2 s 135166 0 135222 800 6 la_data_in[119]
port 23 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 la_data_in[11]
port 24 nsew signal input
rlabel metal2 s 136270 0 136326 800 6 la_data_in[120]
port 25 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 la_data_in[121]
port 26 nsew signal input
rlabel metal2 s 138478 0 138534 800 6 la_data_in[122]
port 27 nsew signal input
rlabel metal2 s 139582 0 139638 800 6 la_data_in[123]
port 28 nsew signal input
rlabel metal2 s 140686 0 140742 800 6 la_data_in[124]
port 29 nsew signal input
rlabel metal2 s 141790 0 141846 800 6 la_data_in[125]
port 30 nsew signal input
rlabel metal2 s 142894 0 142950 800 6 la_data_in[126]
port 31 nsew signal input
rlabel metal2 s 143998 0 144054 800 6 la_data_in[127]
port 32 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 la_data_in[12]
port 33 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 la_data_in[13]
port 34 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 la_data_in[14]
port 35 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 la_data_in[15]
port 36 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 la_data_in[16]
port 37 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 la_data_in[17]
port 38 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 la_data_in[18]
port 39 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 la_data_in[19]
port 40 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 la_data_in[1]
port 41 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 la_data_in[20]
port 42 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 la_data_in[21]
port 43 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 la_data_in[22]
port 44 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 la_data_in[23]
port 45 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 la_data_in[24]
port 46 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 la_data_in[25]
port 47 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 la_data_in[26]
port 48 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_data_in[27]
port 49 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 la_data_in[28]
port 50 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 la_data_in[29]
port 51 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 la_data_in[2]
port 52 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 la_data_in[30]
port 53 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 la_data_in[31]
port 54 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_data_in[32]
port 55 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_data_in[33]
port 56 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 la_data_in[34]
port 57 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 la_data_in[35]
port 58 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_data_in[36]
port 59 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 la_data_in[37]
port 60 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la_data_in[38]
port 61 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_data_in[39]
port 62 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 la_data_in[3]
port 63 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 la_data_in[40]
port 64 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_data_in[41]
port 65 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 la_data_in[42]
port 66 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 la_data_in[43]
port 67 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 la_data_in[44]
port 68 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 la_data_in[45]
port 69 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 la_data_in[46]
port 70 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_data_in[47]
port 71 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_data_in[48]
port 72 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 la_data_in[49]
port 73 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 la_data_in[4]
port 74 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 la_data_in[50]
port 75 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 la_data_in[51]
port 76 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_data_in[52]
port 77 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_data_in[53]
port 78 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_data_in[54]
port 79 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 la_data_in[55]
port 80 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 la_data_in[56]
port 81 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_data_in[57]
port 82 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_data_in[58]
port 83 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 la_data_in[59]
port 84 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 la_data_in[5]
port 85 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 la_data_in[60]
port 86 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_data_in[61]
port 87 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 la_data_in[62]
port 88 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 la_data_in[63]
port 89 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 la_data_in[64]
port 90 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 la_data_in[65]
port 91 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 la_data_in[66]
port 92 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 la_data_in[67]
port 93 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_data_in[68]
port 94 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_data_in[69]
port 95 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 la_data_in[6]
port 96 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 la_data_in[70]
port 97 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_data_in[71]
port 98 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_data_in[72]
port 99 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_data_in[73]
port 100 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 la_data_in[74]
port 101 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 la_data_in[75]
port 102 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_data_in[76]
port 103 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_data_in[77]
port 104 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_data_in[78]
port 105 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 la_data_in[79]
port 106 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 la_data_in[7]
port 107 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_data_in[80]
port 108 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_data_in[81]
port 109 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 la_data_in[82]
port 110 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_data_in[83]
port 111 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_data_in[84]
port 112 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_data_in[85]
port 113 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 la_data_in[86]
port 114 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_data_in[87]
port 115 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 la_data_in[88]
port 116 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 la_data_in[89]
port 117 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 la_data_in[8]
port 118 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 la_data_in[90]
port 119 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 la_data_in[91]
port 120 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 la_data_in[92]
port 121 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_data_in[93]
port 122 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_data_in[94]
port 123 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 la_data_in[95]
port 124 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 la_data_in[96]
port 125 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 la_data_in[97]
port 126 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 la_data_in[98]
port 127 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 la_data_in[99]
port 128 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 la_data_in[9]
port 129 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 la_data_out[0]
port 130 nsew signal output
rlabel metal2 s 114558 0 114614 800 6 la_data_out[100]
port 131 nsew signal output
rlabel metal2 s 115662 0 115718 800 6 la_data_out[101]
port 132 nsew signal output
rlabel metal2 s 116766 0 116822 800 6 la_data_out[102]
port 133 nsew signal output
rlabel metal2 s 117870 0 117926 800 6 la_data_out[103]
port 134 nsew signal output
rlabel metal2 s 118974 0 119030 800 6 la_data_out[104]
port 135 nsew signal output
rlabel metal2 s 120078 0 120134 800 6 la_data_out[105]
port 136 nsew signal output
rlabel metal2 s 121182 0 121238 800 6 la_data_out[106]
port 137 nsew signal output
rlabel metal2 s 122286 0 122342 800 6 la_data_out[107]
port 138 nsew signal output
rlabel metal2 s 123390 0 123446 800 6 la_data_out[108]
port 139 nsew signal output
rlabel metal2 s 124494 0 124550 800 6 la_data_out[109]
port 140 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 la_data_out[10]
port 141 nsew signal output
rlabel metal2 s 125598 0 125654 800 6 la_data_out[110]
port 142 nsew signal output
rlabel metal2 s 126702 0 126758 800 6 la_data_out[111]
port 143 nsew signal output
rlabel metal2 s 127806 0 127862 800 6 la_data_out[112]
port 144 nsew signal output
rlabel metal2 s 128910 0 128966 800 6 la_data_out[113]
port 145 nsew signal output
rlabel metal2 s 130014 0 130070 800 6 la_data_out[114]
port 146 nsew signal output
rlabel metal2 s 131118 0 131174 800 6 la_data_out[115]
port 147 nsew signal output
rlabel metal2 s 132222 0 132278 800 6 la_data_out[116]
port 148 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 la_data_out[117]
port 149 nsew signal output
rlabel metal2 s 134430 0 134486 800 6 la_data_out[118]
port 150 nsew signal output
rlabel metal2 s 135534 0 135590 800 6 la_data_out[119]
port 151 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 la_data_out[11]
port 152 nsew signal output
rlabel metal2 s 136638 0 136694 800 6 la_data_out[120]
port 153 nsew signal output
rlabel metal2 s 137742 0 137798 800 6 la_data_out[121]
port 154 nsew signal output
rlabel metal2 s 138846 0 138902 800 6 la_data_out[122]
port 155 nsew signal output
rlabel metal2 s 139950 0 140006 800 6 la_data_out[123]
port 156 nsew signal output
rlabel metal2 s 141054 0 141110 800 6 la_data_out[124]
port 157 nsew signal output
rlabel metal2 s 142158 0 142214 800 6 la_data_out[125]
port 158 nsew signal output
rlabel metal2 s 143262 0 143318 800 6 la_data_out[126]
port 159 nsew signal output
rlabel metal2 s 144366 0 144422 800 6 la_data_out[127]
port 160 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 la_data_out[12]
port 161 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 la_data_out[13]
port 162 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 la_data_out[14]
port 163 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 la_data_out[15]
port 164 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 la_data_out[16]
port 165 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 la_data_out[17]
port 166 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 la_data_out[18]
port 167 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 la_data_out[19]
port 168 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 la_data_out[1]
port 169 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 la_data_out[20]
port 170 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 la_data_out[21]
port 171 nsew signal output
rlabel metal2 s 28446 0 28502 800 6 la_data_out[22]
port 172 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 la_data_out[23]
port 173 nsew signal output
rlabel metal2 s 30654 0 30710 800 6 la_data_out[24]
port 174 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 la_data_out[25]
port 175 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 la_data_out[26]
port 176 nsew signal output
rlabel metal2 s 33966 0 34022 800 6 la_data_out[27]
port 177 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 la_data_out[28]
port 178 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 la_data_out[29]
port 179 nsew signal output
rlabel metal2 s 6366 0 6422 800 6 la_data_out[2]
port 180 nsew signal output
rlabel metal2 s 37278 0 37334 800 6 la_data_out[30]
port 181 nsew signal output
rlabel metal2 s 38382 0 38438 800 6 la_data_out[31]
port 182 nsew signal output
rlabel metal2 s 39486 0 39542 800 6 la_data_out[32]
port 183 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 la_data_out[33]
port 184 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 la_data_out[34]
port 185 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 la_data_out[35]
port 186 nsew signal output
rlabel metal2 s 43902 0 43958 800 6 la_data_out[36]
port 187 nsew signal output
rlabel metal2 s 45006 0 45062 800 6 la_data_out[37]
port 188 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 la_data_out[38]
port 189 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 la_data_out[39]
port 190 nsew signal output
rlabel metal2 s 7470 0 7526 800 6 la_data_out[3]
port 191 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 la_data_out[40]
port 192 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 la_data_out[41]
port 193 nsew signal output
rlabel metal2 s 50526 0 50582 800 6 la_data_out[42]
port 194 nsew signal output
rlabel metal2 s 51630 0 51686 800 6 la_data_out[43]
port 195 nsew signal output
rlabel metal2 s 52734 0 52790 800 6 la_data_out[44]
port 196 nsew signal output
rlabel metal2 s 53838 0 53894 800 6 la_data_out[45]
port 197 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 la_data_out[46]
port 198 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 la_data_out[47]
port 199 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 la_data_out[48]
port 200 nsew signal output
rlabel metal2 s 58254 0 58310 800 6 la_data_out[49]
port 201 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 la_data_out[4]
port 202 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 la_data_out[50]
port 203 nsew signal output
rlabel metal2 s 60462 0 60518 800 6 la_data_out[51]
port 204 nsew signal output
rlabel metal2 s 61566 0 61622 800 6 la_data_out[52]
port 205 nsew signal output
rlabel metal2 s 62670 0 62726 800 6 la_data_out[53]
port 206 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 la_data_out[54]
port 207 nsew signal output
rlabel metal2 s 64878 0 64934 800 6 la_data_out[55]
port 208 nsew signal output
rlabel metal2 s 65982 0 66038 800 6 la_data_out[56]
port 209 nsew signal output
rlabel metal2 s 67086 0 67142 800 6 la_data_out[57]
port 210 nsew signal output
rlabel metal2 s 68190 0 68246 800 6 la_data_out[58]
port 211 nsew signal output
rlabel metal2 s 69294 0 69350 800 6 la_data_out[59]
port 212 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 la_data_out[5]
port 213 nsew signal output
rlabel metal2 s 70398 0 70454 800 6 la_data_out[60]
port 214 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 la_data_out[61]
port 215 nsew signal output
rlabel metal2 s 72606 0 72662 800 6 la_data_out[62]
port 216 nsew signal output
rlabel metal2 s 73710 0 73766 800 6 la_data_out[63]
port 217 nsew signal output
rlabel metal2 s 74814 0 74870 800 6 la_data_out[64]
port 218 nsew signal output
rlabel metal2 s 75918 0 75974 800 6 la_data_out[65]
port 219 nsew signal output
rlabel metal2 s 77022 0 77078 800 6 la_data_out[66]
port 220 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 la_data_out[67]
port 221 nsew signal output
rlabel metal2 s 79230 0 79286 800 6 la_data_out[68]
port 222 nsew signal output
rlabel metal2 s 80334 0 80390 800 6 la_data_out[69]
port 223 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 la_data_out[6]
port 224 nsew signal output
rlabel metal2 s 81438 0 81494 800 6 la_data_out[70]
port 225 nsew signal output
rlabel metal2 s 82542 0 82598 800 6 la_data_out[71]
port 226 nsew signal output
rlabel metal2 s 83646 0 83702 800 6 la_data_out[72]
port 227 nsew signal output
rlabel metal2 s 84750 0 84806 800 6 la_data_out[73]
port 228 nsew signal output
rlabel metal2 s 85854 0 85910 800 6 la_data_out[74]
port 229 nsew signal output
rlabel metal2 s 86958 0 87014 800 6 la_data_out[75]
port 230 nsew signal output
rlabel metal2 s 88062 0 88118 800 6 la_data_out[76]
port 231 nsew signal output
rlabel metal2 s 89166 0 89222 800 6 la_data_out[77]
port 232 nsew signal output
rlabel metal2 s 90270 0 90326 800 6 la_data_out[78]
port 233 nsew signal output
rlabel metal2 s 91374 0 91430 800 6 la_data_out[79]
port 234 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 la_data_out[7]
port 235 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 la_data_out[80]
port 236 nsew signal output
rlabel metal2 s 93582 0 93638 800 6 la_data_out[81]
port 237 nsew signal output
rlabel metal2 s 94686 0 94742 800 6 la_data_out[82]
port 238 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 la_data_out[83]
port 239 nsew signal output
rlabel metal2 s 96894 0 96950 800 6 la_data_out[84]
port 240 nsew signal output
rlabel metal2 s 97998 0 98054 800 6 la_data_out[85]
port 241 nsew signal output
rlabel metal2 s 99102 0 99158 800 6 la_data_out[86]
port 242 nsew signal output
rlabel metal2 s 100206 0 100262 800 6 la_data_out[87]
port 243 nsew signal output
rlabel metal2 s 101310 0 101366 800 6 la_data_out[88]
port 244 nsew signal output
rlabel metal2 s 102414 0 102470 800 6 la_data_out[89]
port 245 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 la_data_out[8]
port 246 nsew signal output
rlabel metal2 s 103518 0 103574 800 6 la_data_out[90]
port 247 nsew signal output
rlabel metal2 s 104622 0 104678 800 6 la_data_out[91]
port 248 nsew signal output
rlabel metal2 s 105726 0 105782 800 6 la_data_out[92]
port 249 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 la_data_out[93]
port 250 nsew signal output
rlabel metal2 s 107934 0 107990 800 6 la_data_out[94]
port 251 nsew signal output
rlabel metal2 s 109038 0 109094 800 6 la_data_out[95]
port 252 nsew signal output
rlabel metal2 s 110142 0 110198 800 6 la_data_out[96]
port 253 nsew signal output
rlabel metal2 s 111246 0 111302 800 6 la_data_out[97]
port 254 nsew signal output
rlabel metal2 s 112350 0 112406 800 6 la_data_out[98]
port 255 nsew signal output
rlabel metal2 s 113454 0 113510 800 6 la_data_out[99]
port 256 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 la_data_out[9]
port 257 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 la_oenb[0]
port 258 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 la_oenb[100]
port 259 nsew signal input
rlabel metal2 s 116030 0 116086 800 6 la_oenb[101]
port 260 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 la_oenb[102]
port 261 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 la_oenb[103]
port 262 nsew signal input
rlabel metal2 s 119342 0 119398 800 6 la_oenb[104]
port 263 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 la_oenb[105]
port 264 nsew signal input
rlabel metal2 s 121550 0 121606 800 6 la_oenb[106]
port 265 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 la_oenb[107]
port 266 nsew signal input
rlabel metal2 s 123758 0 123814 800 6 la_oenb[108]
port 267 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 la_oenb[109]
port 268 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 la_oenb[10]
port 269 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 la_oenb[110]
port 270 nsew signal input
rlabel metal2 s 127070 0 127126 800 6 la_oenb[111]
port 271 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 la_oenb[112]
port 272 nsew signal input
rlabel metal2 s 129278 0 129334 800 6 la_oenb[113]
port 273 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 la_oenb[114]
port 274 nsew signal input
rlabel metal2 s 131486 0 131542 800 6 la_oenb[115]
port 275 nsew signal input
rlabel metal2 s 132590 0 132646 800 6 la_oenb[116]
port 276 nsew signal input
rlabel metal2 s 133694 0 133750 800 6 la_oenb[117]
port 277 nsew signal input
rlabel metal2 s 134798 0 134854 800 6 la_oenb[118]
port 278 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 la_oenb[119]
port 279 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 la_oenb[11]
port 280 nsew signal input
rlabel metal2 s 137006 0 137062 800 6 la_oenb[120]
port 281 nsew signal input
rlabel metal2 s 138110 0 138166 800 6 la_oenb[121]
port 282 nsew signal input
rlabel metal2 s 139214 0 139270 800 6 la_oenb[122]
port 283 nsew signal input
rlabel metal2 s 140318 0 140374 800 6 la_oenb[123]
port 284 nsew signal input
rlabel metal2 s 141422 0 141478 800 6 la_oenb[124]
port 285 nsew signal input
rlabel metal2 s 142526 0 142582 800 6 la_oenb[125]
port 286 nsew signal input
rlabel metal2 s 143630 0 143686 800 6 la_oenb[126]
port 287 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 la_oenb[127]
port 288 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 la_oenb[12]
port 289 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 la_oenb[13]
port 290 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 la_oenb[14]
port 291 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 la_oenb[15]
port 292 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 la_oenb[16]
port 293 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 la_oenb[17]
port 294 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 la_oenb[18]
port 295 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 la_oenb[19]
port 296 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 la_oenb[1]
port 297 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 la_oenb[20]
port 298 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_oenb[21]
port 299 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 la_oenb[22]
port 300 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_oenb[23]
port 301 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 la_oenb[24]
port 302 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 la_oenb[25]
port 303 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 la_oenb[26]
port 304 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 la_oenb[27]
port 305 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_oenb[28]
port 306 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_oenb[29]
port 307 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 la_oenb[2]
port 308 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 la_oenb[30]
port 309 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 la_oenb[31]
port 310 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 la_oenb[32]
port 311 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 la_oenb[33]
port 312 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 la_oenb[34]
port 313 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_oenb[35]
port 314 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 la_oenb[36]
port 315 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 la_oenb[37]
port 316 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_oenb[38]
port 317 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_oenb[39]
port 318 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 la_oenb[3]
port 319 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 la_oenb[40]
port 320 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 la_oenb[41]
port 321 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 la_oenb[42]
port 322 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 la_oenb[43]
port 323 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 la_oenb[44]
port 324 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 la_oenb[45]
port 325 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 la_oenb[46]
port 326 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 la_oenb[47]
port 327 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 la_oenb[48]
port 328 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_oenb[49]
port 329 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 la_oenb[4]
port 330 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 la_oenb[50]
port 331 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 la_oenb[51]
port 332 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 la_oenb[52]
port 333 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_oenb[53]
port 334 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 la_oenb[54]
port 335 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 la_oenb[55]
port 336 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 la_oenb[56]
port 337 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 la_oenb[57]
port 338 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_oenb[58]
port 339 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_oenb[59]
port 340 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 la_oenb[5]
port 341 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 la_oenb[60]
port 342 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 la_oenb[61]
port 343 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_oenb[62]
port 344 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_oenb[63]
port 345 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 la_oenb[64]
port 346 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 la_oenb[65]
port 347 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 la_oenb[66]
port 348 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_oenb[67]
port 349 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_oenb[68]
port 350 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 la_oenb[69]
port 351 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 la_oenb[6]
port 352 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_oenb[70]
port 353 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 la_oenb[71]
port 354 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_oenb[72]
port 355 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_oenb[73]
port 356 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_oenb[74]
port 357 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 la_oenb[75]
port 358 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_oenb[76]
port 359 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_oenb[77]
port 360 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_oenb[78]
port 361 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_oenb[79]
port 362 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 la_oenb[7]
port 363 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_oenb[80]
port 364 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 la_oenb[81]
port 365 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 la_oenb[82]
port 366 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 la_oenb[83]
port 367 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_oenb[84]
port 368 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_oenb[85]
port 369 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_oenb[86]
port 370 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 la_oenb[87]
port 371 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_oenb[88]
port 372 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 la_oenb[89]
port 373 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 la_oenb[8]
port 374 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 la_oenb[90]
port 375 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 la_oenb[91]
port 376 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 la_oenb[92]
port 377 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 la_oenb[93]
port 378 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 la_oenb[94]
port 379 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 la_oenb[95]
port 380 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 la_oenb[96]
port 381 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 la_oenb[97]
port 382 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 la_oenb[98]
port 383 nsew signal input
rlabel metal2 s 113822 0 113878 800 6 la_oenb[99]
port 384 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 la_oenb[9]
port 385 nsew signal input
rlabel metal4 s 4208 2128 4528 148560 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 148560 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 148560 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 148560 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 148560 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 148560 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 148560 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 148560 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 148560 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 148560 6 vssd1
port 387 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 148918 151062
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 62159182
string GDS_FILE /home/drewarosa/RISC-V-Single-Cycle-CPU-Core/openlane/RISC_V/runs/22_09_22_09_03/results/signoff/RISC_V.magic.gds
string GDS_START 1104428
<< end >>

