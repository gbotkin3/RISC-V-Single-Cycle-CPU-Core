VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pc
  CLASS BLOCK ;
  FOREIGN pc ;
  ORIGIN 0.000 0.000 ;
  SIZE 277.485 BY 288.205 ;
  PIN alu_branch
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 47.640 277.485 48.240 ;
    END
  END alu_branch
  PIN branch
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 241.440 277.485 242.040 ;
    END
  END branch
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 284.205 158.150 288.205 ;
    END
  END clk
  PIN immediate[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 275.440 277.485 276.040 ;
    END
  END immediate[0]
  PIN immediate[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END immediate[10]
  PIN immediate[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END immediate[11]
  PIN immediate[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END immediate[12]
  PIN immediate[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 284.205 267.630 288.205 ;
    END
  END immediate[13]
  PIN immediate[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END immediate[14]
  PIN immediate[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END immediate[15]
  PIN immediate[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END immediate[16]
  PIN immediate[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END immediate[17]
  PIN immediate[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END immediate[18]
  PIN immediate[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END immediate[19]
  PIN immediate[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END immediate[1]
  PIN immediate[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END immediate[20]
  PIN immediate[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 207.440 277.485 208.040 ;
    END
  END immediate[21]
  PIN immediate[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 284.205 125.950 288.205 ;
    END
  END immediate[22]
  PIN immediate[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END immediate[23]
  PIN immediate[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END immediate[24]
  PIN immediate[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END immediate[25]
  PIN immediate[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END immediate[26]
  PIN immediate[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END immediate[27]
  PIN immediate[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END immediate[28]
  PIN immediate[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 0.040 277.485 0.640 ;
    END
  END immediate[29]
  PIN immediate[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END immediate[2]
  PIN immediate[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 149.640 277.485 150.240 ;
    END
  END immediate[30]
  PIN immediate[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 284.205 171.030 288.205 ;
    END
  END immediate[31]
  PIN immediate[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 284.205 93.750 288.205 ;
    END
  END immediate[3]
  PIN immediate[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 265.240 277.485 265.840 ;
    END
  END immediate[4]
  PIN immediate[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END immediate[5]
  PIN immediate[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END immediate[6]
  PIN immediate[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 251.640 277.485 252.240 ;
    END
  END immediate[7]
  PIN immediate[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 284.205 106.630 288.205 ;
    END
  END immediate[8]
  PIN immediate[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 68.040 277.485 68.640 ;
    END
  END immediate[9]
  PIN jump_jal
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 91.840 277.485 92.440 ;
    END
  END jump_jal
  PIN jump_jalr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 284.205 116.290 288.205 ;
    END
  END jump_jalr
  PIN pc_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 284.205 71.210 288.205 ;
    END
  END pc_out[0]
  PIN pc_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END pc_out[10]
  PIN pc_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END pc_out[11]
  PIN pc_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 217.640 277.485 218.240 ;
    END
  END pc_out[12]
  PIN pc_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END pc_out[13]
  PIN pc_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 115.640 277.485 116.240 ;
    END
  END pc_out[14]
  PIN pc_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 284.205 203.230 288.205 ;
    END
  END pc_out[15]
  PIN pc_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 284.205 84.090 288.205 ;
    END
  END pc_out[16]
  PIN pc_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 13.640 277.485 14.240 ;
    END
  END pc_out[17]
  PIN pc_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 231.240 277.485 231.840 ;
    END
  END pc_out[18]
  PIN pc_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 284.205 257.970 288.205 ;
    END
  END pc_out[19]
  PIN pc_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 284.205 148.490 288.205 ;
    END
  END pc_out[1]
  PIN pc_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END pc_out[20]
  PIN pc_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 57.840 277.485 58.440 ;
    END
  END pc_out[21]
  PIN pc_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END pc_out[22]
  PIN pc_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END pc_out[23]
  PIN pc_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 284.205 180.690 288.205 ;
    END
  END pc_out[24]
  PIN pc_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END pc_out[25]
  PIN pc_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END pc_out[26]
  PIN pc_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 284.205 235.430 288.205 ;
    END
  END pc_out[27]
  PIN pc_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END pc_out[28]
  PIN pc_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END pc_out[29]
  PIN pc_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END pc_out[2]
  PIN pc_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END pc_out[30]
  PIN pc_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 125.840 277.485 126.440 ;
    END
  END pc_out[31]
  PIN pc_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 81.640 277.485 82.240 ;
    END
  END pc_out[3]
  PIN pc_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END pc_out[4]
  PIN pc_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END pc_out[5]
  PIN pc_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 23.840 277.485 24.440 ;
    END
  END pc_out[6]
  PIN pc_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 284.205 29.350 288.205 ;
    END
  END pc_out[7]
  PIN pc_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 105.440 277.485 106.040 ;
    END
  END pc_out[8]
  PIN pc_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 183.640 277.485 184.240 ;
    END
  END pc_out[9]
  PIN rs1_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END rs1_data[0]
  PIN rs1_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 197.240 277.485 197.840 ;
    END
  END rs1_data[10]
  PIN rs1_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 284.205 39.010 288.205 ;
    END
  END rs1_data[11]
  PIN rs1_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END rs1_data[12]
  PIN rs1_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END rs1_data[13]
  PIN rs1_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END rs1_data[14]
  PIN rs1_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END rs1_data[15]
  PIN rs1_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 284.205 51.890 288.205 ;
    END
  END rs1_data[16]
  PIN rs1_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 284.205 138.830 288.205 ;
    END
  END rs1_data[17]
  PIN rs1_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END rs1_data[18]
  PIN rs1_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END rs1_data[19]
  PIN rs1_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END rs1_data[1]
  PIN rs1_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END rs1_data[20]
  PIN rs1_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 284.205 245.090 288.205 ;
    END
  END rs1_data[21]
  PIN rs1_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 284.205 193.570 288.205 ;
    END
  END rs1_data[22]
  PIN rs1_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END rs1_data[23]
  PIN rs1_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 284.205 277.290 288.205 ;
    END
  END rs1_data[24]
  PIN rs1_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 34.040 277.485 34.640 ;
    END
  END rs1_data[25]
  PIN rs1_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 284.205 6.810 288.205 ;
    END
  END rs1_data[26]
  PIN rs1_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 159.840 277.485 160.440 ;
    END
  END rs1_data[27]
  PIN rs1_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END rs1_data[28]
  PIN rs1_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END rs1_data[29]
  PIN rs1_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END rs1_data[2]
  PIN rs1_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 173.440 277.485 174.040 ;
    END
  END rs1_data[30]
  PIN rs1_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END rs1_data[31]
  PIN rs1_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 284.205 225.770 288.205 ;
    END
  END rs1_data[3]
  PIN rs1_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 284.205 212.890 288.205 ;
    END
  END rs1_data[4]
  PIN rs1_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 284.205 19.690 288.205 ;
    END
  END rs1_data[5]
  PIN rs1_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 284.205 61.550 288.205 ;
    END
  END rs1_data[6]
  PIN rs1_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END rs1_data[7]
  PIN rs1_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END rs1_data[8]
  PIN rs1_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END rs1_data[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.485 139.440 277.485 140.040 ;
    END
  END rst_n
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 274.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 274.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 274.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 274.960 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 271.860 274.805 ;
      LAYER met1 ;
        RECT 0.070 9.220 277.310 274.960 ;
      LAYER met2 ;
        RECT 0.100 283.925 6.250 286.125 ;
        RECT 7.090 283.925 19.130 286.125 ;
        RECT 19.970 283.925 28.790 286.125 ;
        RECT 29.630 283.925 38.450 286.125 ;
        RECT 39.290 283.925 51.330 286.125 ;
        RECT 52.170 283.925 60.990 286.125 ;
        RECT 61.830 283.925 70.650 286.125 ;
        RECT 71.490 283.925 83.530 286.125 ;
        RECT 84.370 283.925 93.190 286.125 ;
        RECT 94.030 283.925 106.070 286.125 ;
        RECT 106.910 283.925 115.730 286.125 ;
        RECT 116.570 283.925 125.390 286.125 ;
        RECT 126.230 283.925 138.270 286.125 ;
        RECT 139.110 283.925 147.930 286.125 ;
        RECT 148.770 283.925 157.590 286.125 ;
        RECT 158.430 283.925 170.470 286.125 ;
        RECT 171.310 283.925 180.130 286.125 ;
        RECT 180.970 283.925 193.010 286.125 ;
        RECT 193.850 283.925 202.670 286.125 ;
        RECT 203.510 283.925 212.330 286.125 ;
        RECT 213.170 283.925 225.210 286.125 ;
        RECT 226.050 283.925 234.870 286.125 ;
        RECT 235.710 283.925 244.530 286.125 ;
        RECT 245.370 283.925 257.410 286.125 ;
        RECT 258.250 283.925 267.070 286.125 ;
        RECT 267.910 283.925 276.730 286.125 ;
        RECT 0.100 4.280 277.280 283.925 ;
        RECT 0.650 0.155 9.470 4.280 ;
        RECT 10.310 0.155 19.130 4.280 ;
        RECT 19.970 0.155 32.010 4.280 ;
        RECT 32.850 0.155 41.670 4.280 ;
        RECT 42.510 0.155 51.330 4.280 ;
        RECT 52.170 0.155 64.210 4.280 ;
        RECT 65.050 0.155 73.870 4.280 ;
        RECT 74.710 0.155 83.530 4.280 ;
        RECT 84.370 0.155 96.410 4.280 ;
        RECT 97.250 0.155 106.070 4.280 ;
        RECT 106.910 0.155 118.950 4.280 ;
        RECT 119.790 0.155 128.610 4.280 ;
        RECT 129.450 0.155 138.270 4.280 ;
        RECT 139.110 0.155 151.150 4.280 ;
        RECT 151.990 0.155 160.810 4.280 ;
        RECT 161.650 0.155 170.470 4.280 ;
        RECT 171.310 0.155 183.350 4.280 ;
        RECT 184.190 0.155 193.010 4.280 ;
        RECT 193.850 0.155 205.890 4.280 ;
        RECT 206.730 0.155 215.550 4.280 ;
        RECT 216.390 0.155 225.210 4.280 ;
        RECT 226.050 0.155 238.090 4.280 ;
        RECT 238.930 0.155 247.750 4.280 ;
        RECT 248.590 0.155 257.410 4.280 ;
        RECT 258.250 0.155 270.290 4.280 ;
        RECT 271.130 0.155 277.280 4.280 ;
      LAYER met3 ;
        RECT 4.400 285.240 273.485 286.105 ;
        RECT 4.000 276.440 273.485 285.240 ;
        RECT 4.000 275.040 273.085 276.440 ;
        RECT 4.000 273.040 273.485 275.040 ;
        RECT 4.400 271.640 273.485 273.040 ;
        RECT 4.000 266.240 273.485 271.640 ;
        RECT 4.000 264.840 273.085 266.240 ;
        RECT 4.000 262.840 273.485 264.840 ;
        RECT 4.400 261.440 273.485 262.840 ;
        RECT 4.000 252.640 273.485 261.440 ;
        RECT 4.400 251.240 273.085 252.640 ;
        RECT 4.000 242.440 273.485 251.240 ;
        RECT 4.000 241.040 273.085 242.440 ;
        RECT 4.000 239.040 273.485 241.040 ;
        RECT 4.400 237.640 273.485 239.040 ;
        RECT 4.000 232.240 273.485 237.640 ;
        RECT 4.000 230.840 273.085 232.240 ;
        RECT 4.000 228.840 273.485 230.840 ;
        RECT 4.400 227.440 273.485 228.840 ;
        RECT 4.000 218.640 273.485 227.440 ;
        RECT 4.400 217.240 273.085 218.640 ;
        RECT 4.000 208.440 273.485 217.240 ;
        RECT 4.000 207.040 273.085 208.440 ;
        RECT 4.000 205.040 273.485 207.040 ;
        RECT 4.400 203.640 273.485 205.040 ;
        RECT 4.000 198.240 273.485 203.640 ;
        RECT 4.000 196.840 273.085 198.240 ;
        RECT 4.000 194.840 273.485 196.840 ;
        RECT 4.400 193.440 273.485 194.840 ;
        RECT 4.000 184.640 273.485 193.440 ;
        RECT 4.000 183.240 273.085 184.640 ;
        RECT 4.000 181.240 273.485 183.240 ;
        RECT 4.400 179.840 273.485 181.240 ;
        RECT 4.000 174.440 273.485 179.840 ;
        RECT 4.000 173.040 273.085 174.440 ;
        RECT 4.000 171.040 273.485 173.040 ;
        RECT 4.400 169.640 273.485 171.040 ;
        RECT 4.000 160.840 273.485 169.640 ;
        RECT 4.400 159.440 273.085 160.840 ;
        RECT 4.000 150.640 273.485 159.440 ;
        RECT 4.000 149.240 273.085 150.640 ;
        RECT 4.000 147.240 273.485 149.240 ;
        RECT 4.400 145.840 273.485 147.240 ;
        RECT 4.000 140.440 273.485 145.840 ;
        RECT 4.000 139.040 273.085 140.440 ;
        RECT 4.000 137.040 273.485 139.040 ;
        RECT 4.400 135.640 273.485 137.040 ;
        RECT 4.000 126.840 273.485 135.640 ;
        RECT 4.400 125.440 273.085 126.840 ;
        RECT 4.000 116.640 273.485 125.440 ;
        RECT 4.000 115.240 273.085 116.640 ;
        RECT 4.000 113.240 273.485 115.240 ;
        RECT 4.400 111.840 273.485 113.240 ;
        RECT 4.000 106.440 273.485 111.840 ;
        RECT 4.000 105.040 273.085 106.440 ;
        RECT 4.000 103.040 273.485 105.040 ;
        RECT 4.400 101.640 273.485 103.040 ;
        RECT 4.000 92.840 273.485 101.640 ;
        RECT 4.000 91.440 273.085 92.840 ;
        RECT 4.000 89.440 273.485 91.440 ;
        RECT 4.400 88.040 273.485 89.440 ;
        RECT 4.000 82.640 273.485 88.040 ;
        RECT 4.000 81.240 273.085 82.640 ;
        RECT 4.000 79.240 273.485 81.240 ;
        RECT 4.400 77.840 273.485 79.240 ;
        RECT 4.000 69.040 273.485 77.840 ;
        RECT 4.400 67.640 273.085 69.040 ;
        RECT 4.000 58.840 273.485 67.640 ;
        RECT 4.000 57.440 273.085 58.840 ;
        RECT 4.000 55.440 273.485 57.440 ;
        RECT 4.400 54.040 273.485 55.440 ;
        RECT 4.000 48.640 273.485 54.040 ;
        RECT 4.000 47.240 273.085 48.640 ;
        RECT 4.000 45.240 273.485 47.240 ;
        RECT 4.400 43.840 273.485 45.240 ;
        RECT 4.000 35.040 273.485 43.840 ;
        RECT 4.400 33.640 273.085 35.040 ;
        RECT 4.000 24.840 273.485 33.640 ;
        RECT 4.000 23.440 273.085 24.840 ;
        RECT 4.000 21.440 273.485 23.440 ;
        RECT 4.400 20.040 273.485 21.440 ;
        RECT 4.000 14.640 273.485 20.040 ;
        RECT 4.000 13.240 273.085 14.640 ;
        RECT 4.000 11.240 273.485 13.240 ;
        RECT 4.400 9.840 273.485 11.240 ;
        RECT 4.000 1.040 273.485 9.840 ;
        RECT 4.000 0.175 273.085 1.040 ;
      LAYER met4 ;
        RECT 103.335 11.735 155.185 248.705 ;
  END
END pc
END LIBRARY

