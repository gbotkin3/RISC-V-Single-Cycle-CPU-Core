VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RISC_V
  CLASS BLOCK ;
  FOREIGN RISC_V ;
  ORIGIN 0.000 0.000 ;
  SIZE 1112.575 BY 1123.295 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END clk
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 1119.295 1040.430 1123.295 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 1119.295 914.850 1123.295 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.240 4.000 690.840 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 183.640 1112.575 184.240 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1003.040 4.000 1003.640 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 1119.295 460.830 1123.295 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 1119.295 393.210 1123.295 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 1119.295 766.730 1123.295 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 231.240 1112.575 231.840 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.070 1119.295 995.350 1123.295 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 340.040 1112.575 340.640 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 1119.295 1072.630 1123.295 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 918.040 4.000 918.640 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 1057.440 1112.575 1058.040 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 663.040 1112.575 663.640 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.190 0.000 982.470 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 1119.295 869.770 1123.295 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1122.040 4.000 1122.640 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 1119.295 438.290 1123.295 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 952.040 1112.575 952.640 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 387.640 1112.575 388.240 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1098.240 4.000 1098.840 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 1119.295 834.350 1123.295 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 805.840 1112.575 806.440 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 578.040 1112.575 578.640 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 0.000 1062.970 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 0.000 666.910 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 244.840 1112.575 245.440 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 1047.240 1112.575 1047.840 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 0.000 959.930 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 748.040 1112.575 748.640 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 1118.640 1112.575 1119.240 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 0.000 711.990 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 1119.295 293.390 1123.295 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 1119.295 267.630 1123.295 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 1119.295 573.530 1123.295 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.240 4.000 860.840 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 890.840 1112.575 891.440 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 530.440 1112.575 531.040 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 1119.295 64.770 1123.295 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.610 0.000 1017.890 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 125.840 1112.575 126.440 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 686.840 1112.575 687.440 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 1105.040 1112.575 1105.640 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 482.840 1112.575 483.440 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 999.640 1112.575 1000.240 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 1119.295 721.650 1123.295 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.240 4.000 894.840 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 0.000 937.390 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 1119.295 550.990 1123.295 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 0.000 769.950 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 1119.295 892.310 1123.295 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.030 0.000 1053.310 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 1119.295 654.030 1123.295 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 901.040 1112.575 901.640 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 1119.295 483.370 1123.295 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 567.840 1112.575 568.440 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 0.000 847.230 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 843.240 1112.575 843.840 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 829.640 1112.575 830.240 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 751.440 4.000 752.040 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 197.240 1112.575 197.840 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 1119.295 235.430 1123.295 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 0.000 869.770 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.770 0.000 1108.050 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 1119.295 42.230 1123.295 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 1071.040 1112.575 1071.640 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 1119.295 200.010 1123.295 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 975.840 1112.575 976.440 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 1119.295 303.050 1123.295 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 1119.295 87.310 1123.295 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 1119.295 177.470 1123.295 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 258.440 1112.575 259.040 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 1119.295 518.790 1123.295 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 1119.295 563.870 1123.295 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 88.440 1112.575 89.040 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 1119.295 666.910 1123.295 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 758.240 1112.575 758.840 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 54.440 1112.575 55.040 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.770 1119.295 1108.050 1123.295 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.240 4.000 656.840 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 1119.295 676.570 1123.295 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 1119.295 972.810 1123.295 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 924.840 1112.575 925.440 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 914.640 1112.575 915.240 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.840 4.000 500.440 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 1119.295 132.390 1123.295 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 0.000 950.270 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 1119.295 19.690 1123.295 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 1119.295 348.130 1123.295 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 1119.295 528.450 1123.295 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 411.440 1112.575 412.040 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 159.840 1112.575 160.440 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 1119.295 32.570 1123.295 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 112.240 1112.575 112.840 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.070 0.000 995.350 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 1119.295 937.390 1123.295 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.840 4.000 704.440 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 1119.295 109.850 1123.295 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1088.040 4.000 1088.640 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 1119.295 631.490 1123.295 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 1119.295 689.450 1123.295 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 221.040 1112.575 221.640 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 1009.840 1112.575 1010.440 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 0.000 892.310 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 377.440 1112.575 378.040 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 401.240 1112.575 401.840 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 0.000 702.330 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 282.240 1112.575 282.840 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 877.240 1112.575 877.840 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 724.240 1112.575 724.840 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 353.640 1112.575 354.240 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 1119.295 77.650 1123.295 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 605.240 1112.575 605.840 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 1119.295 699.110 1123.295 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 173.440 1112.575 174.040 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 1119.295 608.950 1123.295 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 1119.295 257.970 1123.295 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 710.640 1112.575 711.240 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 363.840 1112.575 364.440 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 1119.295 370.670 1123.295 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 1119.295 190.350 1123.295 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 78.240 1112.575 78.840 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 0.000 486.590 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.190 1119.295 982.470 1123.295 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 734.440 1112.575 735.040 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1111.840 4.000 1112.440 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 1119.295 280.510 1123.295 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 1119.295 950.270 1123.295 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 782.040 1112.575 782.640 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 965.640 4.000 966.240 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 1119.295 100.190 1123.295 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 1119.295 711.990 1123.295 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 0.000 914.850 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 448.840 1112.575 449.440 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 17.040 1112.575 17.640 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 1119.295 505.910 1123.295 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 1119.295 10.030 1123.295 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 149.640 1112.575 150.240 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.730 1119.295 1005.010 1123.295 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 1119.295 644.370 1123.295 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.810 1119.295 1050.090 1123.295 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 1119.295 212.890 1123.295 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 0.000 1098.390 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1050.640 4.000 1051.240 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 979.240 4.000 979.840 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 425.040 1112.575 425.640 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 316.240 1112.575 316.840 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 1119.295 406.090 1123.295 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 520.240 1112.575 520.840 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 0.000 779.610 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 0.000 757.070 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 0.000 905.190 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.240 4.000 775.840 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 0.000 824.690 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 846.640 4.000 847.240 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 1094.840 1112.575 1095.440 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 591.640 1112.575 592.240 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 1119.295 879.430 1123.295 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 1119.295 245.090 1123.295 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 962.240 1112.575 962.840 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 867.040 1112.575 867.640 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 1119.295 621.830 1123.295 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 513.440 4.000 514.040 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 1119.295 496.250 1123.295 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 1119.295 325.590 1123.295 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.230 0.000 1085.510 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 1081.240 1112.575 1081.840 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 64.640 1112.575 65.240 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 1119.295 541.330 1123.295 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.610 1119.295 1017.890 1123.295 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 931.640 4.000 932.240 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 472.640 1112.575 473.240 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1037.040 4.000 1037.640 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.750 0.000 815.030 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 0.000 1040.430 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 639.240 1112.575 639.840 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 1119.295 847.230 1123.295 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 506.640 1112.575 507.240 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.840 4.000 908.440 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 40.840 1112.575 41.440 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 1119.295 757.070 1123.295 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 0.000 972.810 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 1119.295 154.930 1123.295 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 496.440 1112.575 497.040 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 1119.295 55.110 1123.295 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 676.640 1112.575 677.240 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 0.000 1008.230 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 1119.295 428.630 1123.295 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.270 1119.295 1027.550 1123.295 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 795.640 1112.575 796.240 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 1119.295 383.550 1123.295 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 1119.295 473.710 1123.295 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 136.040 1112.575 136.640 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 608.640 4.000 609.240 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 1119.295 811.810 1123.295 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 1119.295 586.410 1123.295 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 1119.295 167.810 1123.295 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1074.440 4.000 1075.040 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 771.840 1112.575 772.440 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 700.440 1112.575 701.040 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 0.000 679.790 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 629.040 1112.575 629.640 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.490 0.000 1030.770 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 1119.295 779.610 1123.295 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.230 1119.295 1085.510 1123.295 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 207.440 1112.575 208.040 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 1119.295 222.550 1123.295 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 1119.295 451.170 1123.295 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 1033.640 1112.575 1034.240 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.230 1119.295 924.510 1123.295 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 435.240 1112.575 435.840 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 0.000 837.570 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 0.000 802.150 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.570 0.000 1075.850 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 268.640 1112.575 269.240 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 1119.295 415.750 1123.295 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 938.440 1112.575 939.040 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.840 4.000 942.440 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1026.840 4.000 1027.440 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 989.440 4.000 990.040 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 554.240 1112.575 554.840 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 0.000 621.830 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 1119.295 802.150 1123.295 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 1119.295 1062.970 1123.295 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 1119.295 122.730 1123.295 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 1119.295 1095.170 1123.295 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 329.840 1112.575 330.440 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 0.000 747.410 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 1119.295 959.930 1123.295 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 1119.295 315.930 1123.295 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 652.840 1112.575 653.440 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 0.000 882.650 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 306.040 1112.575 306.640 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 6.840 1112.575 7.440 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 459.040 1112.575 459.640 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.690 1119.295 901.970 1123.295 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 986.040 1112.575 986.640 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 30.640 1112.575 31.240 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 615.440 1112.575 616.040 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 1023.440 1112.575 1024.040 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 1119.295 856.890 1123.295 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 102.040 1112.575 102.640 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 1119.295 824.690 1123.295 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 0.000 724.870 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 0.000 860.110 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.240 4.000 1013.840 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 1119.295 338.470 1123.295 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 1119.295 596.070 1123.295 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 1119.295 361.010 1123.295 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 0.000 586.410 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 1119.295 789.270 1123.295 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 292.440 1112.575 293.040 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 853.440 1112.575 854.040 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 819.440 1112.575 820.040 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 1119.295 744.190 1123.295 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 1119.295 734.530 1123.295 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.240 4.000 1064.840 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 1119.295 145.270 1123.295 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 955.440 4.000 956.040 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.575 544.040 1112.575 544.640 ;
    END
  END la_oenb[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1110.000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1110.000 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1106.760 1109.845 ;
      LAYER met1 ;
        RECT 5.520 10.640 1106.760 1110.000 ;
      LAYER met2 ;
        RECT 6.990 1119.015 9.470 1119.295 ;
        RECT 10.310 1119.015 19.130 1119.295 ;
        RECT 19.970 1119.015 32.010 1119.295 ;
        RECT 32.850 1119.015 41.670 1119.295 ;
        RECT 42.510 1119.015 54.550 1119.295 ;
        RECT 55.390 1119.015 64.210 1119.295 ;
        RECT 65.050 1119.015 77.090 1119.295 ;
        RECT 77.930 1119.015 86.750 1119.295 ;
        RECT 87.590 1119.015 99.630 1119.295 ;
        RECT 100.470 1119.015 109.290 1119.295 ;
        RECT 110.130 1119.015 122.170 1119.295 ;
        RECT 123.010 1119.015 131.830 1119.295 ;
        RECT 132.670 1119.015 144.710 1119.295 ;
        RECT 145.550 1119.015 154.370 1119.295 ;
        RECT 155.210 1119.015 167.250 1119.295 ;
        RECT 168.090 1119.015 176.910 1119.295 ;
        RECT 177.750 1119.015 189.790 1119.295 ;
        RECT 190.630 1119.015 199.450 1119.295 ;
        RECT 200.290 1119.015 212.330 1119.295 ;
        RECT 213.170 1119.015 221.990 1119.295 ;
        RECT 222.830 1119.015 234.870 1119.295 ;
        RECT 235.710 1119.015 244.530 1119.295 ;
        RECT 245.370 1119.015 257.410 1119.295 ;
        RECT 258.250 1119.015 267.070 1119.295 ;
        RECT 267.910 1119.015 279.950 1119.295 ;
        RECT 280.790 1119.015 292.830 1119.295 ;
        RECT 293.670 1119.015 302.490 1119.295 ;
        RECT 303.330 1119.015 315.370 1119.295 ;
        RECT 316.210 1119.015 325.030 1119.295 ;
        RECT 325.870 1119.015 337.910 1119.295 ;
        RECT 338.750 1119.015 347.570 1119.295 ;
        RECT 348.410 1119.015 360.450 1119.295 ;
        RECT 361.290 1119.015 370.110 1119.295 ;
        RECT 370.950 1119.015 382.990 1119.295 ;
        RECT 383.830 1119.015 392.650 1119.295 ;
        RECT 393.490 1119.015 405.530 1119.295 ;
        RECT 406.370 1119.015 415.190 1119.295 ;
        RECT 416.030 1119.015 428.070 1119.295 ;
        RECT 428.910 1119.015 437.730 1119.295 ;
        RECT 438.570 1119.015 450.610 1119.295 ;
        RECT 451.450 1119.015 460.270 1119.295 ;
        RECT 461.110 1119.015 473.150 1119.295 ;
        RECT 473.990 1119.015 482.810 1119.295 ;
        RECT 483.650 1119.015 495.690 1119.295 ;
        RECT 496.530 1119.015 505.350 1119.295 ;
        RECT 506.190 1119.015 518.230 1119.295 ;
        RECT 519.070 1119.015 527.890 1119.295 ;
        RECT 528.730 1119.015 540.770 1119.295 ;
        RECT 541.610 1119.015 550.430 1119.295 ;
        RECT 551.270 1119.015 563.310 1119.295 ;
        RECT 564.150 1119.015 572.970 1119.295 ;
        RECT 573.810 1119.015 585.850 1119.295 ;
        RECT 586.690 1119.015 595.510 1119.295 ;
        RECT 596.350 1119.015 608.390 1119.295 ;
        RECT 609.230 1119.015 621.270 1119.295 ;
        RECT 622.110 1119.015 630.930 1119.295 ;
        RECT 631.770 1119.015 643.810 1119.295 ;
        RECT 644.650 1119.015 653.470 1119.295 ;
        RECT 654.310 1119.015 666.350 1119.295 ;
        RECT 667.190 1119.015 676.010 1119.295 ;
        RECT 676.850 1119.015 688.890 1119.295 ;
        RECT 689.730 1119.015 698.550 1119.295 ;
        RECT 699.390 1119.015 711.430 1119.295 ;
        RECT 712.270 1119.015 721.090 1119.295 ;
        RECT 721.930 1119.015 733.970 1119.295 ;
        RECT 734.810 1119.015 743.630 1119.295 ;
        RECT 744.470 1119.015 756.510 1119.295 ;
        RECT 757.350 1119.015 766.170 1119.295 ;
        RECT 767.010 1119.015 779.050 1119.295 ;
        RECT 779.890 1119.015 788.710 1119.295 ;
        RECT 789.550 1119.015 801.590 1119.295 ;
        RECT 802.430 1119.015 811.250 1119.295 ;
        RECT 812.090 1119.015 824.130 1119.295 ;
        RECT 824.970 1119.015 833.790 1119.295 ;
        RECT 834.630 1119.015 846.670 1119.295 ;
        RECT 847.510 1119.015 856.330 1119.295 ;
        RECT 857.170 1119.015 869.210 1119.295 ;
        RECT 870.050 1119.015 878.870 1119.295 ;
        RECT 879.710 1119.015 891.750 1119.295 ;
        RECT 892.590 1119.015 901.410 1119.295 ;
        RECT 902.250 1119.015 914.290 1119.295 ;
        RECT 915.130 1119.015 923.950 1119.295 ;
        RECT 924.790 1119.015 936.830 1119.295 ;
        RECT 937.670 1119.015 949.710 1119.295 ;
        RECT 950.550 1119.015 959.370 1119.295 ;
        RECT 960.210 1119.015 972.250 1119.295 ;
        RECT 973.090 1119.015 981.910 1119.295 ;
        RECT 982.750 1119.015 994.790 1119.295 ;
        RECT 995.630 1119.015 1004.450 1119.295 ;
        RECT 1005.290 1119.015 1017.330 1119.295 ;
        RECT 1018.170 1119.015 1026.990 1119.295 ;
        RECT 1027.830 1119.015 1039.870 1119.295 ;
        RECT 1040.710 1119.015 1049.530 1119.295 ;
        RECT 1050.370 1119.015 1062.410 1119.295 ;
        RECT 1063.250 1119.015 1072.070 1119.295 ;
        RECT 1072.910 1119.015 1084.950 1119.295 ;
        RECT 1085.790 1119.015 1094.610 1119.295 ;
        RECT 1095.450 1119.015 1103.910 1119.295 ;
        RECT 6.990 4.280 1103.910 1119.015 ;
        RECT 6.990 3.670 9.470 4.280 ;
        RECT 10.310 3.670 22.350 4.280 ;
        RECT 23.190 3.670 32.010 4.280 ;
        RECT 32.850 3.670 44.890 4.280 ;
        RECT 45.730 3.670 54.550 4.280 ;
        RECT 55.390 3.670 67.430 4.280 ;
        RECT 68.270 3.670 77.090 4.280 ;
        RECT 77.930 3.670 89.970 4.280 ;
        RECT 90.810 3.670 99.630 4.280 ;
        RECT 100.470 3.670 112.510 4.280 ;
        RECT 113.350 3.670 122.170 4.280 ;
        RECT 123.010 3.670 135.050 4.280 ;
        RECT 135.890 3.670 144.710 4.280 ;
        RECT 145.550 3.670 157.590 4.280 ;
        RECT 158.430 3.670 167.250 4.280 ;
        RECT 168.090 3.670 180.130 4.280 ;
        RECT 180.970 3.670 189.790 4.280 ;
        RECT 190.630 3.670 202.670 4.280 ;
        RECT 203.510 3.670 212.330 4.280 ;
        RECT 213.170 3.670 225.210 4.280 ;
        RECT 226.050 3.670 234.870 4.280 ;
        RECT 235.710 3.670 247.750 4.280 ;
        RECT 248.590 3.670 257.410 4.280 ;
        RECT 258.250 3.670 270.290 4.280 ;
        RECT 271.130 3.670 279.950 4.280 ;
        RECT 280.790 3.670 292.830 4.280 ;
        RECT 293.670 3.670 302.490 4.280 ;
        RECT 303.330 3.670 315.370 4.280 ;
        RECT 316.210 3.670 325.030 4.280 ;
        RECT 325.870 3.670 337.910 4.280 ;
        RECT 338.750 3.670 350.790 4.280 ;
        RECT 351.630 3.670 360.450 4.280 ;
        RECT 361.290 3.670 373.330 4.280 ;
        RECT 374.170 3.670 382.990 4.280 ;
        RECT 383.830 3.670 395.870 4.280 ;
        RECT 396.710 3.670 405.530 4.280 ;
        RECT 406.370 3.670 418.410 4.280 ;
        RECT 419.250 3.670 428.070 4.280 ;
        RECT 428.910 3.670 440.950 4.280 ;
        RECT 441.790 3.670 450.610 4.280 ;
        RECT 451.450 3.670 463.490 4.280 ;
        RECT 464.330 3.670 473.150 4.280 ;
        RECT 473.990 3.670 486.030 4.280 ;
        RECT 486.870 3.670 495.690 4.280 ;
        RECT 496.530 3.670 508.570 4.280 ;
        RECT 509.410 3.670 518.230 4.280 ;
        RECT 519.070 3.670 531.110 4.280 ;
        RECT 531.950 3.670 540.770 4.280 ;
        RECT 541.610 3.670 553.650 4.280 ;
        RECT 554.490 3.670 563.310 4.280 ;
        RECT 564.150 3.670 576.190 4.280 ;
        RECT 577.030 3.670 585.850 4.280 ;
        RECT 586.690 3.670 598.730 4.280 ;
        RECT 599.570 3.670 608.390 4.280 ;
        RECT 609.230 3.670 621.270 4.280 ;
        RECT 622.110 3.670 630.930 4.280 ;
        RECT 631.770 3.670 643.810 4.280 ;
        RECT 644.650 3.670 653.470 4.280 ;
        RECT 654.310 3.670 666.350 4.280 ;
        RECT 667.190 3.670 679.230 4.280 ;
        RECT 680.070 3.670 688.890 4.280 ;
        RECT 689.730 3.670 701.770 4.280 ;
        RECT 702.610 3.670 711.430 4.280 ;
        RECT 712.270 3.670 724.310 4.280 ;
        RECT 725.150 3.670 733.970 4.280 ;
        RECT 734.810 3.670 746.850 4.280 ;
        RECT 747.690 3.670 756.510 4.280 ;
        RECT 757.350 3.670 769.390 4.280 ;
        RECT 770.230 3.670 779.050 4.280 ;
        RECT 779.890 3.670 791.930 4.280 ;
        RECT 792.770 3.670 801.590 4.280 ;
        RECT 802.430 3.670 814.470 4.280 ;
        RECT 815.310 3.670 824.130 4.280 ;
        RECT 824.970 3.670 837.010 4.280 ;
        RECT 837.850 3.670 846.670 4.280 ;
        RECT 847.510 3.670 859.550 4.280 ;
        RECT 860.390 3.670 869.210 4.280 ;
        RECT 870.050 3.670 882.090 4.280 ;
        RECT 882.930 3.670 891.750 4.280 ;
        RECT 892.590 3.670 904.630 4.280 ;
        RECT 905.470 3.670 914.290 4.280 ;
        RECT 915.130 3.670 927.170 4.280 ;
        RECT 928.010 3.670 936.830 4.280 ;
        RECT 937.670 3.670 949.710 4.280 ;
        RECT 950.550 3.670 959.370 4.280 ;
        RECT 960.210 3.670 972.250 4.280 ;
        RECT 973.090 3.670 981.910 4.280 ;
        RECT 982.750 3.670 994.790 4.280 ;
        RECT 995.630 3.670 1007.670 4.280 ;
        RECT 1008.510 3.670 1017.330 4.280 ;
        RECT 1018.170 3.670 1030.210 4.280 ;
        RECT 1031.050 3.670 1039.870 4.280 ;
        RECT 1040.710 3.670 1052.750 4.280 ;
        RECT 1053.590 3.670 1062.410 4.280 ;
        RECT 1063.250 3.670 1075.290 4.280 ;
        RECT 1076.130 3.670 1084.950 4.280 ;
        RECT 1085.790 3.670 1097.830 4.280 ;
        RECT 1098.670 3.670 1103.910 4.280 ;
      LAYER met3 ;
        RECT 4.000 1118.240 1108.175 1119.105 ;
        RECT 4.000 1112.840 1108.575 1118.240 ;
        RECT 4.400 1111.440 1108.575 1112.840 ;
        RECT 4.000 1106.040 1108.575 1111.440 ;
        RECT 4.000 1104.640 1108.175 1106.040 ;
        RECT 4.000 1099.240 1108.575 1104.640 ;
        RECT 4.400 1097.840 1108.575 1099.240 ;
        RECT 4.000 1095.840 1108.575 1097.840 ;
        RECT 4.000 1094.440 1108.175 1095.840 ;
        RECT 4.000 1089.040 1108.575 1094.440 ;
        RECT 4.400 1087.640 1108.575 1089.040 ;
        RECT 4.000 1082.240 1108.575 1087.640 ;
        RECT 4.000 1080.840 1108.175 1082.240 ;
        RECT 4.000 1075.440 1108.575 1080.840 ;
        RECT 4.400 1074.040 1108.575 1075.440 ;
        RECT 4.000 1072.040 1108.575 1074.040 ;
        RECT 4.000 1070.640 1108.175 1072.040 ;
        RECT 4.000 1065.240 1108.575 1070.640 ;
        RECT 4.400 1063.840 1108.575 1065.240 ;
        RECT 4.000 1058.440 1108.575 1063.840 ;
        RECT 4.000 1057.040 1108.175 1058.440 ;
        RECT 4.000 1051.640 1108.575 1057.040 ;
        RECT 4.400 1050.240 1108.575 1051.640 ;
        RECT 4.000 1048.240 1108.575 1050.240 ;
        RECT 4.000 1046.840 1108.175 1048.240 ;
        RECT 4.000 1038.040 1108.575 1046.840 ;
        RECT 4.400 1036.640 1108.575 1038.040 ;
        RECT 4.000 1034.640 1108.575 1036.640 ;
        RECT 4.000 1033.240 1108.175 1034.640 ;
        RECT 4.000 1027.840 1108.575 1033.240 ;
        RECT 4.400 1026.440 1108.575 1027.840 ;
        RECT 4.000 1024.440 1108.575 1026.440 ;
        RECT 4.000 1023.040 1108.175 1024.440 ;
        RECT 4.000 1014.240 1108.575 1023.040 ;
        RECT 4.400 1012.840 1108.575 1014.240 ;
        RECT 4.000 1010.840 1108.575 1012.840 ;
        RECT 4.000 1009.440 1108.175 1010.840 ;
        RECT 4.000 1004.040 1108.575 1009.440 ;
        RECT 4.400 1002.640 1108.575 1004.040 ;
        RECT 4.000 1000.640 1108.575 1002.640 ;
        RECT 4.000 999.240 1108.175 1000.640 ;
        RECT 4.000 990.440 1108.575 999.240 ;
        RECT 4.400 989.040 1108.575 990.440 ;
        RECT 4.000 987.040 1108.575 989.040 ;
        RECT 4.000 985.640 1108.175 987.040 ;
        RECT 4.000 980.240 1108.575 985.640 ;
        RECT 4.400 978.840 1108.575 980.240 ;
        RECT 4.000 976.840 1108.575 978.840 ;
        RECT 4.000 975.440 1108.175 976.840 ;
        RECT 4.000 966.640 1108.575 975.440 ;
        RECT 4.400 965.240 1108.575 966.640 ;
        RECT 4.000 963.240 1108.575 965.240 ;
        RECT 4.000 961.840 1108.175 963.240 ;
        RECT 4.000 956.440 1108.575 961.840 ;
        RECT 4.400 955.040 1108.575 956.440 ;
        RECT 4.000 953.040 1108.575 955.040 ;
        RECT 4.000 951.640 1108.175 953.040 ;
        RECT 4.000 942.840 1108.575 951.640 ;
        RECT 4.400 941.440 1108.575 942.840 ;
        RECT 4.000 939.440 1108.575 941.440 ;
        RECT 4.000 938.040 1108.175 939.440 ;
        RECT 4.000 932.640 1108.575 938.040 ;
        RECT 4.400 931.240 1108.575 932.640 ;
        RECT 4.000 925.840 1108.575 931.240 ;
        RECT 4.000 924.440 1108.175 925.840 ;
        RECT 4.000 919.040 1108.575 924.440 ;
        RECT 4.400 917.640 1108.575 919.040 ;
        RECT 4.000 915.640 1108.575 917.640 ;
        RECT 4.000 914.240 1108.175 915.640 ;
        RECT 4.000 908.840 1108.575 914.240 ;
        RECT 4.400 907.440 1108.575 908.840 ;
        RECT 4.000 902.040 1108.575 907.440 ;
        RECT 4.000 900.640 1108.175 902.040 ;
        RECT 4.000 895.240 1108.575 900.640 ;
        RECT 4.400 893.840 1108.575 895.240 ;
        RECT 4.000 891.840 1108.575 893.840 ;
        RECT 4.000 890.440 1108.175 891.840 ;
        RECT 4.000 885.040 1108.575 890.440 ;
        RECT 4.400 883.640 1108.575 885.040 ;
        RECT 4.000 878.240 1108.575 883.640 ;
        RECT 4.000 876.840 1108.175 878.240 ;
        RECT 4.000 871.440 1108.575 876.840 ;
        RECT 4.400 870.040 1108.575 871.440 ;
        RECT 4.000 868.040 1108.575 870.040 ;
        RECT 4.000 866.640 1108.175 868.040 ;
        RECT 4.000 861.240 1108.575 866.640 ;
        RECT 4.400 859.840 1108.575 861.240 ;
        RECT 4.000 854.440 1108.575 859.840 ;
        RECT 4.000 853.040 1108.175 854.440 ;
        RECT 4.000 847.640 1108.575 853.040 ;
        RECT 4.400 846.240 1108.575 847.640 ;
        RECT 4.000 844.240 1108.575 846.240 ;
        RECT 4.000 842.840 1108.175 844.240 ;
        RECT 4.000 837.440 1108.575 842.840 ;
        RECT 4.400 836.040 1108.575 837.440 ;
        RECT 4.000 830.640 1108.575 836.040 ;
        RECT 4.000 829.240 1108.175 830.640 ;
        RECT 4.000 823.840 1108.575 829.240 ;
        RECT 4.400 822.440 1108.575 823.840 ;
        RECT 4.000 820.440 1108.575 822.440 ;
        RECT 4.000 819.040 1108.175 820.440 ;
        RECT 4.000 813.640 1108.575 819.040 ;
        RECT 4.400 812.240 1108.575 813.640 ;
        RECT 4.000 806.840 1108.575 812.240 ;
        RECT 4.000 805.440 1108.175 806.840 ;
        RECT 4.000 800.040 1108.575 805.440 ;
        RECT 4.400 798.640 1108.575 800.040 ;
        RECT 4.000 796.640 1108.575 798.640 ;
        RECT 4.000 795.240 1108.175 796.640 ;
        RECT 4.000 789.840 1108.575 795.240 ;
        RECT 4.400 788.440 1108.575 789.840 ;
        RECT 4.000 783.040 1108.575 788.440 ;
        RECT 4.000 781.640 1108.175 783.040 ;
        RECT 4.000 776.240 1108.575 781.640 ;
        RECT 4.400 774.840 1108.575 776.240 ;
        RECT 4.000 772.840 1108.575 774.840 ;
        RECT 4.000 771.440 1108.175 772.840 ;
        RECT 4.000 766.040 1108.575 771.440 ;
        RECT 4.400 764.640 1108.575 766.040 ;
        RECT 4.000 759.240 1108.575 764.640 ;
        RECT 4.000 757.840 1108.175 759.240 ;
        RECT 4.000 752.440 1108.575 757.840 ;
        RECT 4.400 751.040 1108.575 752.440 ;
        RECT 4.000 749.040 1108.575 751.040 ;
        RECT 4.000 747.640 1108.175 749.040 ;
        RECT 4.000 742.240 1108.575 747.640 ;
        RECT 4.400 740.840 1108.575 742.240 ;
        RECT 4.000 735.440 1108.575 740.840 ;
        RECT 4.000 734.040 1108.175 735.440 ;
        RECT 4.000 728.640 1108.575 734.040 ;
        RECT 4.400 727.240 1108.575 728.640 ;
        RECT 4.000 725.240 1108.575 727.240 ;
        RECT 4.000 723.840 1108.175 725.240 ;
        RECT 4.000 718.440 1108.575 723.840 ;
        RECT 4.400 717.040 1108.575 718.440 ;
        RECT 4.000 711.640 1108.575 717.040 ;
        RECT 4.000 710.240 1108.175 711.640 ;
        RECT 4.000 704.840 1108.575 710.240 ;
        RECT 4.400 703.440 1108.575 704.840 ;
        RECT 4.000 701.440 1108.575 703.440 ;
        RECT 4.000 700.040 1108.175 701.440 ;
        RECT 4.000 691.240 1108.575 700.040 ;
        RECT 4.400 689.840 1108.575 691.240 ;
        RECT 4.000 687.840 1108.575 689.840 ;
        RECT 4.000 686.440 1108.175 687.840 ;
        RECT 4.000 681.040 1108.575 686.440 ;
        RECT 4.400 679.640 1108.575 681.040 ;
        RECT 4.000 677.640 1108.575 679.640 ;
        RECT 4.000 676.240 1108.175 677.640 ;
        RECT 4.000 667.440 1108.575 676.240 ;
        RECT 4.400 666.040 1108.575 667.440 ;
        RECT 4.000 664.040 1108.575 666.040 ;
        RECT 4.000 662.640 1108.175 664.040 ;
        RECT 4.000 657.240 1108.575 662.640 ;
        RECT 4.400 655.840 1108.575 657.240 ;
        RECT 4.000 653.840 1108.575 655.840 ;
        RECT 4.000 652.440 1108.175 653.840 ;
        RECT 4.000 643.640 1108.575 652.440 ;
        RECT 4.400 642.240 1108.575 643.640 ;
        RECT 4.000 640.240 1108.575 642.240 ;
        RECT 4.000 638.840 1108.175 640.240 ;
        RECT 4.000 633.440 1108.575 638.840 ;
        RECT 4.400 632.040 1108.575 633.440 ;
        RECT 4.000 630.040 1108.575 632.040 ;
        RECT 4.000 628.640 1108.175 630.040 ;
        RECT 4.000 619.840 1108.575 628.640 ;
        RECT 4.400 618.440 1108.575 619.840 ;
        RECT 4.000 616.440 1108.575 618.440 ;
        RECT 4.000 615.040 1108.175 616.440 ;
        RECT 4.000 609.640 1108.575 615.040 ;
        RECT 4.400 608.240 1108.575 609.640 ;
        RECT 4.000 606.240 1108.575 608.240 ;
        RECT 4.000 604.840 1108.175 606.240 ;
        RECT 4.000 596.040 1108.575 604.840 ;
        RECT 4.400 594.640 1108.575 596.040 ;
        RECT 4.000 592.640 1108.575 594.640 ;
        RECT 4.000 591.240 1108.175 592.640 ;
        RECT 4.000 585.840 1108.575 591.240 ;
        RECT 4.400 584.440 1108.575 585.840 ;
        RECT 4.000 579.040 1108.575 584.440 ;
        RECT 4.000 577.640 1108.175 579.040 ;
        RECT 4.000 572.240 1108.575 577.640 ;
        RECT 4.400 570.840 1108.575 572.240 ;
        RECT 4.000 568.840 1108.575 570.840 ;
        RECT 4.000 567.440 1108.175 568.840 ;
        RECT 4.000 562.040 1108.575 567.440 ;
        RECT 4.400 560.640 1108.575 562.040 ;
        RECT 4.000 555.240 1108.575 560.640 ;
        RECT 4.000 553.840 1108.175 555.240 ;
        RECT 4.000 548.440 1108.575 553.840 ;
        RECT 4.400 547.040 1108.575 548.440 ;
        RECT 4.000 545.040 1108.575 547.040 ;
        RECT 4.000 543.640 1108.175 545.040 ;
        RECT 4.000 538.240 1108.575 543.640 ;
        RECT 4.400 536.840 1108.575 538.240 ;
        RECT 4.000 531.440 1108.575 536.840 ;
        RECT 4.000 530.040 1108.175 531.440 ;
        RECT 4.000 524.640 1108.575 530.040 ;
        RECT 4.400 523.240 1108.575 524.640 ;
        RECT 4.000 521.240 1108.575 523.240 ;
        RECT 4.000 519.840 1108.175 521.240 ;
        RECT 4.000 514.440 1108.575 519.840 ;
        RECT 4.400 513.040 1108.575 514.440 ;
        RECT 4.000 507.640 1108.575 513.040 ;
        RECT 4.000 506.240 1108.175 507.640 ;
        RECT 4.000 500.840 1108.575 506.240 ;
        RECT 4.400 499.440 1108.575 500.840 ;
        RECT 4.000 497.440 1108.575 499.440 ;
        RECT 4.000 496.040 1108.175 497.440 ;
        RECT 4.000 490.640 1108.575 496.040 ;
        RECT 4.400 489.240 1108.575 490.640 ;
        RECT 4.000 483.840 1108.575 489.240 ;
        RECT 4.000 482.440 1108.175 483.840 ;
        RECT 4.000 477.040 1108.575 482.440 ;
        RECT 4.400 475.640 1108.575 477.040 ;
        RECT 4.000 473.640 1108.575 475.640 ;
        RECT 4.000 472.240 1108.175 473.640 ;
        RECT 4.000 466.840 1108.575 472.240 ;
        RECT 4.400 465.440 1108.575 466.840 ;
        RECT 4.000 460.040 1108.575 465.440 ;
        RECT 4.000 458.640 1108.175 460.040 ;
        RECT 4.000 453.240 1108.575 458.640 ;
        RECT 4.400 451.840 1108.575 453.240 ;
        RECT 4.000 449.840 1108.575 451.840 ;
        RECT 4.000 448.440 1108.175 449.840 ;
        RECT 4.000 443.040 1108.575 448.440 ;
        RECT 4.400 441.640 1108.575 443.040 ;
        RECT 4.000 436.240 1108.575 441.640 ;
        RECT 4.000 434.840 1108.175 436.240 ;
        RECT 4.000 429.440 1108.575 434.840 ;
        RECT 4.400 428.040 1108.575 429.440 ;
        RECT 4.000 426.040 1108.575 428.040 ;
        RECT 4.000 424.640 1108.175 426.040 ;
        RECT 4.000 419.240 1108.575 424.640 ;
        RECT 4.400 417.840 1108.575 419.240 ;
        RECT 4.000 412.440 1108.575 417.840 ;
        RECT 4.000 411.040 1108.175 412.440 ;
        RECT 4.000 405.640 1108.575 411.040 ;
        RECT 4.400 404.240 1108.575 405.640 ;
        RECT 4.000 402.240 1108.575 404.240 ;
        RECT 4.000 400.840 1108.175 402.240 ;
        RECT 4.000 395.440 1108.575 400.840 ;
        RECT 4.400 394.040 1108.575 395.440 ;
        RECT 4.000 388.640 1108.575 394.040 ;
        RECT 4.000 387.240 1108.175 388.640 ;
        RECT 4.000 381.840 1108.575 387.240 ;
        RECT 4.400 380.440 1108.575 381.840 ;
        RECT 4.000 378.440 1108.575 380.440 ;
        RECT 4.000 377.040 1108.175 378.440 ;
        RECT 4.000 371.640 1108.575 377.040 ;
        RECT 4.400 370.240 1108.575 371.640 ;
        RECT 4.000 364.840 1108.575 370.240 ;
        RECT 4.000 363.440 1108.175 364.840 ;
        RECT 4.000 358.040 1108.575 363.440 ;
        RECT 4.400 356.640 1108.575 358.040 ;
        RECT 4.000 354.640 1108.575 356.640 ;
        RECT 4.000 353.240 1108.175 354.640 ;
        RECT 4.000 344.440 1108.575 353.240 ;
        RECT 4.400 343.040 1108.575 344.440 ;
        RECT 4.000 341.040 1108.575 343.040 ;
        RECT 4.000 339.640 1108.175 341.040 ;
        RECT 4.000 334.240 1108.575 339.640 ;
        RECT 4.400 332.840 1108.575 334.240 ;
        RECT 4.000 330.840 1108.575 332.840 ;
        RECT 4.000 329.440 1108.175 330.840 ;
        RECT 4.000 320.640 1108.575 329.440 ;
        RECT 4.400 319.240 1108.575 320.640 ;
        RECT 4.000 317.240 1108.575 319.240 ;
        RECT 4.000 315.840 1108.175 317.240 ;
        RECT 4.000 310.440 1108.575 315.840 ;
        RECT 4.400 309.040 1108.575 310.440 ;
        RECT 4.000 307.040 1108.575 309.040 ;
        RECT 4.000 305.640 1108.175 307.040 ;
        RECT 4.000 296.840 1108.575 305.640 ;
        RECT 4.400 295.440 1108.575 296.840 ;
        RECT 4.000 293.440 1108.575 295.440 ;
        RECT 4.000 292.040 1108.175 293.440 ;
        RECT 4.000 286.640 1108.575 292.040 ;
        RECT 4.400 285.240 1108.575 286.640 ;
        RECT 4.000 283.240 1108.575 285.240 ;
        RECT 4.000 281.840 1108.175 283.240 ;
        RECT 4.000 273.040 1108.575 281.840 ;
        RECT 4.400 271.640 1108.575 273.040 ;
        RECT 4.000 269.640 1108.575 271.640 ;
        RECT 4.000 268.240 1108.175 269.640 ;
        RECT 4.000 262.840 1108.575 268.240 ;
        RECT 4.400 261.440 1108.575 262.840 ;
        RECT 4.000 259.440 1108.575 261.440 ;
        RECT 4.000 258.040 1108.175 259.440 ;
        RECT 4.000 249.240 1108.575 258.040 ;
        RECT 4.400 247.840 1108.575 249.240 ;
        RECT 4.000 245.840 1108.575 247.840 ;
        RECT 4.000 244.440 1108.175 245.840 ;
        RECT 4.000 239.040 1108.575 244.440 ;
        RECT 4.400 237.640 1108.575 239.040 ;
        RECT 4.000 232.240 1108.575 237.640 ;
        RECT 4.000 230.840 1108.175 232.240 ;
        RECT 4.000 225.440 1108.575 230.840 ;
        RECT 4.400 224.040 1108.575 225.440 ;
        RECT 4.000 222.040 1108.575 224.040 ;
        RECT 4.000 220.640 1108.175 222.040 ;
        RECT 4.000 215.240 1108.575 220.640 ;
        RECT 4.400 213.840 1108.575 215.240 ;
        RECT 4.000 208.440 1108.575 213.840 ;
        RECT 4.000 207.040 1108.175 208.440 ;
        RECT 4.000 201.640 1108.575 207.040 ;
        RECT 4.400 200.240 1108.575 201.640 ;
        RECT 4.000 198.240 1108.575 200.240 ;
        RECT 4.000 196.840 1108.175 198.240 ;
        RECT 4.000 191.440 1108.575 196.840 ;
        RECT 4.400 190.040 1108.575 191.440 ;
        RECT 4.000 184.640 1108.575 190.040 ;
        RECT 4.000 183.240 1108.175 184.640 ;
        RECT 4.000 177.840 1108.575 183.240 ;
        RECT 4.400 176.440 1108.575 177.840 ;
        RECT 4.000 174.440 1108.575 176.440 ;
        RECT 4.000 173.040 1108.175 174.440 ;
        RECT 4.000 167.640 1108.575 173.040 ;
        RECT 4.400 166.240 1108.575 167.640 ;
        RECT 4.000 160.840 1108.575 166.240 ;
        RECT 4.000 159.440 1108.175 160.840 ;
        RECT 4.000 154.040 1108.575 159.440 ;
        RECT 4.400 152.640 1108.575 154.040 ;
        RECT 4.000 150.640 1108.575 152.640 ;
        RECT 4.000 149.240 1108.175 150.640 ;
        RECT 4.000 143.840 1108.575 149.240 ;
        RECT 4.400 142.440 1108.575 143.840 ;
        RECT 4.000 137.040 1108.575 142.440 ;
        RECT 4.000 135.640 1108.175 137.040 ;
        RECT 4.000 130.240 1108.575 135.640 ;
        RECT 4.400 128.840 1108.575 130.240 ;
        RECT 4.000 126.840 1108.575 128.840 ;
        RECT 4.000 125.440 1108.175 126.840 ;
        RECT 4.000 120.040 1108.575 125.440 ;
        RECT 4.400 118.640 1108.575 120.040 ;
        RECT 4.000 113.240 1108.575 118.640 ;
        RECT 4.000 111.840 1108.175 113.240 ;
        RECT 4.000 106.440 1108.575 111.840 ;
        RECT 4.400 105.040 1108.575 106.440 ;
        RECT 4.000 103.040 1108.575 105.040 ;
        RECT 4.000 101.640 1108.175 103.040 ;
        RECT 4.000 96.240 1108.575 101.640 ;
        RECT 4.400 94.840 1108.575 96.240 ;
        RECT 4.000 89.440 1108.575 94.840 ;
        RECT 4.000 88.040 1108.175 89.440 ;
        RECT 4.000 82.640 1108.575 88.040 ;
        RECT 4.400 81.240 1108.575 82.640 ;
        RECT 4.000 79.240 1108.575 81.240 ;
        RECT 4.000 77.840 1108.175 79.240 ;
        RECT 4.000 72.440 1108.575 77.840 ;
        RECT 4.400 71.040 1108.575 72.440 ;
        RECT 4.000 65.640 1108.575 71.040 ;
        RECT 4.000 64.240 1108.175 65.640 ;
        RECT 4.000 58.840 1108.575 64.240 ;
        RECT 4.400 57.440 1108.575 58.840 ;
        RECT 4.000 55.440 1108.575 57.440 ;
        RECT 4.000 54.040 1108.175 55.440 ;
        RECT 4.000 48.640 1108.575 54.040 ;
        RECT 4.400 47.240 1108.575 48.640 ;
        RECT 4.000 41.840 1108.575 47.240 ;
        RECT 4.000 40.440 1108.175 41.840 ;
        RECT 4.000 35.040 1108.575 40.440 ;
        RECT 4.400 33.640 1108.575 35.040 ;
        RECT 4.000 31.640 1108.575 33.640 ;
        RECT 4.000 30.240 1108.175 31.640 ;
        RECT 4.000 24.840 1108.575 30.240 ;
        RECT 4.400 23.440 1108.575 24.840 ;
        RECT 4.000 18.040 1108.575 23.440 ;
        RECT 4.000 16.640 1108.175 18.040 ;
        RECT 4.000 11.240 1108.575 16.640 ;
        RECT 4.400 10.375 1108.575 11.240 ;
      LAYER met4 ;
        RECT 138.295 11.735 174.240 1107.545 ;
        RECT 176.640 11.735 251.040 1107.545 ;
        RECT 253.440 11.735 327.840 1107.545 ;
        RECT 330.240 11.735 404.640 1107.545 ;
        RECT 407.040 11.735 481.440 1107.545 ;
        RECT 483.840 11.735 558.240 1107.545 ;
        RECT 560.640 11.735 635.040 1107.545 ;
        RECT 637.440 11.735 711.840 1107.545 ;
        RECT 714.240 11.735 788.640 1107.545 ;
        RECT 791.040 11.735 801.025 1107.545 ;
  END
END RISC_V
END LIBRARY

