magic
tech sky130B
magscale 1 2
timestamp 1663699768
<< obsli1 >>
rect 1104 2159 48852 47345
<< obsm1 >>
rect 14 2128 48852 47376
<< metal2 >>
rect 7746 49200 7802 50000
rect 17406 49200 17462 50000
rect 26422 49200 26478 50000
rect 36082 49200 36138 50000
rect 45098 49200 45154 50000
rect 18 0 74 800
rect 9034 0 9090 800
rect 18050 0 18106 800
rect 27710 0 27766 800
rect 36726 0 36782 800
rect 46386 0 46442 800
<< obsm2 >>
rect 20 49144 7690 49314
rect 7858 49144 17350 49314
rect 17518 49144 26366 49314
rect 26534 49144 36026 49314
rect 36194 49144 45042 49314
rect 45210 49144 48190 49314
rect 20 856 48190 49144
rect 130 800 8978 856
rect 9146 800 17994 856
rect 18162 800 27654 856
rect 27822 800 36670 856
rect 36838 800 46330 856
rect 46498 800 48190 856
<< metal3 >>
rect 0 48968 800 49088
rect 49200 44888 50000 45008
rect 0 38768 800 38888
rect 49200 35368 50000 35488
rect 0 29248 800 29368
rect 49200 25168 50000 25288
rect 0 19048 800 19168
rect 49200 15648 50000 15768
rect 0 9528 800 9648
rect 49200 5448 50000 5568
<< obsm3 >>
rect 880 48888 49200 49061
rect 800 45088 49200 48888
rect 800 44808 49120 45088
rect 800 38968 49200 44808
rect 880 38688 49200 38968
rect 800 35568 49200 38688
rect 800 35288 49120 35568
rect 800 29448 49200 35288
rect 880 29168 49200 29448
rect 800 25368 49200 29168
rect 800 25088 49120 25368
rect 800 19248 49200 25088
rect 880 18968 49200 19248
rect 800 15848 49200 18968
rect 800 15568 49120 15848
rect 800 9728 49200 15568
rect 880 9448 49200 9728
rect 800 5648 49200 9448
rect 800 5368 49120 5648
rect 800 2143 49200 5368
<< metal4 >>
rect 4208 2128 4528 47376
rect 19568 2128 19888 47376
rect 34928 2128 35248 47376
<< labels >>
rlabel metal2 s 36726 0 36782 800 6 branch_output
port 1 nsew signal output
rlabel metal3 s 49200 44888 50000 45008 6 clk
port 2 nsew signal input
rlabel metal2 s 45098 49200 45154 50000 6 immediate_sel_output
port 3 nsew signal output
rlabel metal2 s 26422 49200 26478 50000 6 instruction_type[0]
port 4 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 instruction_type[1]
port 5 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 instruction_type[2]
port 6 nsew signal input
rlabel metal3 s 49200 5448 50000 5568 6 instruction_type[3]
port 7 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 instruction_type[4]
port 8 nsew signal input
rlabel metal3 s 49200 35368 50000 35488 6 instruction_type[5]
port 9 nsew signal input
rlabel metal2 s 18 0 74 800 6 jump_jal_output
port 10 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 jump_jalr_output
port 11 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 mem_write_output
port 12 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 opcode[0]
port 13 nsew signal input
rlabel metal2 s 17406 49200 17462 50000 6 opcode[1]
port 14 nsew signal input
rlabel metal3 s 49200 25168 50000 25288 6 opcode[2]
port 15 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 opcode[3]
port 16 nsew signal input
rlabel metal2 s 36082 49200 36138 50000 6 opcode[4]
port 17 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 opcode[5]
port 18 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 opcode[6]
port 19 nsew signal input
rlabel metal2 s 7746 49200 7802 50000 6 reg_write_output
port 20 nsew signal output
rlabel metal3 s 49200 15648 50000 15768 6 rst_n
port 21 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 22 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 22 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 23 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 50000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 769662
string GDS_FILE /home/drewarosa/RISC-V-Single-Cycle-CPU-Core/openlane/control/runs/22_09_20_14_48/results/signoff/control.magic.gds
string GDS_START 97384
<< end >>

