magic
tech sky130B
magscale 1 2
timestamp 1663699925
<< viali >>
rect 6469 47209 6503 47243
rect 13461 47209 13495 47243
rect 15117 47209 15151 47243
rect 19625 47209 19659 47243
rect 21189 47209 21223 47243
rect 26433 47209 26467 47243
rect 34069 47209 34103 47243
rect 37473 47209 37507 47243
rect 38301 47209 38335 47243
rect 40233 47209 40267 47243
rect 40785 47209 40819 47243
rect 42809 47209 42843 47243
rect 46673 47209 46707 47243
rect 4169 47141 4203 47175
rect 12173 47141 12207 47175
rect 23305 47141 23339 47175
rect 27721 47141 27755 47175
rect 30941 47141 30975 47175
rect 33517 47141 33551 47175
rect 36093 47141 36127 47175
rect 1961 47073 1995 47107
rect 9781 47073 9815 47107
rect 10057 47073 10091 47107
rect 12725 47073 12759 47107
rect 14473 47073 14507 47107
rect 17785 47073 17819 47107
rect 29561 47073 29595 47107
rect 2237 47005 2271 47039
rect 3985 47005 4019 47039
rect 4629 47005 4663 47039
rect 6653 47005 6687 47039
rect 7389 47005 7423 47039
rect 7849 47005 7883 47039
rect 11989 47005 12023 47039
rect 13277 47005 13311 47039
rect 14289 47005 14323 47039
rect 14933 47005 14967 47039
rect 15761 47005 15795 47039
rect 15853 47005 15887 47039
rect 17049 47005 17083 47039
rect 17509 47005 17543 47039
rect 19441 47005 19475 47039
rect 21925 47005 21959 47039
rect 22201 47005 22235 47039
rect 23489 47005 23523 47039
rect 24409 47005 24443 47039
rect 24593 47005 24627 47039
rect 25053 47005 25087 47039
rect 29837 47005 29871 47039
rect 32137 47005 32171 47039
rect 34713 47005 34747 47039
rect 36645 47005 36679 47039
rect 37289 47005 37323 47039
rect 38945 47005 38979 47039
rect 40877 47005 40911 47039
rect 42625 47005 42659 47039
rect 46489 47005 46523 47039
rect 48053 47005 48087 47039
rect 2789 46937 2823 46971
rect 2973 46937 3007 46971
rect 9321 46937 9355 46971
rect 20361 46937 20395 46971
rect 20913 46937 20947 46971
rect 22017 46937 22051 46971
rect 22385 46937 22419 46971
rect 24501 46937 24535 46971
rect 25320 46937 25354 46971
rect 29009 46937 29043 46971
rect 32382 46937 32416 46971
rect 34980 46937 35014 46971
rect 45385 46937 45419 46971
rect 45569 46937 45603 46971
rect 47869 46937 47903 46971
rect 8033 46869 8067 46903
rect 14105 46869 14139 46903
rect 16037 46869 16071 46903
rect 38761 46869 38795 46903
rect 2513 46665 2547 46699
rect 3065 46665 3099 46699
rect 10425 46665 10459 46699
rect 21097 46665 21131 46699
rect 24409 46665 24443 46699
rect 30481 46665 30515 46699
rect 34253 46665 34287 46699
rect 42441 46665 42475 46699
rect 45201 46665 45235 46699
rect 11805 46597 11839 46631
rect 13001 46597 13035 46631
rect 14657 46597 14691 46631
rect 18153 46597 18187 46631
rect 19809 46597 19843 46631
rect 35265 46597 35299 46631
rect 46949 46597 46983 46631
rect 1409 46529 1443 46563
rect 12909 46529 12943 46563
rect 13093 46529 13127 46563
rect 13737 46529 13771 46563
rect 14565 46529 14599 46563
rect 14749 46529 14783 46563
rect 15393 46529 15427 46563
rect 16865 46529 16899 46563
rect 18061 46529 18095 46563
rect 18245 46529 18279 46563
rect 18889 46529 18923 46563
rect 19717 46529 19751 46563
rect 19993 46529 20027 46563
rect 20913 46529 20947 46563
rect 21097 46529 21131 46563
rect 21925 46529 21959 46563
rect 23857 46529 23891 46563
rect 24317 46529 24351 46563
rect 24501 46529 24535 46563
rect 24961 46529 24995 46563
rect 25228 46529 25262 46563
rect 27261 46529 27295 46563
rect 28365 46529 28399 46563
rect 31401 46529 31435 46563
rect 32137 46529 32171 46563
rect 32404 46529 32438 46563
rect 34069 46529 34103 46563
rect 48053 46529 48087 46563
rect 8769 46461 8803 46495
rect 13645 46461 13679 46495
rect 15301 46461 15335 46495
rect 15761 46461 15795 46495
rect 16773 46461 16807 46495
rect 18797 46461 18831 46495
rect 19257 46461 19291 46495
rect 22937 46461 22971 46495
rect 26985 46461 27019 46495
rect 28641 46461 28675 46495
rect 47869 46461 47903 46495
rect 9873 46393 9907 46427
rect 10977 46393 11011 46427
rect 17233 46393 17267 46427
rect 19993 46393 20027 46427
rect 23397 46393 23431 46427
rect 35081 46393 35115 46427
rect 46765 46393 46799 46427
rect 1593 46325 1627 46359
rect 6837 46325 6871 46359
rect 9321 46325 9355 46359
rect 12449 46325 12483 46359
rect 14013 46325 14047 46359
rect 23765 46325 23799 46359
rect 26341 46325 26375 46359
rect 29929 46325 29963 46359
rect 31585 46325 31619 46359
rect 33517 46325 33551 46359
rect 35909 46325 35943 46359
rect 46213 46325 46247 46359
rect 2513 46121 2547 46155
rect 9137 46121 9171 46155
rect 12909 46121 12943 46155
rect 13461 46121 13495 46155
rect 16313 46121 16347 46155
rect 18705 46121 18739 46155
rect 19901 46121 19935 46155
rect 33517 46121 33551 46155
rect 34069 46121 34103 46155
rect 34897 46121 34931 46155
rect 46673 46121 46707 46155
rect 21741 46053 21775 46087
rect 47225 46053 47259 46087
rect 12449 45985 12483 46019
rect 19625 45985 19659 46019
rect 20913 45985 20947 46019
rect 22017 45985 22051 46019
rect 22293 45985 22327 46019
rect 23305 45985 23339 46019
rect 25605 45985 25639 46019
rect 31401 45985 31435 46019
rect 1869 45917 1903 45951
rect 14105 45917 14139 45951
rect 14289 45917 14323 45951
rect 14565 45917 14599 45951
rect 16497 45917 16531 45951
rect 16773 45917 16807 45951
rect 17693 45917 17727 45951
rect 17877 45917 17911 45951
rect 19717 45917 19751 45951
rect 21097 45917 21131 45951
rect 21925 45917 21959 45951
rect 22385 45917 22419 45951
rect 23673 45917 23707 45951
rect 24501 45917 24535 45951
rect 24685 45917 24719 45951
rect 25861 45917 25895 45951
rect 27537 45917 27571 45951
rect 30021 45917 30055 45951
rect 30297 45917 30331 45951
rect 32137 45917 32171 45951
rect 48053 45917 48087 45951
rect 14381 45849 14415 45883
rect 14473 45849 14507 45883
rect 14749 45849 14783 45883
rect 16681 45849 16715 45883
rect 18337 45849 18371 45883
rect 18521 45849 18555 45883
rect 21281 45849 21315 45883
rect 23581 45849 23615 45883
rect 23857 45849 23891 45883
rect 24409 45849 24443 45883
rect 24869 45849 24903 45883
rect 27804 45849 27838 45883
rect 32382 45849 32416 45883
rect 47869 45849 47903 45883
rect 1961 45781 1995 45815
rect 9689 45781 9723 45815
rect 10241 45781 10275 45815
rect 10793 45781 10827 45815
rect 11253 45781 11287 45815
rect 11897 45781 11931 45815
rect 15853 45781 15887 45815
rect 17785 45781 17819 45815
rect 19257 45781 19291 45815
rect 20453 45781 20487 45815
rect 22201 45781 22235 45815
rect 23489 45781 23523 45815
rect 26985 45781 27019 45815
rect 28917 45781 28951 45815
rect 1685 45577 1719 45611
rect 16957 45577 16991 45611
rect 26157 45577 26191 45611
rect 31493 45577 31527 45611
rect 48053 45577 48087 45611
rect 9689 45509 9723 45543
rect 11897 45509 11931 45543
rect 12541 45509 12575 45543
rect 13185 45509 13219 45543
rect 20913 45509 20947 45543
rect 21971 45509 22005 45543
rect 22201 45509 22235 45543
rect 30941 45509 30975 45543
rect 13001 45441 13035 45475
rect 13277 45441 13311 45475
rect 13921 45441 13955 45475
rect 15485 45441 15519 45475
rect 16681 45441 16715 45475
rect 17417 45441 17451 45475
rect 17601 45441 17635 45475
rect 18245 45441 18279 45475
rect 18337 45441 18371 45475
rect 18521 45441 18555 45475
rect 19349 45441 19383 45475
rect 21097 45441 21131 45475
rect 21281 45441 21315 45475
rect 22109 45441 22143 45475
rect 22293 45441 22327 45475
rect 23121 45441 23155 45475
rect 24133 45441 24167 45475
rect 25251 45441 25285 45475
rect 25973 45441 26007 45475
rect 26249 45441 26283 45475
rect 27169 45441 27203 45475
rect 29653 45441 29687 45475
rect 29929 45441 29963 45475
rect 33250 45441 33284 45475
rect 33517 45441 33551 45475
rect 34621 45441 34655 45475
rect 34805 45441 34839 45475
rect 35265 45441 35299 45475
rect 13829 45373 13863 45407
rect 14289 45373 14323 45407
rect 15577 45373 15611 45407
rect 16957 45373 16991 45407
rect 17509 45373 17543 45407
rect 18981 45373 19015 45407
rect 19441 45373 19475 45407
rect 21833 45373 21867 45407
rect 22477 45373 22511 45407
rect 23029 45373 23063 45407
rect 24041 45373 24075 45407
rect 25421 45373 25455 45407
rect 34713 45373 34747 45407
rect 13001 45305 13035 45339
rect 15853 45305 15887 45339
rect 16773 45305 16807 45339
rect 18521 45305 18555 45339
rect 24501 45305 24535 45339
rect 25973 45305 26007 45339
rect 27353 45305 27387 45339
rect 32137 45305 32171 45339
rect 10425 45237 10459 45271
rect 10977 45237 11011 45271
rect 14749 45237 14783 45271
rect 20453 45237 20487 45271
rect 23489 45237 23523 45271
rect 25053 45237 25087 45271
rect 28365 45237 28399 45271
rect 30481 45237 30515 45271
rect 34069 45237 34103 45271
rect 13001 45033 13035 45067
rect 14749 45033 14783 45067
rect 16037 45033 16071 45067
rect 17509 45033 17543 45067
rect 22109 45033 22143 45067
rect 22661 45033 22695 45067
rect 24777 45033 24811 45067
rect 26249 45033 26283 45067
rect 28457 45033 28491 45067
rect 48145 45033 48179 45067
rect 18061 44965 18095 44999
rect 19993 44965 20027 44999
rect 16589 44897 16623 44931
rect 17049 44897 17083 44931
rect 21649 44897 21683 44931
rect 27077 44897 27111 44931
rect 31217 44897 31251 44931
rect 35541 44897 35575 44931
rect 10609 44829 10643 44863
rect 12817 44829 12851 44863
rect 13001 44829 13035 44863
rect 14129 44829 14163 44863
rect 14289 44829 14323 44863
rect 14400 44826 14434 44860
rect 14519 44829 14553 44863
rect 15301 44829 15335 44863
rect 15485 44829 15519 44863
rect 16674 44829 16708 44863
rect 19257 44829 19291 44863
rect 19441 44829 19475 44863
rect 20545 44829 20579 44863
rect 20729 44829 20763 44863
rect 20913 44829 20947 44863
rect 21741 44829 21775 44863
rect 22569 44829 22603 44863
rect 22753 44829 22787 44863
rect 24961 44829 24995 44863
rect 25053 44829 25087 44863
rect 30941 44829 30975 44863
rect 33701 44829 33735 44863
rect 34897 44829 34931 44863
rect 11713 44761 11747 44795
rect 12357 44761 12391 44795
rect 15393 44761 15427 44795
rect 20821 44761 20855 44795
rect 25697 44761 25731 44795
rect 27344 44761 27378 44795
rect 29561 44761 29595 44795
rect 34713 44761 34747 44795
rect 10057 44693 10091 44727
rect 11253 44693 11287 44727
rect 13553 44693 13587 44727
rect 18613 44693 18647 44727
rect 19349 44693 19383 44727
rect 21097 44693 21131 44727
rect 23305 44693 23339 44727
rect 23765 44693 23799 44727
rect 32137 44693 32171 44727
rect 33241 44693 33275 44727
rect 35081 44693 35115 44727
rect 36093 44693 36127 44727
rect 9873 44489 9907 44523
rect 11897 44489 11931 44523
rect 12725 44489 12759 44523
rect 13277 44489 13311 44523
rect 16037 44489 16071 44523
rect 19901 44489 19935 44523
rect 32229 44489 32263 44523
rect 34345 44489 34379 44523
rect 47961 44489 47995 44523
rect 19441 44421 19475 44455
rect 1409 44353 1443 44387
rect 12541 44353 12575 44387
rect 13185 44353 13219 44387
rect 13369 44353 13403 44387
rect 15209 44353 15243 44387
rect 15393 44353 15427 44387
rect 15577 44353 15611 44387
rect 16865 44353 16899 44387
rect 17509 44353 17543 44387
rect 18061 44353 18095 44387
rect 18153 44353 18187 44387
rect 18337 44353 18371 44387
rect 19257 44353 19291 44387
rect 20085 44353 20119 44387
rect 20269 44353 20303 44387
rect 20729 44353 20763 44387
rect 20913 44353 20947 44387
rect 21833 44353 21867 44387
rect 22017 44353 22051 44387
rect 23765 44353 23799 44387
rect 23949 44353 23983 44387
rect 24593 44353 24627 44387
rect 28282 44353 28316 44387
rect 28549 44353 28583 44387
rect 29285 44353 29319 44387
rect 33342 44353 33376 44387
rect 33609 44353 33643 44387
rect 34529 44353 34563 44387
rect 35449 44353 35483 44387
rect 35541 44353 35575 44387
rect 48053 44353 48087 44387
rect 12357 44285 12391 44319
rect 16681 44285 16715 44319
rect 18981 44285 19015 44319
rect 22293 44285 22327 44319
rect 23305 44285 23339 44319
rect 24777 44285 24811 44319
rect 29009 44285 29043 44319
rect 30665 44285 30699 44319
rect 34805 44285 34839 44319
rect 10425 44217 10459 44251
rect 14657 44217 14691 44251
rect 17049 44217 17083 44251
rect 19073 44217 19107 44251
rect 27169 44217 27203 44251
rect 34713 44217 34747 44251
rect 36185 44217 36219 44251
rect 1593 44149 1627 44183
rect 9321 44149 9355 44183
rect 10977 44149 11011 44183
rect 14105 44149 14139 44183
rect 18521 44149 18555 44183
rect 20821 44149 20855 44183
rect 22201 44149 22235 44183
rect 23949 44149 23983 44183
rect 24409 44149 24443 44183
rect 25421 44149 25455 44183
rect 26065 44149 26099 44183
rect 31493 44149 31527 44183
rect 35265 44149 35299 44183
rect 36737 44149 36771 44183
rect 37381 44149 37415 44183
rect 37933 44149 37967 44183
rect 1409 43945 1443 43979
rect 12449 43945 12483 43979
rect 14473 43945 14507 43979
rect 16957 43945 16991 43979
rect 25605 43945 25639 43979
rect 35909 43945 35943 43979
rect 48053 43945 48087 43979
rect 13553 43877 13587 43911
rect 17601 43877 17635 43911
rect 24777 43877 24811 43911
rect 13093 43809 13127 43843
rect 15761 43809 15795 43843
rect 24869 43809 24903 43843
rect 27353 43809 27387 43843
rect 10885 43741 10919 43775
rect 11437 43741 11471 43775
rect 13185 43741 13219 43775
rect 14933 43741 14967 43775
rect 15117 43741 15151 43775
rect 16313 43741 16347 43775
rect 16497 43741 16531 43775
rect 18061 43741 18095 43775
rect 18245 43741 18279 43775
rect 18337 43741 18371 43775
rect 18429 43741 18463 43775
rect 19625 43741 19659 43775
rect 20545 43741 20579 43775
rect 20729 43741 20763 43775
rect 21557 43741 21591 43775
rect 22109 43741 22143 43775
rect 22293 43741 22327 43775
rect 23581 43741 23615 43775
rect 23673 43741 23707 43775
rect 23784 43741 23818 43775
rect 24593 43741 24627 43775
rect 25329 43741 25363 43775
rect 26893 43741 26927 43775
rect 27629 43741 27663 43775
rect 33977 43741 34011 43775
rect 34897 43741 34931 43775
rect 35173 43741 35207 43775
rect 35633 43741 35667 43775
rect 36369 43741 36403 43775
rect 37565 43741 37599 43775
rect 10333 43673 10367 43707
rect 16405 43673 16439 43707
rect 18705 43673 18739 43707
rect 19717 43673 19751 43707
rect 19901 43673 19935 43707
rect 21189 43673 21223 43707
rect 21373 43673 21407 43707
rect 23867 43673 23901 43707
rect 25513 43673 25547 43707
rect 26249 43673 26283 43707
rect 31217 43673 31251 43707
rect 35081 43673 35115 43707
rect 35725 43673 35759 43707
rect 35909 43673 35943 43707
rect 36461 43673 36495 43707
rect 36645 43673 36679 43707
rect 37749 43673 37783 43707
rect 9781 43605 9815 43639
rect 11897 43605 11931 43639
rect 15117 43605 15151 43639
rect 19809 43605 19843 43639
rect 20637 43605 20671 43639
rect 22293 43605 22327 43639
rect 23121 43605 23155 43639
rect 24409 43605 24443 43639
rect 28733 43605 28767 43639
rect 29653 43605 29687 43639
rect 30297 43605 30331 43639
rect 32505 43605 32539 43639
rect 33425 43605 33459 43639
rect 34713 43605 34747 43639
rect 36369 43605 36403 43639
rect 37933 43605 37967 43639
rect 38393 43605 38427 43639
rect 38945 43605 38979 43639
rect 10885 43401 10919 43435
rect 12909 43401 12943 43435
rect 13921 43401 13955 43435
rect 18981 43401 19015 43435
rect 22477 43401 22511 43435
rect 23581 43401 23615 43435
rect 28089 43401 28123 43435
rect 29101 43401 29135 43435
rect 35449 43401 35483 43435
rect 36001 43401 36035 43435
rect 20913 43333 20947 43367
rect 26188 43333 26222 43367
rect 30389 43333 30423 43367
rect 34314 43333 34348 43367
rect 12725 43265 12759 43299
rect 12909 43265 12943 43299
rect 13553 43265 13587 43299
rect 13737 43265 13771 43299
rect 14657 43265 14691 43299
rect 15761 43265 15795 43299
rect 16681 43265 16715 43299
rect 16865 43265 16899 43299
rect 17417 43265 17451 43299
rect 17509 43265 17543 43299
rect 17693 43265 17727 43299
rect 18337 43265 18371 43299
rect 18521 43265 18555 43299
rect 18632 43265 18666 43299
rect 18725 43265 18759 43299
rect 19809 43265 19843 43299
rect 20545 43265 20579 43299
rect 20729 43265 20763 43299
rect 21005 43265 21039 43299
rect 22017 43265 22051 43299
rect 22109 43265 22143 43299
rect 23121 43265 23155 43299
rect 23397 43265 23431 43299
rect 24041 43265 24075 43299
rect 24133 43265 24167 43299
rect 24244 43265 24278 43299
rect 24409 43265 24443 43299
rect 26433 43265 26467 43299
rect 33342 43265 33376 43299
rect 33609 43265 33643 43299
rect 34069 43265 34103 43299
rect 36277 43265 36311 43299
rect 36369 43265 36403 43299
rect 37749 43265 37783 43299
rect 37933 43265 37967 43299
rect 38393 43265 38427 43299
rect 38577 43265 38611 43299
rect 9873 43197 9907 43231
rect 10425 43197 10459 43231
rect 13461 43197 13495 43231
rect 13645 43197 13679 43231
rect 14749 43197 14783 43231
rect 15669 43197 15703 43231
rect 17877 43197 17911 43231
rect 19625 43197 19659 43231
rect 19717 43197 19751 43231
rect 19901 43197 19935 43231
rect 26985 43197 27019 43231
rect 36185 43197 36219 43231
rect 36461 43197 36495 43231
rect 11713 43129 11747 43163
rect 15025 43129 15059 43163
rect 16129 43129 16163 43163
rect 20085 43129 20119 43163
rect 23213 43129 23247 43163
rect 24593 43129 24627 43163
rect 40141 43129 40175 43163
rect 12265 43061 12299 43095
rect 16773 43061 16807 43095
rect 21833 43061 21867 43095
rect 25053 43061 25087 43095
rect 27629 43061 27663 43095
rect 30849 43061 30883 43095
rect 31401 43061 31435 43095
rect 32229 43061 32263 43095
rect 37841 43061 37875 43095
rect 38485 43061 38519 43095
rect 39129 43061 39163 43095
rect 39681 43061 39715 43095
rect 10149 42857 10183 42891
rect 10701 42857 10735 42891
rect 12817 42857 12851 42891
rect 15761 42857 15795 42891
rect 18061 42857 18095 42891
rect 19717 42857 19751 42891
rect 20453 42857 20487 42891
rect 21465 42857 21499 42891
rect 21649 42857 21683 42891
rect 33977 42857 34011 42891
rect 40417 42857 40451 42891
rect 12357 42721 12391 42755
rect 13553 42721 13587 42755
rect 15853 42721 15887 42755
rect 20361 42721 20395 42755
rect 23489 42721 23523 42755
rect 25513 42721 25547 42755
rect 27353 42721 27387 42755
rect 29561 42721 29595 42755
rect 33333 42721 33367 42755
rect 34713 42721 34747 42755
rect 35081 42721 35115 42755
rect 37013 42721 37047 42755
rect 37289 42721 37323 42755
rect 38117 42721 38151 42755
rect 38301 42721 38335 42755
rect 1685 42653 1719 42687
rect 2237 42653 2271 42687
rect 12449 42653 12483 42687
rect 14841 42653 14875 42687
rect 15577 42653 15611 42687
rect 16957 42653 16991 42687
rect 17969 42653 18003 42687
rect 18153 42653 18187 42687
rect 19349 42653 19383 42687
rect 19441 42653 19475 42687
rect 19533 42653 19567 42687
rect 20637 42653 20671 42687
rect 21281 42653 21315 42687
rect 21557 42653 21591 42687
rect 21741 42653 21775 42687
rect 23673 42653 23707 42687
rect 23857 42653 23891 42687
rect 24593 42653 24627 42687
rect 24777 42653 24811 42687
rect 24869 42653 24903 42687
rect 25329 42653 25363 42687
rect 25697 42653 25731 42687
rect 27629 42653 27663 42687
rect 29837 42653 29871 42687
rect 33057 42653 33091 42687
rect 34897 42653 34931 42687
rect 35173 42653 35207 42687
rect 35265 42653 35299 42687
rect 35449 42653 35483 42687
rect 35909 42653 35943 42687
rect 36277 42653 36311 42687
rect 36369 42653 36403 42687
rect 37381 42653 37415 42687
rect 38025 42653 38059 42687
rect 47501 42653 47535 42687
rect 48145 42653 48179 42687
rect 16773 42585 16807 42619
rect 17141 42585 17175 42619
rect 22017 42585 22051 42619
rect 22753 42585 22787 42619
rect 22937 42585 22971 42619
rect 34161 42585 34195 42619
rect 38761 42585 38795 42619
rect 1501 42517 1535 42551
rect 9597 42517 9631 42551
rect 11161 42517 11195 42551
rect 11805 42517 11839 42551
rect 14381 42517 14415 42551
rect 15393 42517 15427 42551
rect 18613 42517 18647 42551
rect 20821 42517 20855 42551
rect 22569 42517 22603 42551
rect 24409 42517 24443 42551
rect 25421 42517 25455 42551
rect 25605 42517 25639 42551
rect 26157 42517 26191 42551
rect 26709 42517 26743 42551
rect 28733 42517 28767 42551
rect 31125 42517 31159 42551
rect 31769 42517 31803 42551
rect 33793 42517 33827 42551
rect 33961 42517 33995 42551
rect 36001 42517 36035 42551
rect 36185 42517 36219 42551
rect 36553 42517 36587 42551
rect 38301 42517 38335 42551
rect 39957 42517 39991 42551
rect 47961 42517 47995 42551
rect 11713 42313 11747 42347
rect 12357 42313 12391 42347
rect 13185 42313 13219 42347
rect 14105 42313 14139 42347
rect 15209 42313 15243 42347
rect 17325 42313 17359 42347
rect 20545 42313 20579 42347
rect 21189 42313 21223 42347
rect 21833 42313 21867 42347
rect 24041 42313 24075 42347
rect 24869 42313 24903 42347
rect 35357 42313 35391 42347
rect 35449 42313 35483 42347
rect 36001 42313 36035 42347
rect 14565 42245 14599 42279
rect 34069 42245 34103 42279
rect 12817 42177 12851 42211
rect 13001 42177 13035 42211
rect 15669 42177 15703 42211
rect 16037 42177 16071 42211
rect 16681 42177 16715 42211
rect 16865 42177 16899 42211
rect 17969 42177 18003 42211
rect 18613 42177 18647 42211
rect 21097 42177 21131 42211
rect 21281 42177 21315 42211
rect 22017 42177 22051 42211
rect 22293 42177 22327 42211
rect 22477 42177 22511 42211
rect 22937 42177 22971 42211
rect 23121 42177 23155 42211
rect 23765 42177 23799 42211
rect 23857 42177 23891 42211
rect 24501 42177 24535 42211
rect 24593 42177 24627 42211
rect 25513 42177 25547 42211
rect 28293 42177 28327 42211
rect 28549 42177 28583 42211
rect 29009 42177 29043 42211
rect 32393 42177 32427 42211
rect 35081 42177 35115 42211
rect 35541 42177 35575 42211
rect 36185 42177 36219 42211
rect 37473 42177 37507 42211
rect 37749 42177 37783 42211
rect 38301 42177 38335 42211
rect 38485 42177 38519 42211
rect 38577 42177 38611 42211
rect 39037 42177 39071 42211
rect 39221 42177 39255 42211
rect 15945 42109 15979 42143
rect 18521 42109 18555 42143
rect 22109 42109 22143 42143
rect 24041 42109 24075 42143
rect 29285 42109 29319 42143
rect 31125 42109 31159 42143
rect 32137 42109 32171 42143
rect 36369 42109 36403 42143
rect 37565 42109 37599 42143
rect 16129 42041 16163 42075
rect 18981 42041 19015 42075
rect 19993 42041 20027 42075
rect 22201 42041 22235 42075
rect 23029 42041 23063 42075
rect 37657 42041 37691 42075
rect 38301 42041 38335 42075
rect 10425 41973 10459 42007
rect 10885 41973 10919 42007
rect 15761 41973 15795 42007
rect 16773 41973 16807 42007
rect 19533 41973 19567 42007
rect 24685 41973 24719 42007
rect 25421 41973 25455 42007
rect 26065 41973 26099 42007
rect 27169 41973 27203 42007
rect 30389 41973 30423 42007
rect 33517 41973 33551 42007
rect 37289 41973 37323 42007
rect 39129 41973 39163 42007
rect 39773 41973 39807 42007
rect 40233 41973 40267 42007
rect 40785 41973 40819 42007
rect 12449 41769 12483 41803
rect 14197 41769 14231 41803
rect 15577 41769 15611 41803
rect 17417 41769 17451 41803
rect 18429 41769 18463 41803
rect 19809 41769 19843 41803
rect 20729 41769 20763 41803
rect 22017 41769 22051 41803
rect 23857 41769 23891 41803
rect 26525 41769 26559 41803
rect 28273 41769 28307 41803
rect 32597 41769 32631 41803
rect 35449 41769 35483 41803
rect 36369 41769 36403 41803
rect 38301 41769 38335 41803
rect 38485 41769 38519 41803
rect 15025 41701 15059 41735
rect 22753 41701 22787 41735
rect 25513 41701 25547 41735
rect 34805 41701 34839 41735
rect 39865 41701 39899 41735
rect 19349 41633 19383 41667
rect 24501 41633 24535 41667
rect 29561 41633 29595 41667
rect 31217 41633 31251 41667
rect 33977 41633 34011 41667
rect 37749 41633 37783 41667
rect 39221 41633 39255 41667
rect 14752 41565 14786 41599
rect 15025 41565 15059 41599
rect 15485 41565 15519 41599
rect 15761 41565 15795 41599
rect 16773 41565 16807 41599
rect 16957 41565 16991 41599
rect 17049 41565 17083 41599
rect 17141 41565 17175 41599
rect 18337 41565 18371 41599
rect 18521 41565 18555 41599
rect 19441 41565 19475 41599
rect 19625 41565 19659 41599
rect 21833 41565 21867 41599
rect 22109 41565 22143 41599
rect 24409 41565 24443 41599
rect 24593 41565 24627 41599
rect 27813 41565 27847 41599
rect 29837 41565 29871 41599
rect 32413 41565 32447 41599
rect 32597 41565 32631 41599
rect 33609 41565 33643 41599
rect 34069 41565 34103 41599
rect 35817 41565 35851 41599
rect 36277 41565 36311 41599
rect 36461 41565 36495 41599
rect 37657 41565 37691 41599
rect 39129 41565 39163 41599
rect 39313 41565 39347 41599
rect 11805 41497 11839 41531
rect 21925 41497 21959 41531
rect 33701 41497 33735 41531
rect 35633 41497 35667 41531
rect 38469 41497 38503 41531
rect 38669 41497 38703 41531
rect 40969 41497 41003 41531
rect 11253 41429 11287 41463
rect 13001 41429 13035 41463
rect 13461 41429 13495 41463
rect 14841 41429 14875 41463
rect 15945 41429 15979 41463
rect 21281 41429 21315 41463
rect 23305 41429 23339 41463
rect 28917 41429 28951 41463
rect 31769 41429 31803 41463
rect 33333 41429 33367 41463
rect 33793 41429 33827 41463
rect 37289 41429 37323 41463
rect 40509 41429 40543 41463
rect 12541 41225 12575 41259
rect 13645 41225 13679 41259
rect 14197 41225 14231 41259
rect 15117 41225 15151 41259
rect 16129 41225 16163 41259
rect 17693 41225 17727 41259
rect 19809 41225 19843 41259
rect 20361 41225 20395 41259
rect 22753 41225 22787 41259
rect 23397 41225 23431 41259
rect 23949 41225 23983 41259
rect 26249 41225 26283 41259
rect 27813 41225 27847 41259
rect 29101 41225 29135 41259
rect 34345 41225 34379 41259
rect 36553 41225 36587 41259
rect 38669 41225 38703 41259
rect 40785 41225 40819 41259
rect 14933 41157 14967 41191
rect 18705 41157 18739 41191
rect 19441 41157 19475 41191
rect 21281 41157 21315 41191
rect 26985 41157 27019 41191
rect 30389 41157 30423 41191
rect 32382 41157 32416 41191
rect 38485 41157 38519 41191
rect 14105 41089 14139 41123
rect 14289 41089 14323 41123
rect 14749 41089 14783 41123
rect 15761 41089 15795 41123
rect 15853 41089 15887 41123
rect 15945 41089 15979 41123
rect 16865 41089 16899 41123
rect 17693 41089 17727 41123
rect 17877 41089 17911 41123
rect 18429 41089 18463 41123
rect 18521 41089 18555 41123
rect 19165 41089 19199 41123
rect 19258 41089 19292 41123
rect 19533 41089 19567 41123
rect 19649 41089 19683 41123
rect 20269 41089 20303 41123
rect 20453 41089 20487 41123
rect 21833 41089 21867 41123
rect 22017 41089 22051 41123
rect 22201 41089 22235 41123
rect 22661 41089 22695 41123
rect 22845 41089 22879 41123
rect 24409 41089 24443 41123
rect 24501 41089 24535 41123
rect 24685 41089 24719 41123
rect 25421 41089 25455 41123
rect 32137 41089 32171 41123
rect 34069 41089 34103 41123
rect 34805 41089 34839 41123
rect 34989 41089 35023 41123
rect 35725 41089 35759 41123
rect 36461 41089 36495 41123
rect 36645 41089 36679 41123
rect 38301 41089 38335 41123
rect 11989 41021 12023 41055
rect 15669 41021 15703 41055
rect 16773 41021 16807 41055
rect 25697 41021 25731 41055
rect 34345 41021 34379 41055
rect 36001 41021 36035 41055
rect 40233 41021 40267 41055
rect 17233 40953 17267 40987
rect 24685 40953 24719 40987
rect 25605 40953 25639 40987
rect 39221 40953 39255 40987
rect 10977 40885 11011 40919
rect 13001 40885 13035 40919
rect 18705 40885 18739 40919
rect 25513 40885 25547 40919
rect 30849 40885 30883 40919
rect 31401 40885 31435 40919
rect 33517 40885 33551 40919
rect 34161 40885 34195 40919
rect 34897 40885 34931 40919
rect 35817 40885 35851 40919
rect 35909 40885 35943 40919
rect 37289 40885 37323 40919
rect 39681 40885 39715 40919
rect 41429 40885 41463 40919
rect 12449 40681 12483 40715
rect 12909 40681 12943 40715
rect 13553 40681 13587 40715
rect 15853 40681 15887 40715
rect 16497 40681 16531 40715
rect 18705 40681 18739 40715
rect 19809 40681 19843 40715
rect 20453 40681 20487 40715
rect 22293 40681 22327 40715
rect 25145 40681 25179 40715
rect 25789 40681 25823 40715
rect 25973 40681 26007 40715
rect 28917 40681 28951 40715
rect 32413 40681 32447 40715
rect 32597 40681 32631 40715
rect 34161 40681 34195 40715
rect 37749 40681 37783 40715
rect 40417 40681 40451 40715
rect 15209 40613 15243 40647
rect 20269 40613 20303 40647
rect 22845 40613 22879 40647
rect 23857 40613 23891 40647
rect 26709 40613 26743 40647
rect 30941 40613 30975 40647
rect 19257 40545 19291 40579
rect 22017 40545 22051 40579
rect 22753 40545 22787 40579
rect 27537 40545 27571 40579
rect 29561 40545 29595 40579
rect 33425 40545 33459 40579
rect 36369 40545 36403 40579
rect 38669 40545 38703 40579
rect 39865 40545 39899 40579
rect 11897 40477 11931 40511
rect 15025 40477 15059 40511
rect 15761 40477 15795 40511
rect 17601 40477 17635 40511
rect 18050 40477 18084 40511
rect 18154 40477 18188 40511
rect 18526 40477 18560 40511
rect 19533 40477 19567 40511
rect 19625 40477 19659 40511
rect 21097 40477 21131 40511
rect 21281 40477 21315 40511
rect 21925 40477 21959 40511
rect 22937 40477 22971 40511
rect 23029 40477 23063 40511
rect 23581 40477 23615 40511
rect 23857 40477 23891 40511
rect 24501 40477 24535 40511
rect 24594 40477 24628 40511
rect 25005 40477 25039 40511
rect 26433 40477 26467 40511
rect 26709 40477 26743 40511
rect 27804 40477 27838 40511
rect 31769 40477 31803 40511
rect 33241 40477 33275 40511
rect 33885 40477 33919 40511
rect 34713 40477 34747 40511
rect 34897 40477 34931 40511
rect 35541 40477 35575 40511
rect 35633 40477 35667 40511
rect 36277 40477 36311 40511
rect 36461 40477 36495 40511
rect 37933 40477 37967 40511
rect 38025 40477 38059 40511
rect 47869 40477 47903 40511
rect 1869 40409 1903 40443
rect 2053 40409 2087 40443
rect 18337 40409 18371 40443
rect 18429 40409 18463 40443
rect 20637 40409 20671 40443
rect 21189 40409 21223 40443
rect 24777 40409 24811 40443
rect 24869 40409 24903 40443
rect 25605 40409 25639 40443
rect 26525 40409 26559 40443
rect 29828 40409 29862 40443
rect 32229 40409 32263 40443
rect 32429 40409 32463 40443
rect 33057 40409 33091 40443
rect 34161 40409 34195 40443
rect 35817 40409 35851 40443
rect 36921 40409 36955 40443
rect 37105 40409 37139 40443
rect 47317 40409 47351 40443
rect 14473 40341 14507 40375
rect 17049 40341 17083 40375
rect 19441 40341 19475 40375
rect 20427 40341 20461 40375
rect 23673 40341 23707 40375
rect 25805 40341 25839 40375
rect 31585 40341 31619 40375
rect 33977 40341 34011 40375
rect 35081 40341 35115 40375
rect 35718 40341 35752 40375
rect 37289 40341 37323 40375
rect 39129 40341 39163 40375
rect 41061 40341 41095 40375
rect 41521 40341 41555 40375
rect 42073 40341 42107 40375
rect 48053 40341 48087 40375
rect 1593 40137 1627 40171
rect 13829 40137 13863 40171
rect 15485 40137 15519 40171
rect 23121 40137 23155 40171
rect 23489 40137 23523 40171
rect 24501 40137 24535 40171
rect 25513 40137 25547 40171
rect 27162 40137 27196 40171
rect 35541 40137 35575 40171
rect 36645 40137 36679 40171
rect 38754 40137 38788 40171
rect 41613 40137 41647 40171
rect 13277 40069 13311 40103
rect 19165 40069 19199 40103
rect 19349 40069 19383 40103
rect 20545 40069 20579 40103
rect 32597 40069 32631 40103
rect 38669 40069 38703 40103
rect 12081 40001 12115 40035
rect 12633 40001 12667 40035
rect 14473 40001 14507 40035
rect 17325 40001 17359 40035
rect 20269 40001 20303 40035
rect 20361 40001 20395 40035
rect 21005 40001 21039 40035
rect 21189 40001 21223 40035
rect 21990 40001 22024 40035
rect 23029 40001 23063 40035
rect 23305 40001 23339 40035
rect 24133 40001 24167 40035
rect 25881 40001 25915 40035
rect 26985 40001 27019 40035
rect 27077 40001 27111 40035
rect 27261 40001 27295 40035
rect 27721 40001 27755 40035
rect 27905 40001 27939 40035
rect 29193 40001 29227 40035
rect 29377 40001 29411 40035
rect 30113 40001 30147 40035
rect 30297 40001 30331 40035
rect 30849 40001 30883 40035
rect 33425 40001 33459 40035
rect 33609 40001 33643 40035
rect 34253 40001 34287 40035
rect 34621 40001 34655 40035
rect 34805 40001 34839 40035
rect 35725 40001 35759 40035
rect 36001 40001 36035 40035
rect 36553 40001 36587 40035
rect 36737 40001 36771 40035
rect 37473 40001 37507 40035
rect 37749 40001 37783 40035
rect 38577 40001 38611 40035
rect 38853 40001 38887 40035
rect 39313 40001 39347 40035
rect 39497 40001 39531 40035
rect 40509 40001 40543 40035
rect 14381 39933 14415 39967
rect 14841 39933 14875 39967
rect 17233 39933 17267 39967
rect 18981 39933 19015 39967
rect 22109 39933 22143 39967
rect 24041 39933 24075 39967
rect 25789 39933 25823 39967
rect 27813 39933 27847 39967
rect 34069 39933 34103 39967
rect 34437 39933 34471 39967
rect 34529 39933 34563 39967
rect 35817 39933 35851 39967
rect 37289 39933 37323 39967
rect 37565 39933 37599 39967
rect 17693 39865 17727 39899
rect 20545 39865 20579 39899
rect 22385 39865 22419 39899
rect 29377 39865 29411 39899
rect 33425 39865 33459 39899
rect 35909 39865 35943 39899
rect 37657 39865 37691 39899
rect 40049 39865 40083 39899
rect 16129 39797 16163 39831
rect 18429 39797 18463 39831
rect 21189 39797 21223 39831
rect 24961 39797 24995 39831
rect 25881 39797 25915 39831
rect 26433 39797 26467 39831
rect 28365 39797 28399 39831
rect 30205 39797 30239 39831
rect 31309 39797 31343 39831
rect 32873 39797 32907 39831
rect 39405 39797 39439 39831
rect 41061 39797 41095 39831
rect 42441 39797 42475 39831
rect 43085 39797 43119 39831
rect 11161 39593 11195 39627
rect 12817 39593 12851 39627
rect 20913 39593 20947 39627
rect 22293 39593 22327 39627
rect 23857 39593 23891 39627
rect 26709 39593 26743 39627
rect 28641 39593 28675 39627
rect 33333 39593 33367 39627
rect 36277 39593 36311 39627
rect 38761 39593 38795 39627
rect 38945 39593 38979 39627
rect 39957 39593 39991 39627
rect 15577 39525 15611 39559
rect 17877 39525 17911 39559
rect 27261 39525 27295 39559
rect 27997 39525 28031 39559
rect 33793 39525 33827 39559
rect 15117 39457 15151 39491
rect 20545 39457 20579 39491
rect 21833 39457 21867 39491
rect 21925 39457 21959 39491
rect 25789 39457 25823 39491
rect 29653 39457 29687 39491
rect 30113 39457 30147 39491
rect 32873 39457 32907 39491
rect 34713 39457 34747 39491
rect 37105 39457 37139 39491
rect 42165 39457 42199 39491
rect 43821 39457 43855 39491
rect 13369 39389 13403 39423
rect 13553 39389 13587 39423
rect 14105 39389 14139 39423
rect 15209 39389 15243 39423
rect 16221 39389 16255 39423
rect 16405 39389 16439 39423
rect 17785 39389 17819 39423
rect 18061 39389 18095 39423
rect 18153 39389 18187 39423
rect 20453 39389 20487 39423
rect 20637 39389 20671 39423
rect 20729 39389 20763 39423
rect 22109 39389 22143 39423
rect 22937 39389 22971 39423
rect 23489 39389 23523 39423
rect 24777 39389 24811 39423
rect 25513 39389 25547 39423
rect 25605 39389 25639 39423
rect 26249 39389 26283 39423
rect 26525 39389 26559 39423
rect 27445 39389 27479 39423
rect 27997 39389 28031 39423
rect 28181 39389 28215 39423
rect 28641 39389 28675 39423
rect 28825 39389 28859 39423
rect 29745 39389 29779 39423
rect 29929 39389 29963 39423
rect 31401 39389 31435 39423
rect 31585 39389 31619 39423
rect 32965 39389 32999 39423
rect 33977 39389 34011 39423
rect 34161 39389 34195 39423
rect 34871 39389 34905 39423
rect 35081 39389 35115 39423
rect 35173 39389 35207 39423
rect 36461 39389 36495 39423
rect 36553 39389 36587 39423
rect 38117 39389 38151 39423
rect 38301 39389 38335 39423
rect 39865 39389 39899 39423
rect 40049 39389 40083 39423
rect 41153 39389 41187 39423
rect 43269 39389 43303 39423
rect 11713 39321 11747 39355
rect 14289 39321 14323 39355
rect 14473 39321 14507 39355
rect 18337 39321 18371 39355
rect 23673 39321 23707 39355
rect 25789 39321 25823 39355
rect 34989 39321 35023 39355
rect 39129 39321 39163 39355
rect 41613 39321 41647 39355
rect 12265 39253 12299 39287
rect 13461 39253 13495 39287
rect 16221 39253 16255 39287
rect 17233 39253 17267 39287
rect 19349 39253 19383 39287
rect 19809 39253 19843 39287
rect 24961 39253 24995 39287
rect 26341 39253 26375 39287
rect 30849 39253 30883 39287
rect 35357 39253 35391 39287
rect 38301 39253 38335 39287
rect 38929 39253 38963 39287
rect 40601 39253 40635 39287
rect 42717 39253 42751 39287
rect 11805 39049 11839 39083
rect 13461 39049 13495 39083
rect 14289 39049 14323 39083
rect 15301 39049 15335 39083
rect 16129 39049 16163 39083
rect 18521 39049 18555 39083
rect 21097 39049 21131 39083
rect 21925 39049 21959 39083
rect 23581 39049 23615 39083
rect 28365 39049 28399 39083
rect 30389 39049 30423 39083
rect 31125 39049 31159 39083
rect 37565 39049 37599 39083
rect 38209 39049 38243 39083
rect 38377 39049 38411 39083
rect 39037 39049 39071 39083
rect 39865 39049 39899 39083
rect 43545 39049 43579 39083
rect 15945 38981 15979 39015
rect 18429 38981 18463 39015
rect 20453 38981 20487 39015
rect 22753 38981 22787 39015
rect 22937 38981 22971 39015
rect 24653 38981 24687 39015
rect 24869 38981 24903 39015
rect 25513 38981 25547 39015
rect 31033 38981 31067 39015
rect 32597 38981 32631 39015
rect 33517 38981 33551 39015
rect 33885 38981 33919 39015
rect 37749 38981 37783 39015
rect 38577 38981 38611 39015
rect 39221 38981 39255 39015
rect 40049 38981 40083 39015
rect 13369 38913 13403 38947
rect 13553 38913 13587 38947
rect 14473 38913 14507 38947
rect 14565 38913 14599 38947
rect 15117 38913 15151 38947
rect 15301 38913 15335 38947
rect 15761 38913 15795 38947
rect 16865 38913 16899 38947
rect 19441 38913 19475 38947
rect 20085 38913 20119 38947
rect 20269 38913 20303 38947
rect 20913 38913 20947 38947
rect 21097 38913 21131 38947
rect 21833 38913 21867 38947
rect 22201 38913 22235 38947
rect 23029 38913 23063 38947
rect 23765 38913 23799 38947
rect 23857 38913 23891 38947
rect 25329 38913 25363 38947
rect 25605 38913 25639 38947
rect 28549 38913 28583 38947
rect 28641 38913 28675 38947
rect 28917 38913 28951 38947
rect 29745 38913 29779 38947
rect 32965 38913 32999 38947
rect 34345 38913 34379 38947
rect 34529 38913 34563 38947
rect 34621 38913 34655 38947
rect 36185 38913 36219 38947
rect 36369 38913 36403 38947
rect 37473 38913 37507 38947
rect 39405 38913 39439 38947
rect 40233 38913 40267 38947
rect 12909 38845 12943 38879
rect 14289 38845 14323 38879
rect 16681 38845 16715 38879
rect 19257 38845 19291 38879
rect 22017 38845 22051 38879
rect 23581 38845 23615 38879
rect 29653 38845 29687 38879
rect 41797 38845 41831 38879
rect 17877 38777 17911 38811
rect 22201 38777 22235 38811
rect 25329 38777 25363 38811
rect 27445 38777 27479 38811
rect 41245 38777 41279 38811
rect 10885 38709 10919 38743
rect 12265 38709 12299 38743
rect 17049 38709 17083 38743
rect 19625 38709 19659 38743
rect 22753 38709 22787 38743
rect 24501 38709 24535 38743
rect 24685 38709 24719 38743
rect 26341 38709 26375 38743
rect 28825 38709 28859 38743
rect 29377 38709 29411 38743
rect 34345 38709 34379 38743
rect 35173 38709 35207 38743
rect 35725 38709 35759 38743
rect 36277 38709 36311 38743
rect 37749 38709 37783 38743
rect 38393 38709 38427 38743
rect 40693 38709 40727 38743
rect 42533 38709 42567 38743
rect 42993 38709 43027 38743
rect 11253 38505 11287 38539
rect 14197 38505 14231 38539
rect 14749 38505 14783 38539
rect 15945 38505 15979 38539
rect 16681 38505 16715 38539
rect 17693 38505 17727 38539
rect 19901 38505 19935 38539
rect 20545 38505 20579 38539
rect 22017 38505 22051 38539
rect 22247 38505 22281 38539
rect 23121 38505 23155 38539
rect 23857 38505 23891 38539
rect 25145 38505 25179 38539
rect 27997 38505 28031 38539
rect 28917 38505 28951 38539
rect 32505 38505 32539 38539
rect 34713 38505 34747 38539
rect 40417 38505 40451 38539
rect 42625 38505 42659 38539
rect 13553 38437 13587 38471
rect 18613 38437 18647 38471
rect 21373 38437 21407 38471
rect 22109 38437 22143 38471
rect 23305 38437 23339 38471
rect 28825 38437 28859 38471
rect 29837 38437 29871 38471
rect 33793 38437 33827 38471
rect 37749 38437 37783 38471
rect 38853 38437 38887 38471
rect 42165 38437 42199 38471
rect 15761 38369 15795 38403
rect 16589 38369 16623 38403
rect 24685 38369 24719 38403
rect 25697 38369 25731 38403
rect 26525 38369 26559 38403
rect 27537 38369 27571 38403
rect 29009 38369 29043 38403
rect 31309 38369 31343 38403
rect 32965 38369 32999 38403
rect 34897 38369 34931 38403
rect 35081 38369 35115 38403
rect 35173 38369 35207 38403
rect 36001 38369 36035 38403
rect 37197 38369 37231 38403
rect 38025 38369 38059 38403
rect 2053 38301 2087 38335
rect 14933 38301 14967 38335
rect 15209 38301 15243 38335
rect 15945 38301 15979 38335
rect 16865 38301 16899 38335
rect 17601 38301 17635 38335
rect 17785 38301 17819 38335
rect 18429 38301 18463 38335
rect 19809 38301 19843 38335
rect 19993 38301 20027 38335
rect 20453 38301 20487 38335
rect 20637 38301 20671 38335
rect 21925 38301 21959 38335
rect 22385 38301 22419 38335
rect 24409 38301 24443 38335
rect 24593 38301 24627 38335
rect 24777 38301 24811 38335
rect 24961 38301 24995 38335
rect 26433 38301 26467 38335
rect 27261 38301 27295 38335
rect 27445 38301 27479 38335
rect 27629 38301 27663 38335
rect 27813 38301 27847 38335
rect 28733 38301 28767 38335
rect 29653 38301 29687 38335
rect 29745 38301 29779 38335
rect 29929 38301 29963 38335
rect 31217 38301 31251 38335
rect 32689 38301 32723 38335
rect 32781 38301 32815 38335
rect 33057 38301 33091 38335
rect 33517 38301 33551 38335
rect 33609 38301 33643 38335
rect 34989 38301 35023 38335
rect 36093 38301 36127 38335
rect 37105 38301 37139 38335
rect 37933 38301 37967 38335
rect 38117 38301 38151 38335
rect 38209 38301 38243 38335
rect 38761 38301 38795 38335
rect 38945 38301 38979 38335
rect 41613 38301 41647 38335
rect 47409 38301 47443 38335
rect 47869 38301 47903 38335
rect 1869 38233 1903 38267
rect 11897 38233 11931 38267
rect 13001 38233 13035 38267
rect 15669 38233 15703 38267
rect 18245 38233 18279 38267
rect 22937 38233 22971 38267
rect 33793 38233 33827 38267
rect 40969 38233 41003 38267
rect 12449 38165 12483 38199
rect 15117 38165 15151 38199
rect 16129 38165 16163 38199
rect 17049 38165 17083 38199
rect 19349 38165 19383 38199
rect 23137 38165 23171 38199
rect 26801 38165 26835 38199
rect 30113 38165 30147 38199
rect 31585 38165 31619 38199
rect 35725 38165 35759 38199
rect 36737 38165 36771 38199
rect 39865 38165 39899 38199
rect 43177 38165 43211 38199
rect 48053 38165 48087 38199
rect 1593 37961 1627 37995
rect 12357 37961 12391 37995
rect 16858 37961 16892 37995
rect 18705 37961 18739 37995
rect 22017 37961 22051 37995
rect 23397 37961 23431 37995
rect 23489 37961 23523 37995
rect 24869 37961 24903 37995
rect 25421 37961 25455 37995
rect 26433 37961 26467 37995
rect 30113 37961 30147 37995
rect 34897 37961 34931 37995
rect 36001 37961 36035 37995
rect 38209 37961 38243 37995
rect 41153 37961 41187 37995
rect 41705 37961 41739 37995
rect 42533 37961 42567 37995
rect 13461 37893 13495 37927
rect 14565 37893 14599 37927
rect 16773 37893 16807 37927
rect 27169 37893 27203 37927
rect 28181 37893 28215 37927
rect 28273 37893 28307 37927
rect 31033 37893 31067 37927
rect 35081 37893 35115 37927
rect 37381 37893 37415 37927
rect 13921 37825 13955 37859
rect 14105 37825 14139 37859
rect 14197 37825 14231 37859
rect 14289 37825 14323 37859
rect 15209 37825 15243 37859
rect 15485 37825 15519 37859
rect 16681 37825 16715 37859
rect 16957 37825 16991 37859
rect 17877 37825 17911 37859
rect 18981 37825 19015 37859
rect 20361 37825 20395 37859
rect 22109 37825 22143 37859
rect 22293 37825 22327 37859
rect 23581 37825 23615 37859
rect 24225 37825 24259 37859
rect 24501 37825 24535 37859
rect 24685 37825 24719 37859
rect 25973 37825 26007 37859
rect 26249 37825 26283 37859
rect 27537 37825 27571 37859
rect 27997 37825 28031 37859
rect 28365 37825 28399 37859
rect 29377 37825 29411 37859
rect 30297 37825 30331 37859
rect 30481 37825 30515 37859
rect 30941 37825 30975 37859
rect 31125 37825 31159 37859
rect 32413 37825 32447 37859
rect 32505 37825 32539 37859
rect 32597 37825 32631 37859
rect 32781 37825 32815 37859
rect 33609 37825 33643 37859
rect 33793 37825 33827 37859
rect 35265 37825 35299 37859
rect 36185 37825 36219 37859
rect 36461 37825 36495 37859
rect 37289 37825 37323 37859
rect 37473 37825 37507 37859
rect 38577 37825 38611 37859
rect 40509 37825 40543 37859
rect 15301 37757 15335 37791
rect 17785 37757 17819 37791
rect 18705 37757 18739 37791
rect 23765 37757 23799 37791
rect 24409 37757 24443 37791
rect 24593 37757 24627 37791
rect 26065 37757 26099 37791
rect 32137 37757 32171 37791
rect 38485 37757 38519 37791
rect 40601 37757 40635 37791
rect 12817 37689 12851 37723
rect 15025 37689 15059 37723
rect 18245 37689 18279 37723
rect 23213 37689 23247 37723
rect 26157 37689 26191 37723
rect 26985 37689 27019 37723
rect 28549 37689 28583 37723
rect 29561 37689 29595 37723
rect 36369 37689 36403 37723
rect 39221 37689 39255 37723
rect 10885 37621 10919 37655
rect 11713 37621 11747 37655
rect 15485 37621 15519 37655
rect 16037 37621 16071 37655
rect 18889 37621 18923 37655
rect 19901 37621 19935 37655
rect 20637 37621 20671 37655
rect 20821 37621 20855 37655
rect 21833 37621 21867 37655
rect 27169 37621 27203 37655
rect 33609 37621 33643 37655
rect 33977 37621 34011 37655
rect 40141 37621 40175 37655
rect 11529 37417 11563 37451
rect 14381 37417 14415 37451
rect 16037 37417 16071 37451
rect 18613 37417 18647 37451
rect 19625 37417 19659 37451
rect 20913 37417 20947 37451
rect 24961 37417 24995 37451
rect 25697 37417 25731 37451
rect 26249 37417 26283 37451
rect 27445 37417 27479 37451
rect 27997 37417 28031 37451
rect 32137 37417 32171 37451
rect 32873 37417 32907 37451
rect 35817 37417 35851 37451
rect 38485 37417 38519 37451
rect 41153 37417 41187 37451
rect 41705 37417 41739 37451
rect 42809 37417 42843 37451
rect 43361 37417 43395 37451
rect 10977 37349 11011 37383
rect 21649 37349 21683 37383
rect 31309 37349 31343 37383
rect 37381 37349 37415 37383
rect 37841 37349 37875 37383
rect 42165 37349 42199 37383
rect 10333 37281 10367 37315
rect 18061 37281 18095 37315
rect 19533 37281 19567 37315
rect 21557 37281 21591 37315
rect 23213 37281 23247 37315
rect 24501 37281 24535 37315
rect 27077 37281 27111 37315
rect 27169 37281 27203 37315
rect 27261 37281 27295 37315
rect 39221 37281 39255 37315
rect 40969 37281 41003 37315
rect 12541 37213 12575 37247
rect 12725 37213 12759 37247
rect 13369 37213 13403 37247
rect 14197 37213 14231 37247
rect 14381 37213 14415 37247
rect 14841 37213 14875 37247
rect 15025 37213 15059 37247
rect 15209 37213 15243 37247
rect 15853 37213 15887 37247
rect 17325 37213 17359 37247
rect 17509 37213 17543 37247
rect 19441 37213 19475 37247
rect 20269 37213 20303 37247
rect 20453 37213 20487 37247
rect 20564 37207 20598 37241
rect 20683 37213 20717 37247
rect 21465 37213 21499 37247
rect 21741 37213 21775 37247
rect 23029 37213 23063 37247
rect 23673 37213 23707 37247
rect 23857 37213 23891 37247
rect 24409 37213 24443 37247
rect 24685 37213 24719 37247
rect 24777 37213 24811 37247
rect 26985 37213 27019 37247
rect 28457 37213 28491 37247
rect 28641 37213 28675 37247
rect 30205 37213 30239 37247
rect 30294 37213 30328 37247
rect 30389 37213 30423 37247
rect 30573 37213 30607 37247
rect 31217 37213 31251 37247
rect 31401 37213 31435 37247
rect 32045 37213 32079 37247
rect 32229 37213 32263 37247
rect 33517 37213 33551 37247
rect 33701 37213 33735 37247
rect 33793 37213 33827 37247
rect 33885 37213 33919 37247
rect 34713 37213 34747 37247
rect 36461 37213 36495 37247
rect 36829 37213 36863 37247
rect 39129 37213 39163 37247
rect 39313 37213 39347 37247
rect 39865 37213 39899 37247
rect 40049 37213 40083 37247
rect 40877 37213 40911 37247
rect 13185 37145 13219 37179
rect 15669 37145 15703 37179
rect 23765 37145 23799 37179
rect 32689 37145 32723 37179
rect 32889 37145 32923 37179
rect 34161 37145 34195 37179
rect 36001 37145 36035 37179
rect 36645 37145 36679 37179
rect 12081 37077 12115 37111
rect 12725 37077 12759 37111
rect 13553 37077 13587 37111
rect 16865 37077 16899 37111
rect 17509 37077 17543 37111
rect 19809 37077 19843 37111
rect 21925 37077 21959 37111
rect 22845 37077 22879 37111
rect 28549 37077 28583 37111
rect 29929 37077 29963 37111
rect 33057 37077 33091 37111
rect 34805 37077 34839 37111
rect 35633 37077 35667 37111
rect 35801 37077 35835 37111
rect 40049 37077 40083 37111
rect 40509 37077 40543 37111
rect 48053 37077 48087 37111
rect 10977 36873 11011 36907
rect 12449 36873 12483 36907
rect 13553 36873 13587 36907
rect 14289 36873 14323 36907
rect 19073 36873 19107 36907
rect 20729 36873 20763 36907
rect 22937 36873 22971 36907
rect 24409 36873 24443 36907
rect 26065 36873 26099 36907
rect 28273 36873 28307 36907
rect 33609 36873 33643 36907
rect 35725 36873 35759 36907
rect 40233 36873 40267 36907
rect 42533 36873 42567 36907
rect 43085 36873 43119 36907
rect 11897 36805 11931 36839
rect 15393 36805 15427 36839
rect 19809 36805 19843 36839
rect 23673 36805 23707 36839
rect 25145 36805 25179 36839
rect 25345 36805 25379 36839
rect 29837 36805 29871 36839
rect 32781 36805 32815 36839
rect 33761 36805 33795 36839
rect 33977 36805 34011 36839
rect 36093 36805 36127 36839
rect 38301 36805 38335 36839
rect 46673 36805 46707 36839
rect 47593 36805 47627 36839
rect 13461 36737 13495 36771
rect 13645 36737 13679 36771
rect 14105 36737 14139 36771
rect 14289 36737 14323 36771
rect 15117 36737 15151 36771
rect 15209 36737 15243 36771
rect 17417 36737 17451 36771
rect 17509 36737 17543 36771
rect 17693 36737 17727 36771
rect 18337 36737 18371 36771
rect 18521 36737 18555 36771
rect 18613 36737 18647 36771
rect 18889 36737 18923 36771
rect 19717 36737 19751 36771
rect 19901 36737 19935 36771
rect 20361 36737 20395 36771
rect 20545 36737 20579 36771
rect 22661 36737 22695 36771
rect 23397 36737 23431 36771
rect 24317 36737 24351 36771
rect 24501 36737 24535 36771
rect 27445 36737 27479 36771
rect 28457 36737 28491 36771
rect 28641 36737 28675 36771
rect 28733 36737 28767 36771
rect 28917 36737 28951 36771
rect 29561 36737 29595 36771
rect 29653 36737 29687 36771
rect 30389 36737 30423 36771
rect 30573 36737 30607 36771
rect 31217 36737 31251 36771
rect 31309 36737 31343 36771
rect 32505 36737 32539 36771
rect 32653 36737 32687 36771
rect 32870 36737 32904 36771
rect 32970 36737 33004 36771
rect 34529 36737 34563 36771
rect 34805 36737 34839 36771
rect 35817 36737 35851 36771
rect 35909 36737 35943 36771
rect 36553 36737 36587 36771
rect 36737 36737 36771 36771
rect 37933 36737 37967 36771
rect 38393 36737 38427 36771
rect 39129 36737 39163 36771
rect 39313 36737 39347 36771
rect 39773 36737 39807 36771
rect 41245 36737 41279 36771
rect 41429 36737 41463 36771
rect 46857 36737 46891 36771
rect 47777 36737 47811 36771
rect 47961 36737 47995 36771
rect 18705 36669 18739 36703
rect 21189 36669 21223 36703
rect 22293 36669 22327 36703
rect 22385 36669 22419 36703
rect 22753 36669 22787 36703
rect 23489 36669 23523 36703
rect 23673 36669 23707 36703
rect 27353 36669 27387 36703
rect 36645 36669 36679 36703
rect 40785 36669 40819 36703
rect 47041 36669 47075 36703
rect 15393 36601 15427 36635
rect 25513 36601 25547 36635
rect 28549 36601 28583 36635
rect 29837 36601 29871 36635
rect 34529 36601 34563 36635
rect 37289 36601 37323 36635
rect 38071 36601 38105 36635
rect 39313 36601 39347 36635
rect 13001 36533 13035 36567
rect 16129 36533 16163 36567
rect 16957 36533 16991 36567
rect 17877 36533 17911 36567
rect 25329 36533 25363 36567
rect 27813 36533 27847 36567
rect 30573 36533 30607 36567
rect 31309 36533 31343 36567
rect 33149 36533 33183 36567
rect 33793 36533 33827 36567
rect 35541 36533 35575 36567
rect 38209 36533 38243 36567
rect 39865 36533 39899 36567
rect 11897 36329 11931 36363
rect 15945 36329 15979 36363
rect 18245 36329 18279 36363
rect 18613 36329 18647 36363
rect 19349 36329 19383 36363
rect 20545 36329 20579 36363
rect 26985 36329 27019 36363
rect 27537 36329 27571 36363
rect 28365 36329 28399 36363
rect 31861 36329 31895 36363
rect 32873 36329 32907 36363
rect 35265 36329 35299 36363
rect 35633 36329 35667 36363
rect 38209 36329 38243 36363
rect 41981 36329 42015 36363
rect 47225 36329 47259 36363
rect 2237 36261 2271 36295
rect 25329 36261 25363 36295
rect 28825 36261 28859 36295
rect 36093 36261 36127 36295
rect 38485 36261 38519 36295
rect 40141 36261 40175 36295
rect 42441 36261 42475 36295
rect 15577 36193 15611 36227
rect 16589 36193 16623 36227
rect 17233 36193 17267 36227
rect 18337 36193 18371 36227
rect 22845 36193 22879 36227
rect 34805 36193 34839 36227
rect 35541 36193 35575 36227
rect 1685 36125 1719 36159
rect 13001 36125 13035 36159
rect 15669 36125 15703 36159
rect 16497 36125 16531 36159
rect 16681 36125 16715 36159
rect 17601 36125 17635 36159
rect 17693 36125 17727 36159
rect 18245 36125 18279 36159
rect 19257 36125 19291 36159
rect 19441 36125 19475 36159
rect 20453 36125 20487 36159
rect 20637 36125 20671 36159
rect 22109 36125 22143 36159
rect 22753 36125 22787 36159
rect 25053 36125 25087 36159
rect 25789 36125 25823 36159
rect 25973 36125 26007 36159
rect 27721 36125 27755 36159
rect 27905 36125 27939 36159
rect 28549 36125 28583 36159
rect 28641 36125 28675 36159
rect 28917 36125 28951 36159
rect 30297 36125 30331 36159
rect 30573 36125 30607 36159
rect 31401 36125 31435 36159
rect 31953 36125 31987 36159
rect 33057 36125 33091 36159
rect 33701 36125 33735 36159
rect 33885 36125 33919 36159
rect 35633 36125 35667 36159
rect 36277 36125 36311 36159
rect 36369 36125 36403 36159
rect 37013 36125 37047 36159
rect 37197 36125 37231 36159
rect 38025 36125 38059 36159
rect 38209 36125 38243 36159
rect 38945 36125 38979 36159
rect 39129 36125 39163 36159
rect 40049 36125 40083 36159
rect 40233 36125 40267 36159
rect 40325 36125 40359 36159
rect 40509 36125 40543 36159
rect 41153 36125 41187 36159
rect 41245 36103 41279 36137
rect 41373 36125 41407 36159
rect 11345 36057 11379 36091
rect 12449 36057 12483 36091
rect 14473 36057 14507 36091
rect 19993 36057 20027 36091
rect 25329 36057 25363 36091
rect 26433 36057 26467 36091
rect 30757 36057 30791 36091
rect 33241 36057 33275 36091
rect 33793 36057 33827 36091
rect 36093 36057 36127 36091
rect 36829 36057 36863 36091
rect 40969 36057 41003 36091
rect 47869 36057 47903 36091
rect 48053 36057 48087 36091
rect 1501 35989 1535 36023
rect 13553 35989 13587 36023
rect 15025 35989 15059 36023
rect 17509 35989 17543 36023
rect 21465 35989 21499 36023
rect 23121 35989 23155 36023
rect 23765 35989 23799 36023
rect 24593 35989 24627 36023
rect 25145 35989 25179 36023
rect 25881 35989 25915 36023
rect 39037 35989 39071 36023
rect 39865 35989 39899 36023
rect 42993 35989 43027 36023
rect 10885 35785 10919 35819
rect 12173 35785 12207 35819
rect 12725 35785 12759 35819
rect 13277 35785 13311 35819
rect 15761 35785 15795 35819
rect 17049 35785 17083 35819
rect 20637 35785 20671 35819
rect 21005 35785 21039 35819
rect 24041 35785 24075 35819
rect 25145 35785 25179 35819
rect 31125 35785 31159 35819
rect 32413 35785 32447 35819
rect 33609 35785 33643 35819
rect 35541 35785 35575 35819
rect 36185 35785 36219 35819
rect 38485 35785 38519 35819
rect 48053 35785 48087 35819
rect 17877 35717 17911 35751
rect 28273 35717 28307 35751
rect 29193 35717 29227 35751
rect 34069 35717 34103 35751
rect 38117 35717 38151 35751
rect 38317 35717 38351 35751
rect 39221 35717 39255 35751
rect 14289 35649 14323 35683
rect 14473 35649 14507 35683
rect 15393 35649 15427 35683
rect 16681 35649 16715 35683
rect 16865 35649 16899 35683
rect 18153 35649 18187 35683
rect 18613 35649 18647 35683
rect 19073 35649 19107 35683
rect 19717 35649 19751 35683
rect 19901 35649 19935 35683
rect 20545 35649 20579 35683
rect 20821 35649 20855 35683
rect 22569 35649 22603 35683
rect 24501 35649 24535 35683
rect 24685 35649 24719 35683
rect 24777 35649 24811 35683
rect 24869 35649 24903 35683
rect 25789 35649 25823 35683
rect 25882 35649 25916 35683
rect 26157 35649 26191 35683
rect 26985 35649 27019 35683
rect 29377 35649 29411 35683
rect 30389 35649 30423 35683
rect 30573 35649 30607 35683
rect 30665 35649 30699 35683
rect 30941 35649 30975 35683
rect 32229 35649 32263 35683
rect 32413 35649 32447 35683
rect 33425 35649 33459 35683
rect 34345 35649 34379 35683
rect 35449 35649 35483 35683
rect 35633 35649 35667 35683
rect 36277 35649 36311 35683
rect 37289 35649 37323 35683
rect 37473 35649 37507 35683
rect 38945 35649 38979 35683
rect 39037 35649 39071 35683
rect 40171 35649 40205 35683
rect 40325 35649 40359 35683
rect 15485 35581 15519 35615
rect 18797 35581 18831 35615
rect 18889 35581 18923 35615
rect 19257 35581 19291 35615
rect 25605 35581 25639 35615
rect 26065 35581 26099 35615
rect 27261 35581 27295 35615
rect 27813 35581 27847 35615
rect 29653 35581 29687 35615
rect 30757 35581 30791 35615
rect 33241 35581 33275 35615
rect 37381 35581 37415 35615
rect 18061 35513 18095 35547
rect 18153 35513 18187 35547
rect 18981 35513 19015 35547
rect 39221 35513 39255 35547
rect 10333 35445 10367 35479
rect 11621 35445 11655 35479
rect 13829 35445 13863 35479
rect 14473 35445 14507 35479
rect 19717 35445 19751 35479
rect 22477 35445 22511 35479
rect 23489 35445 23523 35479
rect 27077 35445 27111 35479
rect 27169 35445 27203 35479
rect 29561 35445 29595 35479
rect 34805 35445 34839 35479
rect 38301 35445 38335 35479
rect 40141 35445 40175 35479
rect 40877 35445 40911 35479
rect 41429 35445 41463 35479
rect 42441 35445 42475 35479
rect 43085 35445 43119 35479
rect 43545 35445 43579 35479
rect 10241 35241 10275 35275
rect 10793 35241 10827 35275
rect 11345 35241 11379 35275
rect 13553 35241 13587 35275
rect 15301 35241 15335 35275
rect 17785 35241 17819 35275
rect 18337 35241 18371 35275
rect 18705 35241 18739 35275
rect 19349 35241 19383 35275
rect 19993 35241 20027 35275
rect 21097 35241 21131 35275
rect 28089 35241 28123 35275
rect 30389 35241 30423 35275
rect 32505 35241 32539 35275
rect 33241 35241 33275 35275
rect 34897 35241 34931 35275
rect 39957 35241 39991 35275
rect 41521 35241 41555 35275
rect 42625 35241 42659 35275
rect 12817 35173 12851 35207
rect 24501 35173 24535 35207
rect 25329 35173 25363 35207
rect 29653 35173 29687 35207
rect 36553 35173 36587 35207
rect 15117 35105 15151 35139
rect 17417 35105 17451 35139
rect 18245 35105 18279 35139
rect 19901 35105 19935 35139
rect 20085 35105 20119 35139
rect 20821 35105 20855 35139
rect 21833 35105 21867 35139
rect 22753 35105 22787 35139
rect 23029 35105 23063 35139
rect 23857 35105 23891 35139
rect 25513 35105 25547 35139
rect 29005 35105 29039 35139
rect 33701 35105 33735 35139
rect 34713 35105 34747 35139
rect 36277 35105 36311 35139
rect 40141 35105 40175 35139
rect 11805 35037 11839 35071
rect 11989 35037 12023 35071
rect 12725 35037 12759 35071
rect 12817 35037 12851 35071
rect 13461 35037 13495 35071
rect 13553 35037 13587 35071
rect 14105 35037 14139 35071
rect 14381 35037 14415 35071
rect 15577 35037 15611 35071
rect 16221 35037 16255 35071
rect 16313 35037 16347 35071
rect 17601 35037 17635 35071
rect 18521 35037 18555 35071
rect 19809 35037 19843 35071
rect 20729 35037 20763 35071
rect 21557 35037 21591 35071
rect 21649 35037 21683 35071
rect 22385 35037 22419 35071
rect 22569 35037 22603 35071
rect 23121 35037 23155 35071
rect 24501 35037 24535 35071
rect 24685 35037 24719 35071
rect 25237 35037 25271 35071
rect 25973 35037 26007 35071
rect 26157 35037 26191 35071
rect 26341 35037 26375 35071
rect 26985 35037 27019 35071
rect 27261 35037 27295 35071
rect 28733 35037 28767 35071
rect 28825 35037 28859 35071
rect 30568 35037 30602 35071
rect 30940 35037 30974 35071
rect 31033 35037 31067 35071
rect 33425 35037 33459 35071
rect 33517 35037 33551 35071
rect 33793 35037 33827 35071
rect 34989 35037 35023 35071
rect 36185 35037 36219 35071
rect 37933 35037 37967 35071
rect 38117 35037 38151 35071
rect 38761 35037 38795 35071
rect 40233 35037 40267 35071
rect 40969 35037 41003 35071
rect 11897 34969 11931 35003
rect 12541 34969 12575 35003
rect 13277 34969 13311 35003
rect 14197 34969 14231 35003
rect 21833 34969 21867 35003
rect 27905 34969 27939 35003
rect 30665 34969 30699 35003
rect 30757 34969 30791 35003
rect 31493 34969 31527 35003
rect 31677 34969 31711 35003
rect 31861 34969 31895 35003
rect 32413 34969 32447 35003
rect 34713 34969 34747 35003
rect 38025 34969 38059 35003
rect 42073 34969 42107 35003
rect 14565 34901 14599 34935
rect 15485 34901 15519 34935
rect 16037 34901 16071 34935
rect 16957 34901 16991 34935
rect 25513 34901 25547 34935
rect 27077 34901 27111 34935
rect 27445 34901 27479 34935
rect 28105 34901 28139 34935
rect 28273 34901 28307 34935
rect 29009 34901 29043 34935
rect 35449 34901 35483 34935
rect 37013 34901 37047 34935
rect 38669 34901 38703 34935
rect 39313 34901 39347 34935
rect 43085 34901 43119 34935
rect 1961 34697 1995 34731
rect 9137 34697 9171 34731
rect 10241 34697 10275 34731
rect 10977 34697 11011 34731
rect 12541 34697 12575 34731
rect 12909 34697 12943 34731
rect 15577 34697 15611 34731
rect 15761 34697 15795 34731
rect 18077 34697 18111 34731
rect 18245 34697 18279 34731
rect 19717 34697 19751 34731
rect 21189 34697 21223 34731
rect 23121 34697 23155 34731
rect 24409 34697 24443 34731
rect 30389 34697 30423 34731
rect 31493 34697 31527 34731
rect 32229 34697 32263 34731
rect 33425 34697 33459 34731
rect 34161 34697 34195 34731
rect 36467 34697 36501 34731
rect 38209 34697 38243 34731
rect 38577 34697 38611 34731
rect 39221 34697 39255 34731
rect 39865 34697 39899 34731
rect 41429 34697 41463 34731
rect 11529 34629 11563 34663
rect 14933 34629 14967 34663
rect 17877 34629 17911 34663
rect 18797 34629 18831 34663
rect 23489 34629 23523 34663
rect 26341 34629 26375 34663
rect 32689 34629 32723 34663
rect 36553 34629 36587 34663
rect 37381 34629 37415 34663
rect 1869 34561 1903 34595
rect 10793 34561 10827 34595
rect 10977 34561 11011 34595
rect 11713 34561 11747 34595
rect 12449 34561 12483 34595
rect 12725 34561 12759 34595
rect 13829 34561 13863 34595
rect 13921 34561 13955 34595
rect 14105 34561 14139 34595
rect 14565 34561 14599 34595
rect 14749 34561 14783 34595
rect 15669 34561 15703 34595
rect 16865 34561 16899 34595
rect 19257 34561 19291 34595
rect 19349 34561 19383 34595
rect 19533 34561 19567 34595
rect 21005 34561 21039 34595
rect 22293 34561 22327 34595
rect 23259 34561 23293 34595
rect 23397 34561 23431 34595
rect 23672 34561 23706 34595
rect 23765 34561 23799 34595
rect 24225 34561 24259 34595
rect 24409 34561 24443 34595
rect 25053 34561 25087 34595
rect 25237 34561 25271 34595
rect 25329 34561 25363 34595
rect 25789 34561 25823 34595
rect 26065 34561 26099 34595
rect 26157 34561 26191 34595
rect 27169 34561 27203 34595
rect 27353 34561 27387 34595
rect 28641 34561 28675 34595
rect 28917 34561 28951 34595
rect 29101 34561 29135 34595
rect 29561 34561 29595 34595
rect 29745 34561 29779 34595
rect 29929 34561 29963 34595
rect 30757 34561 30791 34595
rect 31585 34561 31619 34595
rect 33333 34561 33367 34595
rect 33609 34561 33643 34595
rect 33701 34561 33735 34595
rect 34437 34561 34471 34595
rect 35541 34561 35575 34595
rect 36369 34561 36403 34595
rect 36645 34561 36679 34595
rect 37289 34561 37323 34595
rect 37565 34561 37599 34595
rect 38393 34561 38427 34595
rect 38669 34561 38703 34595
rect 39129 34561 39163 34595
rect 39313 34561 39347 34595
rect 40417 34561 40451 34595
rect 40601 34561 40635 34595
rect 15945 34493 15979 34527
rect 16773 34493 16807 34527
rect 20821 34493 20855 34527
rect 22201 34493 22235 34527
rect 25881 34493 25915 34527
rect 27077 34493 27111 34527
rect 27261 34493 27295 34527
rect 27537 34493 27571 34527
rect 28825 34493 28859 34527
rect 30849 34493 30883 34527
rect 33517 34493 33551 34527
rect 34161 34493 34195 34527
rect 35633 34493 35667 34527
rect 37749 34493 37783 34527
rect 42533 34493 42567 34527
rect 42993 34493 43027 34527
rect 15393 34425 15427 34459
rect 17233 34425 17267 34459
rect 22661 34425 22695 34459
rect 28733 34425 28767 34459
rect 35909 34425 35943 34459
rect 9781 34357 9815 34391
rect 11897 34357 11931 34391
rect 14105 34357 14139 34391
rect 18061 34357 18095 34391
rect 20361 34357 20395 34391
rect 25053 34357 25087 34391
rect 28457 34357 28491 34391
rect 34345 34357 34379 34391
rect 10333 34153 10367 34187
rect 14657 34153 14691 34187
rect 15393 34153 15427 34187
rect 16129 34153 16163 34187
rect 17969 34153 18003 34187
rect 21649 34153 21683 34187
rect 21833 34153 21867 34187
rect 25145 34153 25179 34187
rect 25329 34153 25363 34187
rect 25881 34153 25915 34187
rect 27629 34153 27663 34187
rect 28733 34153 28767 34187
rect 29837 34153 29871 34187
rect 31861 34153 31895 34187
rect 32413 34153 32447 34187
rect 33701 34153 33735 34187
rect 34713 34153 34747 34187
rect 35633 34153 35667 34187
rect 36461 34153 36495 34187
rect 39865 34153 39899 34187
rect 42073 34153 42107 34187
rect 1593 34085 1627 34119
rect 13553 34085 13587 34119
rect 16957 34085 16991 34119
rect 23213 34085 23247 34119
rect 27445 34085 27479 34119
rect 35725 34085 35759 34119
rect 37197 34085 37231 34119
rect 38853 34085 38887 34119
rect 42533 34085 42567 34119
rect 11529 34017 11563 34051
rect 11989 34017 12023 34051
rect 13277 34017 13311 34051
rect 19533 34017 19567 34051
rect 20637 34017 20671 34051
rect 22937 34017 22971 34051
rect 23765 34017 23799 34051
rect 25053 34017 25087 34051
rect 35541 34017 35575 34051
rect 38209 34017 38243 34051
rect 38485 34017 38519 34051
rect 38694 34017 38728 34051
rect 40509 34017 40543 34051
rect 48145 34017 48179 34051
rect 10885 33949 10919 33983
rect 11069 33949 11103 33983
rect 11897 33949 11931 33983
rect 13185 33949 13219 33983
rect 14289 33949 14323 33983
rect 14473 33949 14507 33983
rect 15117 33949 15151 33983
rect 15209 33949 15243 33983
rect 16037 33949 16071 33983
rect 16221 33949 16255 33983
rect 16681 33949 16715 33983
rect 17785 33949 17819 33983
rect 18613 33949 18647 33983
rect 19625 33949 19659 33983
rect 20545 33949 20579 33983
rect 21465 33949 21499 33983
rect 21557 33949 21591 33983
rect 22845 33949 22879 33983
rect 24777 33949 24811 33983
rect 26801 33949 26835 33983
rect 26985 33949 27019 33983
rect 27997 33949 28031 33983
rect 28457 33949 28491 33983
rect 30021 33949 30055 33983
rect 30205 33949 30239 33983
rect 30481 33949 30515 33983
rect 31309 33949 31343 33983
rect 33517 33949 33551 33983
rect 34897 33949 34931 33983
rect 35081 33949 35115 33983
rect 35817 33949 35851 33983
rect 36277 33949 36311 33983
rect 36461 33949 36495 33983
rect 37381 33949 37415 33983
rect 37473 33949 37507 33983
rect 38577 33949 38611 33983
rect 41429 33949 41463 33983
rect 47869 33949 47903 33983
rect 10977 33881 11011 33915
rect 15393 33881 15427 33915
rect 17601 33881 17635 33915
rect 20821 33881 20855 33915
rect 28733 33881 28767 33915
rect 30113 33881 30147 33915
rect 30323 33881 30357 33915
rect 31125 33881 31159 33915
rect 37565 33881 37599 33915
rect 9781 33813 9815 33847
rect 12173 33813 12207 33847
rect 17141 33813 17175 33847
rect 19257 33813 19291 33847
rect 20545 33813 20579 33847
rect 26985 33813 27019 33847
rect 27629 33813 27663 33847
rect 28549 33813 28583 33847
rect 30941 33813 30975 33847
rect 32873 33813 32907 33847
rect 33977 33813 34011 33847
rect 37749 33813 37783 33847
rect 43177 33813 43211 33847
rect 11897 33609 11931 33643
rect 13730 33609 13764 33643
rect 15577 33609 15611 33643
rect 16865 33609 16899 33643
rect 17509 33609 17543 33643
rect 19257 33609 19291 33643
rect 21005 33609 21039 33643
rect 21189 33609 21223 33643
rect 24317 33609 24351 33643
rect 28181 33609 28215 33643
rect 28733 33609 28767 33643
rect 29745 33609 29779 33643
rect 31309 33609 31343 33643
rect 34253 33609 34287 33643
rect 36185 33609 36219 33643
rect 37289 33609 37323 33643
rect 38669 33609 38703 33643
rect 48145 33609 48179 33643
rect 10425 33541 10459 33575
rect 11713 33541 11747 33575
rect 12725 33541 12759 33575
rect 12909 33541 12943 33575
rect 13645 33541 13679 33575
rect 16681 33541 16715 33575
rect 19717 33541 19751 33575
rect 20361 33541 20395 33575
rect 22385 33541 22419 33575
rect 22937 33541 22971 33575
rect 24225 33541 24259 33575
rect 33701 33541 33735 33575
rect 35633 33541 35667 33575
rect 37657 33541 37691 33575
rect 38485 33541 38519 33575
rect 39497 33541 39531 33575
rect 42993 33541 43027 33575
rect 9873 33473 9907 33507
rect 10977 33473 11011 33507
rect 11529 33473 11563 33507
rect 13553 33473 13587 33507
rect 13829 33473 13863 33507
rect 14841 33473 14875 33507
rect 15025 33473 15059 33507
rect 15485 33473 15519 33507
rect 15669 33473 15703 33507
rect 16957 33473 16991 33507
rect 17969 33473 18003 33507
rect 18153 33473 18187 33507
rect 19073 33473 19107 33507
rect 20821 33473 20855 33507
rect 20913 33473 20947 33507
rect 22845 33473 22879 33507
rect 23029 33473 23063 33507
rect 24133 33473 24167 33507
rect 24409 33473 24443 33507
rect 24869 33473 24903 33507
rect 24961 33473 24995 33507
rect 25145 33473 25179 33507
rect 25605 33473 25639 33507
rect 25789 33473 25823 33507
rect 27353 33473 27387 33507
rect 27445 33473 27479 33507
rect 27721 33473 27755 33507
rect 30389 33473 30423 33507
rect 31217 33473 31251 33507
rect 31401 33473 31435 33507
rect 32321 33473 32355 33507
rect 32413 33473 32447 33507
rect 32597 33473 32631 33507
rect 34621 33473 34655 33507
rect 35449 33473 35483 33507
rect 36093 33473 36127 33507
rect 36277 33473 36311 33507
rect 37473 33473 37507 33507
rect 37565 33473 37599 33507
rect 37841 33473 37875 33507
rect 38301 33473 38335 33507
rect 39129 33473 39163 33507
rect 39313 33473 39347 33507
rect 39589 33473 39623 33507
rect 39957 33473 39991 33507
rect 40693 33473 40727 33507
rect 40782 33473 40816 33507
rect 40877 33473 40911 33507
rect 41061 33473 41095 33507
rect 14381 33405 14415 33439
rect 18613 33405 18647 33439
rect 18981 33405 19015 33439
rect 20085 33405 20119 33439
rect 20177 33405 20211 33439
rect 21189 33405 21223 33439
rect 27537 33405 27571 33439
rect 30481 33405 30515 33439
rect 30757 33405 30791 33439
rect 34529 33405 34563 33439
rect 35265 33405 35299 33439
rect 16681 33337 16715 33371
rect 23581 33337 23615 33371
rect 25145 33337 25179 33371
rect 27721 33337 27755 33371
rect 41521 33337 41555 33371
rect 13093 33269 13127 33303
rect 15025 33269 15059 33303
rect 18061 33269 18095 33303
rect 25697 33269 25731 33303
rect 26433 33269 26467 33303
rect 32597 33269 32631 33303
rect 33149 33269 33183 33303
rect 34529 33269 34563 33303
rect 40417 33269 40451 33303
rect 42441 33269 42475 33303
rect 43637 33269 43671 33303
rect 11621 33065 11655 33099
rect 12633 33065 12667 33099
rect 14933 33065 14967 33099
rect 20177 33065 20211 33099
rect 20729 33065 20763 33099
rect 22477 33065 22511 33099
rect 22845 33065 22879 33099
rect 23397 33065 23431 33099
rect 24869 33065 24903 33099
rect 30297 33065 30331 33099
rect 33517 33065 33551 33099
rect 36185 33065 36219 33099
rect 36737 33065 36771 33099
rect 37473 33065 37507 33099
rect 38117 33065 38151 33099
rect 40877 33065 40911 33099
rect 16313 32997 16347 33031
rect 25973 32997 26007 33031
rect 31217 32997 31251 33031
rect 32321 32997 32355 33031
rect 35633 32997 35667 33031
rect 41429 32997 41463 33031
rect 42533 32997 42567 33031
rect 10517 32929 10551 32963
rect 19809 32929 19843 32963
rect 21833 32929 21867 32963
rect 25697 32929 25731 32963
rect 31677 32929 31711 32963
rect 11529 32861 11563 32895
rect 11713 32861 11747 32895
rect 12817 32861 12851 32895
rect 12909 32861 12943 32895
rect 13093 32861 13127 32895
rect 13185 32861 13219 32895
rect 15393 32861 15427 32895
rect 15577 32861 15611 32895
rect 15945 32861 15979 32895
rect 16129 32861 16163 32895
rect 16405 32861 16439 32895
rect 17049 32861 17083 32895
rect 17325 32861 17359 32895
rect 17509 32861 17543 32895
rect 17969 32861 18003 32895
rect 18153 32861 18187 32895
rect 19993 32861 20027 32895
rect 20729 32861 20763 32895
rect 20913 32861 20947 32895
rect 21747 32861 21781 32895
rect 21925 32861 21959 32895
rect 22385 32861 22419 32895
rect 22661 32861 22695 32895
rect 23305 32861 23339 32895
rect 23489 32861 23523 32895
rect 24777 32861 24811 32895
rect 24961 32861 24995 32895
rect 25605 32861 25639 32895
rect 26709 32861 26743 32895
rect 26893 32861 26927 32895
rect 27537 32861 27571 32895
rect 28365 32861 28399 32895
rect 28549 32861 28583 32895
rect 30481 32861 30515 32895
rect 30573 32861 30607 32895
rect 31585 32861 31619 32895
rect 32505 32861 32539 32895
rect 32597 32861 32631 32895
rect 32781 32861 32815 32895
rect 32873 32861 32907 32895
rect 34989 32861 35023 32895
rect 35173 32861 35207 32895
rect 37473 32861 37507 32895
rect 37657 32861 37691 32895
rect 38117 32861 38151 32895
rect 38301 32861 38335 32895
rect 40049 32861 40083 32895
rect 40141 32861 40175 32895
rect 40325 32861 40359 32895
rect 40417 32861 40451 32895
rect 33471 32827 33505 32861
rect 16865 32793 16899 32827
rect 18705 32793 18739 32827
rect 27353 32793 27387 32827
rect 33701 32793 33735 32827
rect 39865 32793 39899 32827
rect 11069 32725 11103 32759
rect 14381 32725 14415 32759
rect 18061 32725 18095 32759
rect 19349 32725 19383 32759
rect 26801 32725 26835 32759
rect 27721 32725 27755 32759
rect 28733 32725 28767 32759
rect 29653 32725 29687 32759
rect 33333 32725 33367 32759
rect 35081 32725 35115 32759
rect 38761 32725 38795 32759
rect 41981 32725 42015 32759
rect 10425 32521 10459 32555
rect 16681 32521 16715 32555
rect 18261 32521 18295 32555
rect 18429 32521 18463 32555
rect 22569 32521 22603 32555
rect 24593 32521 24627 32555
rect 25973 32521 26007 32555
rect 28917 32521 28951 32555
rect 29561 32521 29595 32555
rect 31493 32521 31527 32555
rect 32505 32521 32539 32555
rect 33609 32521 33643 32555
rect 33977 32521 34011 32555
rect 34989 32521 35023 32555
rect 36461 32521 36495 32555
rect 38117 32521 38151 32555
rect 40049 32521 40083 32555
rect 14473 32453 14507 32487
rect 15301 32453 15335 32487
rect 18061 32453 18095 32487
rect 23213 32453 23247 32487
rect 24685 32453 24719 32487
rect 29837 32453 29871 32487
rect 30757 32453 30791 32487
rect 30941 32453 30975 32487
rect 32664 32453 32698 32487
rect 39497 32453 39531 32487
rect 1869 32385 1903 32419
rect 12633 32385 12667 32419
rect 12725 32385 12759 32419
rect 12909 32385 12943 32419
rect 13737 32385 13771 32419
rect 14381 32385 14415 32419
rect 14565 32385 14599 32419
rect 16865 32385 16899 32419
rect 19073 32385 19107 32419
rect 19257 32385 19291 32419
rect 19901 32385 19935 32419
rect 20085 32385 20119 32419
rect 21097 32385 21131 32419
rect 21281 32385 21315 32419
rect 21925 32385 21959 32419
rect 22385 32385 22419 32419
rect 22569 32385 22603 32419
rect 23397 32385 23431 32419
rect 23489 32385 23523 32419
rect 24593 32385 24627 32419
rect 24869 32385 24903 32419
rect 25513 32385 25547 32419
rect 25973 32385 26007 32419
rect 26157 32385 26191 32419
rect 26985 32385 27019 32419
rect 27169 32385 27203 32419
rect 27905 32385 27939 32419
rect 28089 32385 28123 32419
rect 28641 32385 28675 32419
rect 28825 32385 28859 32419
rect 29745 32385 29779 32419
rect 29929 32385 29963 32419
rect 30113 32385 30147 32419
rect 30205 32385 30239 32419
rect 30665 32385 30699 32419
rect 32781 32385 32815 32419
rect 33793 32385 33827 32419
rect 34069 32385 34103 32419
rect 34805 32385 34839 32419
rect 35081 32385 35115 32419
rect 35725 32385 35759 32419
rect 36369 32385 36403 32419
rect 36553 32385 36587 32419
rect 37473 32385 37507 32419
rect 37657 32385 37691 32419
rect 38301 32385 38335 32419
rect 40601 32385 40635 32419
rect 47869 32385 47903 32419
rect 13921 32317 13955 32351
rect 15853 32317 15887 32351
rect 17049 32317 17083 32351
rect 25421 32317 25455 32351
rect 27813 32317 27847 32351
rect 27997 32317 28031 32351
rect 32873 32317 32907 32351
rect 33149 32317 33183 32351
rect 34621 32317 34655 32351
rect 35909 32317 35943 32351
rect 38485 32317 38519 32351
rect 41705 32317 41739 32351
rect 12817 32249 12851 32283
rect 13093 32249 13127 32283
rect 18889 32249 18923 32283
rect 23673 32249 23707 32283
rect 27077 32249 27111 32283
rect 30941 32249 30975 32283
rect 38945 32249 38979 32283
rect 1961 32181 1995 32215
rect 10885 32181 10919 32215
rect 11989 32181 12023 32215
rect 13553 32181 13587 32215
rect 17509 32181 17543 32215
rect 18245 32181 18279 32215
rect 19993 32181 20027 32215
rect 20913 32181 20947 32215
rect 21097 32181 21131 32215
rect 23213 32181 23247 32215
rect 27629 32181 27663 32215
rect 29101 32181 29135 32215
rect 35541 32181 35575 32215
rect 37289 32181 37323 32215
rect 41153 32181 41187 32215
rect 48053 32181 48087 32215
rect 1593 31977 1627 32011
rect 10701 31977 10735 32011
rect 11345 31977 11379 32011
rect 11805 31977 11839 32011
rect 12633 31977 12667 32011
rect 14289 31977 14323 32011
rect 15025 31977 15059 32011
rect 15945 31977 15979 32011
rect 16589 31977 16623 32011
rect 19257 31977 19291 32011
rect 20453 31977 20487 32011
rect 22845 31977 22879 32011
rect 23397 31977 23431 32011
rect 24501 31977 24535 32011
rect 25605 31977 25639 32011
rect 27905 31977 27939 32011
rect 29009 31977 29043 32011
rect 30113 31977 30147 32011
rect 31861 31977 31895 32011
rect 32781 31977 32815 32011
rect 34161 31977 34195 32011
rect 34805 31977 34839 32011
rect 39865 31977 39899 32011
rect 40417 31977 40451 32011
rect 40969 31977 41003 32011
rect 47685 31977 47719 32011
rect 17141 31909 17175 31943
rect 20821 31909 20855 31943
rect 22017 31909 22051 31943
rect 25145 31909 25179 31943
rect 20729 31841 20763 31875
rect 22477 31841 22511 31875
rect 23581 31841 23615 31875
rect 24409 31841 24443 31875
rect 25973 31841 26007 31875
rect 27169 31841 27203 31875
rect 28641 31841 28675 31875
rect 28733 31841 28767 31875
rect 29653 31841 29687 31875
rect 29745 31841 29779 31875
rect 29929 31841 29963 31875
rect 30665 31841 30699 31875
rect 32229 31841 32263 31875
rect 33885 31841 33919 31875
rect 34069 31841 34103 31875
rect 36553 31841 36587 31875
rect 38209 31841 38243 31875
rect 38669 31841 38703 31875
rect 10241 31773 10275 31807
rect 12357 31773 12391 31807
rect 12449 31773 12483 31807
rect 12633 31773 12667 31807
rect 13369 31773 13403 31807
rect 14105 31773 14139 31807
rect 14197 31773 14231 31807
rect 14381 31773 14415 31807
rect 15669 31773 15703 31807
rect 15761 31773 15795 31807
rect 17141 31773 17175 31807
rect 17417 31773 17451 31807
rect 18245 31773 18279 31807
rect 18337 31773 18371 31807
rect 18521 31773 18555 31807
rect 19257 31773 19291 31807
rect 19441 31773 19475 31807
rect 20637 31773 20671 31807
rect 20913 31773 20947 31807
rect 21097 31773 21131 31807
rect 21649 31773 21683 31807
rect 22661 31773 22695 31807
rect 23305 31773 23339 31807
rect 24869 31773 24903 31807
rect 25789 31773 25823 31807
rect 26985 31773 27019 31807
rect 27629 31773 27663 31807
rect 27905 31773 27939 31807
rect 28549 31773 28583 31807
rect 28825 31773 28859 31807
rect 29837 31773 29871 31807
rect 30573 31773 30607 31807
rect 30757 31773 30791 31807
rect 32137 31773 32171 31807
rect 32965 31773 32999 31807
rect 33057 31773 33091 31807
rect 34161 31773 34195 31807
rect 35061 31773 35095 31807
rect 35154 31773 35188 31807
rect 35265 31773 35299 31807
rect 35449 31773 35483 31807
rect 36737 31773 36771 31807
rect 37197 31773 37231 31807
rect 37473 31773 37507 31807
rect 39221 31773 39255 31807
rect 13185 31705 13219 31739
rect 15009 31705 15043 31739
rect 15209 31705 15243 31739
rect 15945 31705 15979 31739
rect 21833 31705 21867 31739
rect 24685 31705 24719 31739
rect 26801 31705 26835 31739
rect 36277 31705 36311 31739
rect 13553 31637 13587 31671
rect 14841 31637 14875 31671
rect 17325 31637 17359 31671
rect 17877 31637 17911 31671
rect 19993 31637 20027 31671
rect 23857 31637 23891 31671
rect 24777 31637 24811 31671
rect 27721 31637 27755 31671
rect 31309 31637 31343 31671
rect 10977 31433 11011 31467
rect 13553 31433 13587 31467
rect 13921 31433 13955 31467
rect 16865 31433 16899 31467
rect 17877 31433 17911 31467
rect 19809 31433 19843 31467
rect 21097 31433 21131 31467
rect 23397 31433 23431 31467
rect 24225 31433 24259 31467
rect 25513 31433 25547 31467
rect 27635 31433 27669 31467
rect 28365 31433 28399 31467
rect 29009 31433 29043 31467
rect 29469 31433 29503 31467
rect 31033 31433 31067 31467
rect 32321 31433 32355 31467
rect 35541 31433 35575 31467
rect 37657 31433 37691 31467
rect 38853 31433 38887 31467
rect 40509 31433 40543 31467
rect 12357 31365 12391 31399
rect 20637 31365 20671 31399
rect 22477 31365 22511 31399
rect 22845 31365 22879 31399
rect 24685 31365 24719 31399
rect 25053 31365 25087 31399
rect 27721 31365 27755 31399
rect 32597 31365 32631 31399
rect 11897 31297 11931 31331
rect 12541 31297 12575 31331
rect 13461 31297 13495 31331
rect 13737 31297 13771 31331
rect 14841 31297 14875 31331
rect 15025 31297 15059 31331
rect 15117 31297 15151 31331
rect 15761 31297 15795 31331
rect 17417 31297 17451 31331
rect 17509 31297 17543 31331
rect 17693 31297 17727 31331
rect 18797 31297 18831 31331
rect 18981 31297 19015 31331
rect 19717 31297 19751 31331
rect 19901 31297 19935 31331
rect 20913 31297 20947 31331
rect 22661 31297 22695 31331
rect 23305 31297 23339 31331
rect 23489 31297 23523 31331
rect 24869 31297 24903 31331
rect 25513 31297 25547 31331
rect 25697 31297 25731 31331
rect 26157 31297 26191 31331
rect 26341 31297 26375 31331
rect 27537 31297 27571 31331
rect 27813 31297 27847 31331
rect 28273 31297 28307 31331
rect 28457 31297 28491 31331
rect 29929 31297 29963 31331
rect 30389 31297 30423 31331
rect 30573 31297 30607 31331
rect 31033 31297 31067 31331
rect 31217 31297 31251 31331
rect 32505 31297 32539 31331
rect 32689 31297 32723 31331
rect 32807 31297 32841 31331
rect 33425 31297 33459 31331
rect 34069 31297 34103 31331
rect 35173 31297 35207 31331
rect 37473 31297 37507 31331
rect 37749 31297 37783 31331
rect 15577 31229 15611 31263
rect 19257 31229 19291 31263
rect 20729 31229 20763 31263
rect 32965 31229 32999 31263
rect 33517 31229 33551 31263
rect 34253 31229 34287 31263
rect 35265 31229 35299 31263
rect 15117 31161 15151 31195
rect 18981 31161 19015 31195
rect 12725 31093 12759 31127
rect 15945 31093 15979 31127
rect 20637 31093 20671 31127
rect 22017 31093 22051 31127
rect 26157 31093 26191 31127
rect 27077 31093 27111 31127
rect 29653 31093 29687 31127
rect 30389 31093 30423 31127
rect 36093 31093 36127 31127
rect 36553 31093 36587 31127
rect 37289 31093 37323 31127
rect 38301 31093 38335 31127
rect 39313 31093 39347 31127
rect 39865 31093 39899 31127
rect 14105 30889 14139 30923
rect 15209 30889 15243 30923
rect 16589 30889 16623 30923
rect 17417 30889 17451 30923
rect 18705 30889 18739 30923
rect 19993 30889 20027 30923
rect 20637 30889 20671 30923
rect 20821 30889 20855 30923
rect 21373 30889 21407 30923
rect 22385 30889 22419 30923
rect 27537 30889 27571 30923
rect 29653 30889 29687 30923
rect 30757 30889 30791 30923
rect 33517 30889 33551 30923
rect 37105 30889 37139 30923
rect 38209 30889 38243 30923
rect 38761 30889 38795 30923
rect 14473 30821 14507 30855
rect 16497 30821 16531 30855
rect 28365 30821 28399 30855
rect 11897 30753 11931 30787
rect 13093 30753 13127 30787
rect 14197 30753 14231 30787
rect 21741 30753 21775 30787
rect 22293 30753 22327 30787
rect 32045 30753 32079 30787
rect 36553 30753 36587 30787
rect 11345 30685 11379 30719
rect 12357 30685 12391 30719
rect 12541 30685 12575 30719
rect 13001 30685 13035 30719
rect 13185 30685 13219 30719
rect 14105 30685 14139 30719
rect 15393 30685 15427 30719
rect 15669 30685 15703 30719
rect 17417 30685 17451 30719
rect 17693 30685 17727 30719
rect 19717 30685 19751 30719
rect 21649 30685 21683 30719
rect 22477 30685 22511 30719
rect 22569 30685 22603 30719
rect 24409 30685 24443 30719
rect 24593 30685 24627 30719
rect 26801 30685 26835 30719
rect 29561 30685 29595 30719
rect 29745 30685 29779 30719
rect 31125 30685 31159 30719
rect 32965 30685 32999 30719
rect 33517 30685 33551 30719
rect 33701 30685 33735 30719
rect 37657 30685 37691 30719
rect 12449 30617 12483 30651
rect 15577 30617 15611 30651
rect 16129 30617 16163 30651
rect 17509 30617 17543 30651
rect 19993 30617 20027 30651
rect 20453 30617 20487 30651
rect 20653 30617 20687 30651
rect 27721 30617 27755 30651
rect 27905 30617 27939 30651
rect 30941 30617 30975 30651
rect 35173 30617 35207 30651
rect 35357 30617 35391 30651
rect 19809 30549 19843 30583
rect 23121 30549 23155 30583
rect 23765 30549 23799 30583
rect 24501 30549 24535 30583
rect 25145 30549 25179 30583
rect 26065 30549 26099 30583
rect 26893 30549 26927 30583
rect 29009 30549 29043 30583
rect 30205 30549 30239 30583
rect 35541 30549 35575 30583
rect 36001 30549 36035 30583
rect 12081 30345 12115 30379
rect 12541 30345 12575 30379
rect 13737 30345 13771 30379
rect 15393 30345 15427 30379
rect 17141 30345 17175 30379
rect 19625 30345 19659 30379
rect 20637 30345 20671 30379
rect 22293 30345 22327 30379
rect 24961 30345 24995 30379
rect 32321 30345 32355 30379
rect 32689 30345 32723 30379
rect 35265 30345 35299 30379
rect 37289 30345 37323 30379
rect 2053 30277 2087 30311
rect 17601 30277 17635 30311
rect 21143 30277 21177 30311
rect 27813 30277 27847 30311
rect 31585 30277 31619 30311
rect 33517 30277 33551 30311
rect 1869 30209 1903 30243
rect 13185 30209 13219 30243
rect 14289 30209 14323 30243
rect 15301 30209 15335 30243
rect 15577 30209 15611 30243
rect 16681 30209 16715 30243
rect 16773 30209 16807 30243
rect 16957 30209 16991 30243
rect 17785 30209 17819 30243
rect 18889 30209 18923 30243
rect 19073 30209 19107 30243
rect 19533 30209 19567 30243
rect 19717 30209 19751 30243
rect 19809 30209 19843 30243
rect 20821 30209 20855 30243
rect 20913 30209 20947 30243
rect 21005 30209 21039 30243
rect 21281 30209 21315 30243
rect 23029 30209 23063 30243
rect 24041 30209 24075 30243
rect 24869 30209 24903 30243
rect 25145 30209 25179 30243
rect 25789 30209 25823 30243
rect 25973 30209 26007 30243
rect 27537 30209 27571 30243
rect 28273 30209 28307 30243
rect 28365 30209 28399 30243
rect 28549 30209 28583 30243
rect 29101 30209 29135 30243
rect 29837 30209 29871 30243
rect 30297 30209 30331 30243
rect 30481 30209 30515 30243
rect 31401 30209 31435 30243
rect 32229 30209 32263 30243
rect 32505 30209 32539 30243
rect 33425 30209 33459 30243
rect 33609 30209 33643 30243
rect 34069 30209 34103 30243
rect 34253 30209 34287 30243
rect 34897 30209 34931 30243
rect 36369 30209 36403 30243
rect 15761 30141 15795 30175
rect 23949 30141 23983 30175
rect 24409 30141 24443 30175
rect 27813 30141 27847 30175
rect 29561 30141 29595 30175
rect 31217 30141 31251 30175
rect 34805 30141 34839 30175
rect 36461 30141 36495 30175
rect 36737 30141 36771 30175
rect 18981 30073 19015 30107
rect 25881 30073 25915 30107
rect 28549 30073 28583 30107
rect 14841 30005 14875 30039
rect 17969 30005 18003 30039
rect 25329 30005 25363 30039
rect 26985 30005 27019 30039
rect 27629 30005 27663 30039
rect 29653 30005 29687 30039
rect 29745 30005 29779 30039
rect 30297 30005 30331 30039
rect 34161 30005 34195 30039
rect 1593 29801 1627 29835
rect 15025 29801 15059 29835
rect 16037 29801 16071 29835
rect 16221 29801 16255 29835
rect 16957 29801 16991 29835
rect 17785 29801 17819 29835
rect 18521 29801 18555 29835
rect 18705 29801 18739 29835
rect 19809 29801 19843 29835
rect 21189 29801 21223 29835
rect 22845 29801 22879 29835
rect 23029 29801 23063 29835
rect 26893 29801 26927 29835
rect 27721 29801 27755 29835
rect 28917 29801 28951 29835
rect 29561 29801 29595 29835
rect 30481 29801 30515 29835
rect 30665 29801 30699 29835
rect 31309 29801 31343 29835
rect 34161 29801 34195 29835
rect 34805 29801 34839 29835
rect 36093 29801 36127 29835
rect 14473 29733 14507 29767
rect 25513 29733 25547 29767
rect 35357 29733 35391 29767
rect 25237 29665 25271 29699
rect 26985 29665 27019 29699
rect 33149 29665 33183 29699
rect 35909 29665 35943 29699
rect 48145 29665 48179 29699
rect 16865 29597 16899 29631
rect 17049 29597 17083 29631
rect 19349 29597 19383 29631
rect 19625 29597 19659 29631
rect 20453 29597 20487 29631
rect 20637 29597 20671 29631
rect 21189 29597 21223 29631
rect 21373 29597 21407 29631
rect 21833 29597 21867 29631
rect 22017 29597 22051 29631
rect 23489 29597 23523 29631
rect 23581 29597 23615 29631
rect 23765 29597 23799 29631
rect 25145 29597 25179 29631
rect 26525 29597 26559 29631
rect 26801 29597 26835 29631
rect 27905 29597 27939 29631
rect 28181 29597 28215 29631
rect 28365 29597 28399 29631
rect 29009 29597 29043 29631
rect 29561 29597 29595 29631
rect 29837 29597 29871 29631
rect 31309 29597 31343 29631
rect 31493 29597 31527 29631
rect 32505 29597 32539 29631
rect 32689 29597 32723 29631
rect 33609 29597 33643 29631
rect 35817 29597 35851 29631
rect 36737 29597 36771 29631
rect 36829 29597 36863 29631
rect 47869 29597 47903 29631
rect 16175 29563 16209 29597
rect 16405 29529 16439 29563
rect 18337 29529 18371 29563
rect 22661 29529 22695 29563
rect 30297 29529 30331 29563
rect 32597 29529 32631 29563
rect 35357 29529 35391 29563
rect 15485 29461 15519 29495
rect 18537 29461 18571 29495
rect 19441 29461 19475 29495
rect 20269 29461 20303 29495
rect 21925 29461 21959 29495
rect 22861 29461 22895 29495
rect 23666 29461 23700 29495
rect 24409 29461 24443 29495
rect 25973 29461 26007 29495
rect 26617 29461 26651 29495
rect 27261 29461 27295 29495
rect 29745 29461 29779 29495
rect 30507 29461 30541 29495
rect 32045 29461 32079 29495
rect 33425 29461 33459 29495
rect 33517 29461 33551 29495
rect 36553 29461 36587 29495
rect 16129 29257 16163 29291
rect 17049 29257 17083 29291
rect 17693 29257 17727 29291
rect 18889 29257 18923 29291
rect 19257 29257 19291 29291
rect 19809 29257 19843 29291
rect 21005 29257 21039 29291
rect 22569 29257 22603 29291
rect 23305 29257 23339 29291
rect 23857 29257 23891 29291
rect 27077 29257 27111 29291
rect 27169 29257 27203 29291
rect 28273 29257 28307 29291
rect 28457 29257 28491 29291
rect 30481 29257 30515 29291
rect 30941 29257 30975 29291
rect 33241 29257 33275 29291
rect 35173 29257 35207 29291
rect 35817 29257 35851 29291
rect 48145 29257 48179 29291
rect 16681 29189 16715 29223
rect 20637 29189 20671 29223
rect 20853 29189 20887 29223
rect 29469 29189 29503 29223
rect 32873 29189 32907 29223
rect 36277 29189 36311 29223
rect 15945 29121 15979 29155
rect 16129 29121 16163 29155
rect 16865 29121 16899 29155
rect 17601 29121 17635 29155
rect 17969 29121 18003 29155
rect 18797 29121 18831 29155
rect 19073 29121 19107 29155
rect 19717 29121 19751 29155
rect 19993 29121 20027 29155
rect 22201 29121 22235 29155
rect 23029 29121 23063 29155
rect 23765 29121 23799 29155
rect 23949 29121 23983 29155
rect 24501 29121 24535 29155
rect 24593 29121 24627 29155
rect 24777 29121 24811 29155
rect 25605 29121 25639 29155
rect 25697 29121 25731 29155
rect 26985 29121 27019 29155
rect 28089 29121 28123 29155
rect 28181 29121 28215 29155
rect 29377 29121 29411 29155
rect 29653 29121 29687 29155
rect 30113 29121 30147 29155
rect 30205 29121 30239 29155
rect 31217 29121 31251 29155
rect 33057 29121 33091 29155
rect 34345 29121 34379 29155
rect 35449 29121 35483 29155
rect 17877 29053 17911 29087
rect 22293 29053 22327 29087
rect 23305 29053 23339 29087
rect 24961 29053 24995 29087
rect 25421 29053 25455 29087
rect 27445 29053 27479 29087
rect 30941 29053 30975 29087
rect 34253 29053 34287 29087
rect 34437 29053 34471 29087
rect 34529 29053 34563 29087
rect 35357 29053 35391 29087
rect 14841 28985 14875 29019
rect 15393 28985 15427 29019
rect 18061 28985 18095 29019
rect 25513 28985 25547 29019
rect 27905 28985 27939 29019
rect 31125 28985 31159 29019
rect 18337 28917 18371 28951
rect 19993 28917 20027 28951
rect 20821 28917 20855 28951
rect 22385 28917 22419 28951
rect 23121 28917 23155 28951
rect 26433 28917 26467 28951
rect 29653 28917 29687 28951
rect 30113 28917 30147 28951
rect 32137 28917 32171 28951
rect 34713 28917 34747 28951
rect 15301 28713 15335 28747
rect 18061 28713 18095 28747
rect 19441 28713 19475 28747
rect 20085 28713 20119 28747
rect 23397 28713 23431 28747
rect 25053 28713 25087 28747
rect 26341 28713 26375 28747
rect 29653 28713 29687 28747
rect 30297 28713 30331 28747
rect 32965 28713 32999 28747
rect 35817 28713 35851 28747
rect 18613 28645 18647 28679
rect 21005 28645 21039 28679
rect 25973 28645 26007 28679
rect 35265 28645 35299 28679
rect 20545 28577 20579 28611
rect 21097 28577 21131 28611
rect 21649 28577 21683 28611
rect 22477 28577 22511 28611
rect 24593 28577 24627 28611
rect 27905 28577 27939 28611
rect 28089 28577 28123 28611
rect 28181 28577 28215 28611
rect 28365 28577 28399 28611
rect 30665 28577 30699 28611
rect 32597 28577 32631 28611
rect 34805 28577 34839 28611
rect 17601 28509 17635 28543
rect 17693 28509 17727 28543
rect 17877 28509 17911 28543
rect 19349 28509 19383 28543
rect 19533 28509 19567 28543
rect 20729 28509 20763 28543
rect 22017 28509 22051 28543
rect 22661 28509 22695 28543
rect 24685 28509 24719 28543
rect 26249 28509 26283 28543
rect 26341 28509 26375 28543
rect 26985 28509 27019 28543
rect 27997 28509 28031 28543
rect 29561 28509 29595 28543
rect 29745 28509 29779 28543
rect 30481 28509 30515 28543
rect 31723 28509 31757 28543
rect 31861 28509 31895 28543
rect 31974 28509 32008 28543
rect 32137 28509 32171 28543
rect 33057 28509 33091 28543
rect 34897 28509 34931 28543
rect 35725 28509 35759 28543
rect 21833 28441 21867 28475
rect 22845 28441 22879 28475
rect 26801 28441 26835 28475
rect 31493 28441 31527 28475
rect 33517 28441 33551 28475
rect 15761 28373 15795 28407
rect 16497 28373 16531 28407
rect 17141 28373 17175 28407
rect 27169 28373 27203 28407
rect 28825 28373 28859 28407
rect 34161 28373 34195 28407
rect 18429 28169 18463 28203
rect 19073 28169 19107 28203
rect 27997 28169 28031 28203
rect 28641 28169 28675 28203
rect 30297 28169 30331 28203
rect 30941 28169 30975 28203
rect 32229 28169 32263 28203
rect 34069 28169 34103 28203
rect 35173 28169 35207 28203
rect 18337 28101 18371 28135
rect 18521 28101 18555 28135
rect 21281 28101 21315 28135
rect 25145 28101 25179 28135
rect 26065 28101 26099 28135
rect 31493 28101 31527 28135
rect 33793 28101 33827 28135
rect 33977 28101 34011 28135
rect 34529 28101 34563 28135
rect 1685 28033 1719 28067
rect 18245 28033 18279 28067
rect 19257 28033 19291 28067
rect 19349 28033 19383 28067
rect 19533 28033 19567 28067
rect 19717 28033 19751 28067
rect 20637 28033 20671 28067
rect 22293 28033 22327 28067
rect 22845 28033 22879 28067
rect 23029 28033 23063 28067
rect 23673 28033 23707 28067
rect 23857 28033 23891 28067
rect 24869 28033 24903 28067
rect 25973 28033 26007 28067
rect 26249 28033 26283 28067
rect 27629 28033 27663 28067
rect 28457 28033 28491 28067
rect 28641 28033 28675 28067
rect 30205 28033 30239 28067
rect 30389 28033 30423 28067
rect 30849 28033 30883 28067
rect 31033 28033 31067 28067
rect 32873 28033 32907 28067
rect 33241 28033 33275 28067
rect 34069 28033 34103 28067
rect 20177 27965 20211 27999
rect 23489 27965 23523 27999
rect 25145 27965 25179 27999
rect 27721 27965 27755 27999
rect 29745 27965 29779 27999
rect 1501 27897 1535 27931
rect 2237 27897 2271 27931
rect 17785 27897 17819 27931
rect 19441 27897 19475 27931
rect 24409 27897 24443 27931
rect 26249 27897 26283 27931
rect 20361 27829 20395 27863
rect 23029 27829 23063 27863
rect 24961 27829 24995 27863
rect 29101 27829 29135 27863
rect 19809 27625 19843 27659
rect 21833 27625 21867 27659
rect 26249 27625 26283 27659
rect 26433 27625 26467 27659
rect 28089 27625 28123 27659
rect 30573 27625 30607 27659
rect 32229 27625 32263 27659
rect 18613 27557 18647 27591
rect 21005 27557 21039 27591
rect 22017 27557 22051 27591
rect 23121 27557 23155 27591
rect 33517 27557 33551 27591
rect 27537 27489 27571 27523
rect 27997 27489 28031 27523
rect 33333 27489 33367 27523
rect 48145 27489 48179 27523
rect 19717 27421 19751 27455
rect 19901 27421 19935 27455
rect 21557 27421 21591 27455
rect 22477 27421 22511 27455
rect 22661 27421 22695 27455
rect 22753 27421 22787 27455
rect 22845 27421 22879 27455
rect 23581 27421 23615 27455
rect 23765 27421 23799 27455
rect 25145 27421 25179 27455
rect 25329 27421 25363 27455
rect 27077 27421 27111 27455
rect 27353 27421 27387 27455
rect 28181 27421 28215 27455
rect 28273 27421 28307 27455
rect 28733 27421 28767 27455
rect 29561 27421 29595 27455
rect 31217 27421 31251 27455
rect 31401 27421 31435 27455
rect 32137 27421 32171 27455
rect 32321 27421 32355 27455
rect 33241 27421 33275 27455
rect 47869 27421 47903 27455
rect 23673 27353 23707 27387
rect 24501 27353 24535 27387
rect 26065 27353 26099 27387
rect 31033 27353 31067 27387
rect 20545 27285 20579 27319
rect 24961 27285 24995 27319
rect 26265 27285 26299 27319
rect 27169 27285 27203 27319
rect 32873 27285 32907 27319
rect 33977 27285 34011 27319
rect 18797 27081 18831 27115
rect 20177 27081 20211 27115
rect 21925 27081 21959 27115
rect 23397 27081 23431 27115
rect 26065 27081 26099 27115
rect 27077 27081 27111 27115
rect 31125 27081 31159 27115
rect 32321 27081 32355 27115
rect 48145 27081 48179 27115
rect 19717 27013 19751 27047
rect 20361 27013 20395 27047
rect 21189 27013 21223 27047
rect 24133 27013 24167 27047
rect 34161 27013 34195 27047
rect 20545 26945 20579 26979
rect 21097 26945 21131 26979
rect 21281 26945 21315 26979
rect 22109 26945 22143 26979
rect 23029 26945 23063 26979
rect 24041 26945 24075 26979
rect 24225 26945 24259 26979
rect 24869 26945 24903 26979
rect 25145 26945 25179 26979
rect 25697 26945 25731 26979
rect 25789 26945 25823 26979
rect 27445 26945 27479 26979
rect 28457 26945 28491 26979
rect 29469 26945 29503 26979
rect 30297 26945 30331 26979
rect 30481 26945 30515 26979
rect 30941 26945 30975 26979
rect 31125 26945 31159 26979
rect 32321 26945 32355 26979
rect 32505 26945 32539 26979
rect 22293 26877 22327 26911
rect 23121 26877 23155 26911
rect 27353 26877 27387 26911
rect 28549 26877 28583 26911
rect 29377 26877 29411 26911
rect 33333 26877 33367 26911
rect 24961 26809 24995 26843
rect 25053 26809 25087 26843
rect 28825 26809 28859 26843
rect 29837 26809 29871 26843
rect 24685 26741 24719 26775
rect 25697 26741 25731 26775
rect 30389 26741 30423 26775
rect 34713 26741 34747 26775
rect 19625 26537 19659 26571
rect 20177 26537 20211 26571
rect 20913 26537 20947 26571
rect 22937 26537 22971 26571
rect 23029 26537 23063 26571
rect 25053 26537 25087 26571
rect 26525 26537 26559 26571
rect 29837 26537 29871 26571
rect 31953 26537 31987 26571
rect 33609 26537 33643 26571
rect 25881 26469 25915 26503
rect 27169 26469 27203 26503
rect 22385 26401 22419 26435
rect 23121 26401 23155 26435
rect 30113 26401 30147 26435
rect 31125 26401 31159 26435
rect 33149 26401 33183 26435
rect 20085 26333 20119 26367
rect 20269 26333 20303 26367
rect 22201 26333 22235 26367
rect 22845 26333 22879 26367
rect 25421 26333 25455 26367
rect 25881 26333 25915 26367
rect 26065 26333 26099 26367
rect 30021 26333 30055 26367
rect 31493 26333 31527 26367
rect 32597 26333 32631 26367
rect 47869 26333 47903 26367
rect 48145 26333 48179 26367
rect 1869 26265 1903 26299
rect 2053 26265 2087 26299
rect 21465 26265 21499 26299
rect 22017 26265 22051 26299
rect 24593 26265 24627 26299
rect 25237 26265 25271 26299
rect 27721 26265 27755 26299
rect 28365 26265 28399 26299
rect 31309 26265 31343 26299
rect 30481 26197 30515 26231
rect 21833 25993 21867 26027
rect 30297 25993 30331 26027
rect 31033 25993 31067 26027
rect 32781 25993 32815 26027
rect 1593 25925 1627 25959
rect 48145 25925 48179 25959
rect 24593 25857 24627 25891
rect 24777 25857 24811 25891
rect 27261 25857 27295 25891
rect 29929 25857 29963 25891
rect 31033 25857 31067 25891
rect 31217 25857 31251 25891
rect 27169 25789 27203 25823
rect 27629 25789 27663 25823
rect 29837 25789 29871 25823
rect 20545 25653 20579 25687
rect 22477 25653 22511 25687
rect 24685 25653 24719 25687
rect 25513 25653 25547 25687
rect 26249 25653 26283 25687
rect 32137 25653 32171 25687
rect 25145 25449 25179 25483
rect 28181 25449 28215 25483
rect 28825 25449 28859 25483
rect 31309 25449 31343 25483
rect 31861 25449 31895 25483
rect 25789 25381 25823 25415
rect 27445 25381 27479 25415
rect 27537 25381 27571 25415
rect 24961 25313 24995 25347
rect 26801 25313 26835 25347
rect 27629 25313 27663 25347
rect 24869 25245 24903 25279
rect 26709 25245 26743 25279
rect 26893 25245 26927 25279
rect 27353 25245 27387 25279
rect 28089 25245 28123 25279
rect 28273 25245 28307 25279
rect 23489 25109 23523 25143
rect 24869 24905 24903 24939
rect 28089 24905 28123 24939
rect 23765 24769 23799 24803
rect 23949 24769 23983 24803
rect 24593 24769 24627 24803
rect 24961 24769 24995 24803
rect 25053 24769 25087 24803
rect 26433 24769 26467 24803
rect 27169 24769 27203 24803
rect 27353 24769 27387 24803
rect 27997 24769 28031 24803
rect 28181 24769 28215 24803
rect 28641 24769 28675 24803
rect 23305 24701 23339 24735
rect 24133 24701 24167 24735
rect 27537 24701 27571 24735
rect 2237 24361 2271 24395
rect 24501 24361 24535 24395
rect 25145 24361 25179 24395
rect 27721 24361 27755 24395
rect 28273 24361 28307 24395
rect 47777 24361 47811 24395
rect 1685 24157 1719 24191
rect 24409 24157 24443 24191
rect 24593 24157 24627 24191
rect 48053 24089 48087 24123
rect 1501 24021 1535 24055
rect 23765 24021 23799 24055
rect 27077 24021 27111 24055
rect 48145 23817 48179 23851
rect 47317 21981 47351 22015
rect 47869 21981 47903 22015
rect 1869 21913 1903 21947
rect 1961 21845 1995 21879
rect 48053 21845 48087 21879
rect 1593 21641 1627 21675
rect 47317 20009 47351 20043
rect 47869 19805 47903 19839
rect 1869 19737 1903 19771
rect 2145 19669 2179 19703
rect 48053 19669 48087 19703
rect 1685 19465 1719 19499
rect 1869 18241 1903 18275
rect 47869 18241 47903 18275
rect 1961 18037 1995 18071
rect 48053 18037 48087 18071
rect 47685 17833 47719 17867
rect 1593 17765 1627 17799
rect 47961 16201 47995 16235
rect 1869 16065 1903 16099
rect 48145 16065 48179 16099
rect 2145 15861 2179 15895
rect 1593 15657 1627 15691
rect 48145 15657 48179 15691
rect 1409 13889 1443 13923
rect 47869 13889 47903 13923
rect 1593 13753 1627 13787
rect 48053 13685 48087 13719
rect 1409 13481 1443 13515
rect 47777 13481 47811 13515
rect 47961 11849 47995 11883
rect 1685 11713 1719 11747
rect 48145 11713 48179 11747
rect 1501 11577 1535 11611
rect 2237 11577 2271 11611
rect 48145 11305 48179 11339
rect 47317 10013 47351 10047
rect 47869 10013 47903 10047
rect 1869 9945 1903 9979
rect 2145 9877 2179 9911
rect 48053 9877 48087 9911
rect 1593 9605 1627 9639
rect 47961 8041 47995 8075
rect 1685 7837 1719 7871
rect 2237 7837 2271 7871
rect 47409 7769 47443 7803
rect 48053 7769 48087 7803
rect 1501 7701 1535 7735
rect 1869 5593 1903 5627
rect 47869 5593 47903 5627
rect 48053 5593 48087 5627
rect 1961 5525 1995 5559
rect 47409 5525 47443 5559
rect 1593 5321 1627 5355
rect 47593 4097 47627 4131
rect 47317 3553 47351 3587
rect 1685 3485 1719 3519
rect 47869 3485 47903 3519
rect 2237 3417 2271 3451
rect 46857 3417 46891 3451
rect 1501 3349 1535 3383
rect 48053 3349 48087 3383
rect 32229 3145 32263 3179
rect 1409 3009 1443 3043
rect 2697 3009 2731 3043
rect 48145 3009 48179 3043
rect 4261 2941 4295 2975
rect 46581 2941 46615 2975
rect 1593 2873 1627 2907
rect 11989 2873 12023 2907
rect 47961 2873 47995 2907
rect 2145 2805 2179 2839
rect 9137 2805 9171 2839
rect 16865 2805 16899 2839
rect 19441 2805 19475 2839
rect 20637 2805 20671 2839
rect 24593 2805 24627 2839
rect 28365 2805 28399 2839
rect 39957 2805 39991 2839
rect 20913 2601 20947 2635
rect 28549 2601 28583 2635
rect 36369 2601 36403 2635
rect 45293 2601 45327 2635
rect 5457 2533 5491 2567
rect 7481 2533 7515 2567
rect 13277 2533 13311 2567
rect 19901 2533 19935 2567
rect 34897 2533 34931 2567
rect 37565 2533 37599 2567
rect 44189 2533 44223 2567
rect 1685 2465 1719 2499
rect 9597 2465 9631 2499
rect 22937 2465 22971 2499
rect 27261 2465 27295 2499
rect 30665 2465 30699 2499
rect 2145 2397 2179 2431
rect 4077 2397 4111 2431
rect 4813 2397 4847 2431
rect 5273 2397 5307 2431
rect 11805 2397 11839 2431
rect 15209 2397 15243 2431
rect 15669 2397 15703 2431
rect 19717 2397 19751 2431
rect 20729 2397 20763 2431
rect 22201 2397 22235 2431
rect 22661 2397 22695 2431
rect 26985 2397 27019 2431
rect 29929 2397 29963 2431
rect 30389 2397 30423 2431
rect 32597 2397 32631 2431
rect 34713 2397 34747 2431
rect 38117 2397 38151 2431
rect 40049 2397 40083 2431
rect 42441 2397 42475 2431
rect 45845 2397 45879 2431
rect 46765 2397 46799 2431
rect 47777 2397 47811 2431
rect 1501 2329 1535 2363
rect 2881 2329 2915 2363
rect 6745 2329 6779 2363
rect 7297 2329 7331 2363
rect 9413 2329 9447 2363
rect 12541 2329 12575 2363
rect 13093 2329 13127 2363
rect 17141 2329 17175 2363
rect 24869 2329 24903 2363
rect 28641 2329 28675 2363
rect 35725 2329 35759 2363
rect 36277 2329 36311 2363
rect 43453 2329 43487 2363
rect 44005 2329 44039 2363
rect 2329 2261 2363 2295
rect 3893 2261 3927 2295
rect 11621 2261 11655 2295
rect 15025 2261 15059 2295
rect 17233 2261 17267 2295
rect 24961 2261 24995 2295
rect 26433 2261 26467 2295
rect 32413 2261 32447 2295
rect 34161 2261 34195 2295
rect 38301 2261 38335 2295
rect 40233 2261 40267 2295
rect 41889 2261 41923 2295
rect 42625 2261 42659 2295
rect 46029 2261 46063 2295
rect 46949 2261 46983 2295
rect 47961 2261 47995 2295
<< metal1 >>
rect 21082 47744 21088 47796
rect 21140 47784 21146 47796
rect 30834 47784 30840 47796
rect 21140 47756 30840 47784
rect 21140 47744 21146 47756
rect 30834 47744 30840 47756
rect 30892 47744 30898 47796
rect 19150 47676 19156 47728
rect 19208 47716 19214 47728
rect 29822 47716 29828 47728
rect 19208 47688 29828 47716
rect 19208 47676 19214 47688
rect 29822 47676 29828 47688
rect 29880 47676 29886 47728
rect 21174 47608 21180 47660
rect 21232 47648 21238 47660
rect 26234 47648 26240 47660
rect 21232 47620 26240 47648
rect 21232 47608 21238 47620
rect 26234 47608 26240 47620
rect 26292 47608 26298 47660
rect 26418 47608 26424 47660
rect 26476 47648 26482 47660
rect 32490 47648 32496 47660
rect 26476 47620 32496 47648
rect 26476 47608 26482 47620
rect 32490 47608 32496 47620
rect 32548 47608 32554 47660
rect 37366 47648 37372 47660
rect 35866 47620 37372 47648
rect 19610 47540 19616 47592
rect 19668 47580 19674 47592
rect 35866 47580 35894 47620
rect 37366 47608 37372 47620
rect 37424 47608 37430 47660
rect 19668 47552 35894 47580
rect 19668 47540 19674 47552
rect 17218 47472 17224 47524
rect 17276 47512 17282 47524
rect 22002 47512 22008 47524
rect 17276 47484 22008 47512
rect 17276 47472 17282 47484
rect 22002 47472 22008 47484
rect 22060 47472 22066 47524
rect 26234 47472 26240 47524
rect 26292 47512 26298 47524
rect 26878 47512 26884 47524
rect 26292 47484 26884 47512
rect 26292 47472 26298 47484
rect 26878 47472 26884 47484
rect 26936 47472 26942 47524
rect 14274 47404 14280 47456
rect 14332 47444 14338 47456
rect 40770 47444 40776 47456
rect 14332 47416 40776 47444
rect 14332 47404 14338 47416
rect 40770 47404 40776 47416
rect 40828 47404 40834 47456
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 5810 47200 5816 47252
rect 5868 47240 5874 47252
rect 6457 47243 6515 47249
rect 6457 47240 6469 47243
rect 5868 47212 6469 47240
rect 5868 47200 5874 47212
rect 6457 47209 6469 47212
rect 6503 47209 6515 47243
rect 6457 47203 6515 47209
rect 13449 47243 13507 47249
rect 13449 47209 13461 47243
rect 13495 47240 13507 47243
rect 13538 47240 13544 47252
rect 13495 47212 13544 47240
rect 13495 47209 13507 47212
rect 13449 47203 13507 47209
rect 13538 47200 13544 47212
rect 13596 47200 13602 47252
rect 15105 47243 15163 47249
rect 15105 47209 15117 47243
rect 15151 47240 15163 47243
rect 15470 47240 15476 47252
rect 15151 47212 15476 47240
rect 15151 47209 15163 47212
rect 15105 47203 15163 47209
rect 15470 47200 15476 47212
rect 15528 47200 15534 47252
rect 15746 47200 15752 47252
rect 15804 47240 15810 47252
rect 19610 47240 19616 47252
rect 15804 47212 17356 47240
rect 19571 47212 19616 47240
rect 15804 47200 15810 47212
rect 4157 47175 4215 47181
rect 4157 47141 4169 47175
rect 4203 47172 4215 47175
rect 9582 47172 9588 47184
rect 4203 47144 9588 47172
rect 4203 47141 4215 47144
rect 4157 47135 4215 47141
rect 9582 47132 9588 47144
rect 9640 47132 9646 47184
rect 12161 47175 12219 47181
rect 12161 47141 12173 47175
rect 12207 47172 12219 47175
rect 17218 47172 17224 47184
rect 12207 47144 17224 47172
rect 12207 47141 12219 47144
rect 12161 47135 12219 47141
rect 17218 47132 17224 47144
rect 17276 47132 17282 47184
rect 17328 47172 17356 47212
rect 19610 47200 19616 47212
rect 19668 47200 19674 47252
rect 21174 47240 21180 47252
rect 21135 47212 21180 47240
rect 21174 47200 21180 47212
rect 21232 47200 21238 47252
rect 23198 47200 23204 47252
rect 23256 47240 23262 47252
rect 26418 47240 26424 47252
rect 23256 47212 26004 47240
rect 26379 47212 26424 47240
rect 23256 47200 23262 47212
rect 21082 47172 21088 47184
rect 17328 47144 21088 47172
rect 21082 47132 21088 47144
rect 21140 47132 21146 47184
rect 23293 47175 23351 47181
rect 23293 47172 23305 47175
rect 21376 47144 23305 47172
rect 1949 47107 2007 47113
rect 1949 47073 1961 47107
rect 1995 47104 2007 47107
rect 9122 47104 9128 47116
rect 1995 47076 9128 47104
rect 1995 47073 2007 47076
rect 1949 47067 2007 47073
rect 9122 47064 9128 47076
rect 9180 47064 9186 47116
rect 9766 47104 9772 47116
rect 9727 47076 9772 47104
rect 9766 47064 9772 47076
rect 9824 47064 9830 47116
rect 10045 47107 10103 47113
rect 10045 47073 10057 47107
rect 10091 47104 10103 47107
rect 12342 47104 12348 47116
rect 10091 47076 12348 47104
rect 10091 47073 10103 47076
rect 10045 47067 10103 47073
rect 12342 47064 12348 47076
rect 12400 47064 12406 47116
rect 12526 47064 12532 47116
rect 12584 47104 12590 47116
rect 12713 47107 12771 47113
rect 12713 47104 12725 47107
rect 12584 47076 12725 47104
rect 12584 47064 12590 47076
rect 12713 47073 12725 47076
rect 12759 47073 12771 47107
rect 12713 47067 12771 47073
rect 14182 47064 14188 47116
rect 14240 47104 14246 47116
rect 14461 47107 14519 47113
rect 14240 47076 14412 47104
rect 14240 47064 14246 47076
rect 2225 47039 2283 47045
rect 2225 47036 2237 47039
rect 1780 47008 2237 47036
rect 14 46860 20 46912
rect 72 46900 78 46912
rect 1780 46900 1808 47008
rect 2225 47005 2237 47008
rect 2271 47036 2283 47039
rect 2682 47036 2688 47048
rect 2271 47008 2688 47036
rect 2271 47005 2283 47008
rect 2225 46999 2283 47005
rect 2682 46996 2688 47008
rect 2740 46996 2746 47048
rect 3970 47036 3976 47048
rect 3931 47008 3976 47036
rect 3970 46996 3976 47008
rect 4028 47036 4034 47048
rect 4617 47039 4675 47045
rect 4617 47036 4629 47039
rect 4028 47008 4629 47036
rect 4028 46996 4034 47008
rect 4617 47005 4629 47008
rect 4663 47005 4675 47039
rect 4617 46999 4675 47005
rect 6641 47039 6699 47045
rect 6641 47005 6653 47039
rect 6687 47036 6699 47039
rect 6822 47036 6828 47048
rect 6687 47008 6828 47036
rect 6687 47005 6699 47008
rect 6641 46999 6699 47005
rect 6822 46996 6828 47008
rect 6880 46996 6886 47048
rect 7377 47039 7435 47045
rect 7377 47005 7389 47039
rect 7423 47036 7435 47039
rect 7834 47036 7840 47048
rect 7423 47008 7840 47036
rect 7423 47005 7435 47008
rect 7377 46999 7435 47005
rect 7834 46996 7840 47008
rect 7892 46996 7898 47048
rect 11606 46996 11612 47048
rect 11664 47036 11670 47048
rect 11977 47039 12035 47045
rect 11977 47036 11989 47039
rect 11664 47008 11989 47036
rect 11664 46996 11670 47008
rect 11977 47005 11989 47008
rect 12023 47005 12035 47039
rect 13265 47039 13323 47045
rect 13265 47036 13277 47039
rect 11977 46999 12035 47005
rect 12084 47008 13277 47036
rect 2777 46971 2835 46977
rect 2777 46937 2789 46971
rect 2823 46937 2835 46971
rect 2777 46931 2835 46937
rect 72 46872 1808 46900
rect 72 46860 78 46872
rect 1946 46860 1952 46912
rect 2004 46900 2010 46912
rect 2498 46900 2504 46912
rect 2004 46872 2504 46900
rect 2004 46860 2010 46872
rect 2498 46860 2504 46872
rect 2556 46900 2562 46912
rect 2792 46900 2820 46931
rect 2866 46928 2872 46980
rect 2924 46968 2930 46980
rect 2961 46971 3019 46977
rect 2961 46968 2973 46971
rect 2924 46940 2973 46968
rect 2924 46928 2930 46940
rect 2961 46937 2973 46940
rect 3007 46937 3019 46971
rect 2961 46931 3019 46937
rect 9309 46971 9367 46977
rect 9309 46937 9321 46971
rect 9355 46968 9367 46971
rect 9858 46968 9864 46980
rect 9355 46940 9864 46968
rect 9355 46937 9367 46940
rect 9309 46931 9367 46937
rect 9858 46928 9864 46940
rect 9916 46928 9922 46980
rect 10870 46928 10876 46980
rect 10928 46968 10934 46980
rect 12084 46968 12112 47008
rect 13265 47005 13277 47008
rect 13311 47005 13323 47039
rect 14274 47036 14280 47048
rect 14235 47008 14280 47036
rect 13265 46999 13323 47005
rect 14274 46996 14280 47008
rect 14332 46996 14338 47048
rect 14384 47036 14412 47076
rect 14461 47073 14473 47107
rect 14507 47104 14519 47107
rect 14734 47104 14740 47116
rect 14507 47076 14740 47104
rect 14507 47073 14519 47076
rect 14461 47067 14519 47073
rect 14734 47064 14740 47076
rect 14792 47104 14798 47116
rect 16850 47104 16856 47116
rect 14792 47076 16856 47104
rect 14792 47064 14798 47076
rect 16850 47064 16856 47076
rect 16908 47104 16914 47116
rect 17773 47107 17831 47113
rect 17773 47104 17785 47107
rect 16908 47076 17785 47104
rect 16908 47064 16914 47076
rect 17773 47073 17785 47076
rect 17819 47073 17831 47107
rect 17773 47067 17831 47073
rect 20254 47064 20260 47116
rect 20312 47104 20318 47116
rect 21376 47104 21404 47144
rect 23293 47141 23305 47144
rect 23339 47141 23351 47175
rect 23293 47135 23351 47141
rect 20312 47076 21404 47104
rect 20312 47064 20318 47076
rect 14921 47039 14979 47045
rect 14921 47036 14933 47039
rect 14384 47008 14933 47036
rect 14921 47005 14933 47008
rect 14967 47005 14979 47039
rect 15746 47036 15752 47048
rect 15707 47008 15752 47036
rect 14921 46999 14979 47005
rect 15746 46996 15752 47008
rect 15804 46996 15810 47048
rect 15841 47039 15899 47045
rect 15841 47005 15853 47039
rect 15887 47005 15899 47039
rect 17034 47036 17040 47048
rect 16995 47008 17040 47036
rect 15841 46999 15899 47005
rect 10928 46940 12112 46968
rect 12636 46940 12848 46968
rect 10928 46928 10934 46940
rect 8018 46900 8024 46912
rect 2556 46872 2820 46900
rect 7979 46872 8024 46900
rect 2556 46860 2562 46872
rect 8018 46860 8024 46872
rect 8076 46860 8082 46912
rect 10410 46860 10416 46912
rect 10468 46900 10474 46912
rect 12636 46900 12664 46940
rect 10468 46872 12664 46900
rect 12820 46900 12848 46940
rect 13924 46940 14228 46968
rect 13924 46900 13952 46940
rect 14090 46900 14096 46912
rect 12820 46872 13952 46900
rect 14051 46872 14096 46900
rect 10468 46860 10474 46872
rect 14090 46860 14096 46872
rect 14148 46860 14154 46912
rect 14200 46900 14228 46940
rect 15286 46928 15292 46980
rect 15344 46968 15350 46980
rect 15856 46968 15884 46999
rect 17034 46996 17040 47008
rect 17092 46996 17098 47048
rect 17497 47039 17555 47045
rect 17497 47005 17509 47039
rect 17543 47005 17555 47039
rect 19426 47036 19432 47048
rect 19387 47008 19432 47036
rect 17497 46999 17555 47005
rect 17402 46968 17408 46980
rect 15344 46940 15884 46968
rect 15948 46940 17408 46968
rect 15344 46928 15350 46940
rect 15948 46900 15976 46940
rect 17402 46928 17408 46940
rect 17460 46968 17466 46980
rect 17512 46968 17540 46999
rect 19426 46996 19432 47008
rect 19484 46996 19490 47048
rect 21726 46996 21732 47048
rect 21784 47036 21790 47048
rect 21913 47039 21971 47045
rect 21913 47036 21925 47039
rect 21784 47008 21925 47036
rect 21784 46996 21790 47008
rect 21913 47005 21925 47008
rect 21959 47005 21971 47039
rect 22186 47036 22192 47048
rect 22147 47008 22192 47036
rect 21913 46999 21971 47005
rect 22186 46996 22192 47008
rect 22244 46996 22250 47048
rect 23492 47045 23520 47212
rect 25976 47172 26004 47212
rect 26418 47200 26424 47212
rect 26476 47200 26482 47252
rect 34057 47243 34115 47249
rect 34057 47240 34069 47243
rect 26528 47212 34069 47240
rect 26528 47172 26556 47212
rect 34057 47209 34069 47212
rect 34103 47209 34115 47243
rect 34057 47203 34115 47209
rect 34330 47200 34336 47252
rect 34388 47240 34394 47252
rect 34388 47212 35894 47240
rect 34388 47200 34394 47212
rect 25976 47144 26556 47172
rect 27709 47175 27767 47181
rect 27709 47141 27721 47175
rect 27755 47141 27767 47175
rect 27709 47135 27767 47141
rect 27724 47104 27752 47135
rect 30834 47132 30840 47184
rect 30892 47172 30898 47184
rect 30929 47175 30987 47181
rect 30929 47172 30941 47175
rect 30892 47144 30941 47172
rect 30892 47132 30898 47144
rect 30929 47141 30941 47144
rect 30975 47141 30987 47175
rect 30929 47135 30987 47141
rect 33505 47175 33563 47181
rect 33505 47141 33517 47175
rect 33551 47172 33563 47175
rect 33870 47172 33876 47184
rect 33551 47144 33876 47172
rect 33551 47141 33563 47144
rect 33505 47135 33563 47141
rect 33870 47132 33876 47144
rect 33928 47132 33934 47184
rect 35866 47172 35894 47212
rect 37274 47200 37280 47252
rect 37332 47240 37338 47252
rect 37461 47243 37519 47249
rect 37461 47240 37473 47243
rect 37332 47212 37473 47240
rect 37332 47200 37338 47212
rect 37461 47209 37473 47212
rect 37507 47209 37519 47243
rect 37461 47203 37519 47209
rect 38289 47243 38347 47249
rect 38289 47209 38301 47243
rect 38335 47240 38347 47243
rect 38654 47240 38660 47252
rect 38335 47212 38660 47240
rect 38335 47209 38347 47212
rect 38289 47203 38347 47209
rect 38654 47200 38660 47212
rect 38712 47200 38718 47252
rect 40221 47243 40279 47249
rect 40221 47209 40233 47243
rect 40267 47240 40279 47243
rect 40586 47240 40592 47252
rect 40267 47212 40592 47240
rect 40267 47209 40279 47212
rect 40221 47203 40279 47209
rect 40586 47200 40592 47212
rect 40644 47200 40650 47252
rect 40770 47240 40776 47252
rect 40731 47212 40776 47240
rect 40770 47200 40776 47212
rect 40828 47200 40834 47252
rect 42794 47240 42800 47252
rect 42755 47212 42800 47240
rect 42794 47200 42800 47212
rect 42852 47200 42858 47252
rect 46658 47240 46664 47252
rect 46619 47212 46664 47240
rect 46658 47200 46664 47212
rect 46716 47200 46722 47252
rect 36081 47175 36139 47181
rect 36081 47172 36093 47175
rect 35866 47144 36093 47172
rect 36081 47141 36093 47144
rect 36127 47141 36139 47175
rect 36081 47135 36139 47141
rect 28350 47104 28356 47116
rect 27724 47076 28356 47104
rect 23477 47039 23535 47045
rect 23477 47005 23489 47039
rect 23523 47005 23535 47039
rect 24394 47036 24400 47048
rect 24355 47008 24400 47036
rect 23477 46999 23535 47005
rect 24394 46996 24400 47008
rect 24452 46996 24458 47048
rect 24578 47036 24584 47048
rect 24539 47008 24584 47036
rect 24578 46996 24584 47008
rect 24636 46996 24642 47048
rect 24946 46996 24952 47048
rect 25004 47036 25010 47048
rect 25041 47039 25099 47045
rect 25041 47036 25053 47039
rect 25004 47008 25053 47036
rect 25004 46996 25010 47008
rect 25041 47005 25053 47008
rect 25087 47036 25099 47039
rect 27724 47036 27752 47076
rect 28350 47064 28356 47076
rect 28408 47104 28414 47116
rect 29549 47107 29607 47113
rect 29549 47104 29561 47107
rect 28408 47076 29561 47104
rect 28408 47064 28414 47076
rect 29549 47073 29561 47076
rect 29595 47104 29607 47107
rect 36096 47104 36124 47135
rect 42426 47104 42432 47116
rect 29595 47076 32168 47104
rect 36096 47076 42432 47104
rect 29595 47073 29607 47076
rect 29549 47067 29607 47073
rect 32140 47048 32168 47076
rect 42426 47064 42432 47076
rect 42484 47104 42490 47116
rect 42484 47076 42656 47104
rect 42484 47064 42490 47076
rect 29822 47036 29828 47048
rect 25087 47008 27752 47036
rect 29783 47008 29828 47036
rect 25087 47005 25099 47008
rect 25041 46999 25099 47005
rect 29822 46996 29828 47008
rect 29880 46996 29886 47048
rect 32122 47036 32128 47048
rect 32035 47008 32128 47036
rect 32122 46996 32128 47008
rect 32180 47036 32186 47048
rect 34701 47039 34759 47045
rect 34701 47036 34713 47039
rect 32180 47008 34713 47036
rect 32180 46996 32186 47008
rect 34701 47005 34713 47008
rect 34747 47005 34759 47039
rect 36633 47039 36691 47045
rect 36633 47036 36645 47039
rect 34701 46999 34759 47005
rect 34808 47008 36645 47036
rect 20346 46968 20352 46980
rect 17460 46940 17540 46968
rect 20307 46940 20352 46968
rect 17460 46928 17466 46940
rect 20346 46928 20352 46940
rect 20404 46928 20410 46980
rect 20901 46971 20959 46977
rect 20901 46937 20913 46971
rect 20947 46968 20959 46971
rect 20990 46968 20996 46980
rect 20947 46940 20996 46968
rect 20947 46937 20959 46940
rect 20901 46931 20959 46937
rect 20990 46928 20996 46940
rect 21048 46968 21054 46980
rect 21266 46968 21272 46980
rect 21048 46940 21272 46968
rect 21048 46928 21054 46940
rect 21266 46928 21272 46940
rect 21324 46928 21330 46980
rect 22005 46971 22063 46977
rect 22005 46937 22017 46971
rect 22051 46968 22063 46971
rect 22051 46940 22085 46968
rect 22051 46937 22063 46940
rect 22005 46931 22063 46937
rect 14200 46872 15976 46900
rect 16025 46903 16083 46909
rect 16025 46869 16037 46903
rect 16071 46900 16083 46903
rect 16482 46900 16488 46912
rect 16071 46872 16488 46900
rect 16071 46869 16083 46872
rect 16025 46863 16083 46869
rect 16482 46860 16488 46872
rect 16540 46860 16546 46912
rect 20806 46860 20812 46912
rect 20864 46900 20870 46912
rect 22020 46900 22048 46931
rect 22278 46928 22284 46980
rect 22336 46968 22342 46980
rect 22373 46971 22431 46977
rect 22373 46968 22385 46971
rect 22336 46940 22385 46968
rect 22336 46928 22342 46940
rect 22373 46937 22385 46940
rect 22419 46937 22431 46971
rect 22373 46931 22431 46937
rect 24489 46971 24547 46977
rect 24489 46937 24501 46971
rect 24535 46937 24547 46971
rect 24489 46931 24547 46937
rect 25308 46971 25366 46977
rect 25308 46937 25320 46971
rect 25354 46968 25366 46971
rect 28810 46968 28816 46980
rect 25354 46940 28816 46968
rect 25354 46937 25366 46940
rect 25308 46931 25366 46937
rect 24504 46900 24532 46931
rect 28810 46928 28816 46940
rect 28868 46928 28874 46980
rect 28997 46971 29055 46977
rect 28997 46937 29009 46971
rect 29043 46968 29055 46971
rect 29178 46968 29184 46980
rect 29043 46940 29184 46968
rect 29043 46937 29055 46940
rect 28997 46931 29055 46937
rect 29178 46928 29184 46940
rect 29236 46928 29242 46980
rect 31938 46928 31944 46980
rect 31996 46968 32002 46980
rect 32370 46971 32428 46977
rect 32370 46968 32382 46971
rect 31996 46940 32382 46968
rect 31996 46928 32002 46940
rect 32370 46937 32382 46940
rect 32416 46937 32428 46971
rect 32370 46931 32428 46937
rect 32490 46928 32496 46980
rect 32548 46968 32554 46980
rect 34808 46968 34836 47008
rect 36633 47005 36645 47008
rect 36679 47036 36691 47039
rect 37277 47039 37335 47045
rect 37277 47036 37289 47039
rect 36679 47008 37289 47036
rect 36679 47005 36691 47008
rect 36633 46999 36691 47005
rect 37277 47005 37289 47008
rect 37323 47005 37335 47039
rect 37277 46999 37335 47005
rect 38654 46996 38660 47048
rect 38712 47036 38718 47048
rect 38933 47039 38991 47045
rect 38933 47036 38945 47039
rect 38712 47008 38945 47036
rect 38712 46996 38718 47008
rect 38933 47005 38945 47008
rect 38979 47005 38991 47039
rect 38933 46999 38991 47005
rect 40586 46996 40592 47048
rect 40644 47036 40650 47048
rect 42628 47045 42656 47076
rect 40865 47039 40923 47045
rect 40865 47036 40877 47039
rect 40644 47008 40877 47036
rect 40644 46996 40650 47008
rect 40865 47005 40877 47008
rect 40911 47005 40923 47039
rect 40865 46999 40923 47005
rect 42613 47039 42671 47045
rect 42613 47005 42625 47039
rect 42659 47005 42671 47039
rect 42613 46999 42671 47005
rect 46198 46996 46204 47048
rect 46256 47036 46262 47048
rect 46477 47039 46535 47045
rect 46477 47036 46489 47039
rect 46256 47008 46489 47036
rect 46256 46996 46262 47008
rect 46477 47005 46489 47008
rect 46523 47005 46535 47039
rect 46477 46999 46535 47005
rect 48041 47039 48099 47045
rect 48041 47005 48053 47039
rect 48087 47036 48099 47039
rect 48314 47036 48320 47048
rect 48087 47008 48320 47036
rect 48087 47005 48099 47008
rect 48041 46999 48099 47005
rect 48314 46996 48320 47008
rect 48372 46996 48378 47048
rect 32548 46940 34836 46968
rect 34968 46971 35026 46977
rect 32548 46928 32554 46940
rect 34968 46937 34980 46971
rect 35014 46968 35026 46971
rect 35894 46968 35900 46980
rect 35014 46940 35900 46968
rect 35014 46937 35026 46940
rect 34968 46931 35026 46937
rect 35894 46928 35900 46940
rect 35952 46928 35958 46980
rect 45373 46971 45431 46977
rect 45373 46937 45385 46971
rect 45419 46968 45431 46971
rect 45462 46968 45468 46980
rect 45419 46940 45468 46968
rect 45419 46937 45431 46940
rect 45373 46931 45431 46937
rect 45462 46928 45468 46940
rect 45520 46928 45526 46980
rect 45557 46971 45615 46977
rect 45557 46937 45569 46971
rect 45603 46937 45615 46971
rect 45557 46931 45615 46937
rect 26142 46900 26148 46912
rect 20864 46872 26148 46900
rect 20864 46860 20870 46872
rect 26142 46860 26148 46872
rect 26200 46860 26206 46912
rect 38746 46900 38752 46912
rect 38707 46872 38752 46900
rect 38746 46860 38752 46872
rect 38804 46860 38810 46912
rect 44450 46860 44456 46912
rect 44508 46900 44514 46912
rect 45186 46900 45192 46912
rect 44508 46872 45192 46900
rect 44508 46860 44514 46872
rect 45186 46860 45192 46872
rect 45244 46900 45250 46912
rect 45572 46900 45600 46931
rect 47118 46928 47124 46980
rect 47176 46968 47182 46980
rect 47857 46971 47915 46977
rect 47857 46968 47869 46971
rect 47176 46940 47869 46968
rect 47176 46928 47182 46940
rect 47857 46937 47869 46940
rect 47903 46937 47915 46971
rect 47857 46931 47915 46937
rect 45244 46872 45600 46900
rect 45244 46860 45250 46872
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 2498 46696 2504 46708
rect 2459 46668 2504 46696
rect 2498 46656 2504 46668
rect 2556 46656 2562 46708
rect 2682 46656 2688 46708
rect 2740 46696 2746 46708
rect 3053 46699 3111 46705
rect 3053 46696 3065 46699
rect 2740 46668 3065 46696
rect 2740 46656 2746 46668
rect 3053 46665 3065 46668
rect 3099 46665 3111 46699
rect 10410 46696 10416 46708
rect 10371 46668 10416 46696
rect 3053 46659 3111 46665
rect 10410 46656 10416 46668
rect 10468 46656 10474 46708
rect 19426 46696 19432 46708
rect 12820 46668 19432 46696
rect 9582 46588 9588 46640
rect 9640 46628 9646 46640
rect 11793 46631 11851 46637
rect 11793 46628 11805 46631
rect 9640 46600 11805 46628
rect 9640 46588 9646 46600
rect 11793 46597 11805 46600
rect 11839 46628 11851 46631
rect 12710 46628 12716 46640
rect 11839 46600 12716 46628
rect 11839 46597 11851 46600
rect 11793 46591 11851 46597
rect 12710 46588 12716 46600
rect 12768 46588 12774 46640
rect 1394 46560 1400 46572
rect 1355 46532 1400 46560
rect 1394 46520 1400 46532
rect 1452 46520 1458 46572
rect 12820 46560 12848 46668
rect 19426 46656 19432 46668
rect 19484 46656 19490 46708
rect 20898 46656 20904 46708
rect 20956 46696 20962 46708
rect 21085 46699 21143 46705
rect 21085 46696 21097 46699
rect 20956 46668 21097 46696
rect 20956 46656 20962 46668
rect 21085 46665 21097 46668
rect 21131 46696 21143 46699
rect 24394 46696 24400 46708
rect 21131 46668 23888 46696
rect 24355 46668 24400 46696
rect 21131 46665 21143 46668
rect 21085 46659 21143 46665
rect 12986 46628 12992 46640
rect 12947 46600 12992 46628
rect 12986 46588 12992 46600
rect 13044 46588 13050 46640
rect 14645 46631 14703 46637
rect 14645 46628 14657 46631
rect 13090 46600 14657 46628
rect 13090 46569 13118 46600
rect 14645 46597 14657 46600
rect 14691 46597 14703 46631
rect 15746 46628 15752 46640
rect 14645 46591 14703 46597
rect 15396 46600 15752 46628
rect 12406 46532 12848 46560
rect 12897 46563 12955 46569
rect 8757 46495 8815 46501
rect 8757 46461 8769 46495
rect 8803 46492 8815 46495
rect 10870 46492 10876 46504
rect 8803 46464 10876 46492
rect 8803 46461 8815 46464
rect 8757 46455 8815 46461
rect 10870 46452 10876 46464
rect 10928 46452 10934 46504
rect 9858 46424 9864 46436
rect 9771 46396 9864 46424
rect 9858 46384 9864 46396
rect 9916 46424 9922 46436
rect 10778 46424 10784 46436
rect 9916 46396 10784 46424
rect 9916 46384 9922 46396
rect 10778 46384 10784 46396
rect 10836 46384 10842 46436
rect 10965 46427 11023 46433
rect 10965 46393 10977 46427
rect 11011 46424 11023 46427
rect 12406 46424 12434 46532
rect 12897 46529 12909 46563
rect 12943 46529 12955 46563
rect 12897 46523 12955 46529
rect 13081 46563 13139 46569
rect 13081 46529 13093 46563
rect 13127 46529 13139 46563
rect 13081 46523 13139 46529
rect 11011 46396 12434 46424
rect 12912 46424 12940 46523
rect 13170 46520 13176 46572
rect 13228 46560 13234 46572
rect 13722 46560 13728 46572
rect 13228 46532 13728 46560
rect 13228 46520 13234 46532
rect 13722 46520 13728 46532
rect 13780 46520 13786 46572
rect 13814 46520 13820 46572
rect 13872 46560 13878 46572
rect 14274 46560 14280 46572
rect 13872 46532 14280 46560
rect 13872 46520 13878 46532
rect 14274 46520 14280 46532
rect 14332 46560 14338 46572
rect 14553 46563 14611 46569
rect 14553 46560 14565 46563
rect 14332 46532 14565 46560
rect 14332 46520 14338 46532
rect 14553 46529 14565 46532
rect 14599 46529 14611 46563
rect 14734 46560 14740 46572
rect 14695 46532 14740 46560
rect 14553 46523 14611 46529
rect 14734 46520 14740 46532
rect 14792 46520 14798 46572
rect 15396 46569 15424 46600
rect 15746 46588 15752 46600
rect 15804 46628 15810 46640
rect 16942 46628 16948 46640
rect 15804 46600 16948 46628
rect 15804 46588 15810 46600
rect 16942 46588 16948 46600
rect 17000 46588 17006 46640
rect 18141 46631 18199 46637
rect 18141 46597 18153 46631
rect 18187 46628 18199 46631
rect 18187 46600 18920 46628
rect 18187 46597 18199 46600
rect 18141 46591 18199 46597
rect 15381 46563 15439 46569
rect 15381 46529 15393 46563
rect 15427 46529 15439 46563
rect 16666 46560 16672 46572
rect 15381 46523 15439 46529
rect 15764 46532 16672 46560
rect 12986 46452 12992 46504
rect 13044 46492 13050 46504
rect 13633 46495 13691 46501
rect 13633 46492 13645 46495
rect 13044 46464 13645 46492
rect 13044 46452 13050 46464
rect 13633 46461 13645 46464
rect 13679 46461 13691 46495
rect 15286 46492 15292 46504
rect 13633 46455 13691 46461
rect 15120 46464 15292 46492
rect 14090 46424 14096 46436
rect 12912 46396 14096 46424
rect 11011 46393 11023 46396
rect 10965 46387 11023 46393
rect 14090 46384 14096 46396
rect 14148 46384 14154 46436
rect 1581 46359 1639 46365
rect 1581 46325 1593 46359
rect 1627 46356 1639 46359
rect 2682 46356 2688 46368
rect 1627 46328 2688 46356
rect 1627 46325 1639 46328
rect 1581 46319 1639 46325
rect 2682 46316 2688 46328
rect 2740 46316 2746 46368
rect 6822 46356 6828 46368
rect 6783 46328 6828 46356
rect 6822 46316 6828 46328
rect 6880 46316 6886 46368
rect 9306 46356 9312 46368
rect 9267 46328 9312 46356
rect 9306 46316 9312 46328
rect 9364 46316 9370 46368
rect 12434 46316 12440 46368
rect 12492 46356 12498 46368
rect 13446 46356 13452 46368
rect 12492 46328 13452 46356
rect 12492 46316 12498 46328
rect 13446 46316 13452 46328
rect 13504 46316 13510 46368
rect 14001 46359 14059 46365
rect 14001 46325 14013 46359
rect 14047 46356 14059 46359
rect 15120 46356 15148 46464
rect 15286 46452 15292 46464
rect 15344 46452 15350 46504
rect 15764 46501 15792 46532
rect 16666 46520 16672 46532
rect 16724 46560 16730 46572
rect 16853 46563 16911 46569
rect 16853 46560 16865 46563
rect 16724 46532 16865 46560
rect 16724 46520 16730 46532
rect 16853 46529 16865 46532
rect 16899 46529 16911 46563
rect 18046 46560 18052 46572
rect 18007 46532 18052 46560
rect 16853 46523 16911 46529
rect 18046 46520 18052 46532
rect 18104 46520 18110 46572
rect 18233 46563 18291 46569
rect 18233 46529 18245 46563
rect 18279 46560 18291 46563
rect 18690 46560 18696 46572
rect 18279 46532 18696 46560
rect 18279 46529 18291 46532
rect 18233 46523 18291 46529
rect 18690 46520 18696 46532
rect 18748 46520 18754 46572
rect 18892 46569 18920 46600
rect 19334 46588 19340 46640
rect 19392 46628 19398 46640
rect 19797 46631 19855 46637
rect 19797 46628 19809 46631
rect 19392 46600 19809 46628
rect 19392 46588 19398 46600
rect 19797 46597 19809 46600
rect 19843 46597 19855 46631
rect 19797 46591 19855 46597
rect 21634 46588 21640 46640
rect 21692 46628 21698 46640
rect 22094 46628 22100 46640
rect 21692 46600 22100 46628
rect 21692 46588 21698 46600
rect 18877 46563 18935 46569
rect 18877 46529 18889 46563
rect 18923 46529 18935 46563
rect 19705 46563 19763 46569
rect 19705 46560 19717 46563
rect 18877 46523 18935 46529
rect 19260 46532 19717 46560
rect 15749 46495 15807 46501
rect 15749 46461 15761 46495
rect 15795 46461 15807 46495
rect 16758 46492 16764 46504
rect 16719 46464 16764 46492
rect 15749 46455 15807 46461
rect 16758 46452 16764 46464
rect 16816 46452 16822 46504
rect 18506 46452 18512 46504
rect 18564 46492 18570 46504
rect 19260 46501 19288 46532
rect 19705 46529 19717 46532
rect 19751 46529 19763 46563
rect 19705 46523 19763 46529
rect 19981 46563 20039 46569
rect 19981 46529 19993 46563
rect 20027 46560 20039 46563
rect 20070 46560 20076 46572
rect 20027 46532 20076 46560
rect 20027 46529 20039 46532
rect 19981 46523 20039 46529
rect 20070 46520 20076 46532
rect 20128 46520 20134 46572
rect 20714 46520 20720 46572
rect 20772 46560 20778 46572
rect 20901 46563 20959 46569
rect 20901 46560 20913 46563
rect 20772 46532 20913 46560
rect 20772 46520 20778 46532
rect 20901 46529 20913 46532
rect 20947 46529 20959 46563
rect 20901 46523 20959 46529
rect 21085 46563 21143 46569
rect 21085 46529 21097 46563
rect 21131 46560 21143 46563
rect 21174 46560 21180 46572
rect 21131 46532 21180 46560
rect 21131 46529 21143 46532
rect 21085 46523 21143 46529
rect 21174 46520 21180 46532
rect 21232 46520 21238 46572
rect 21818 46520 21824 46572
rect 21876 46560 21882 46572
rect 21913 46563 21971 46569
rect 21913 46560 21925 46563
rect 21876 46532 21925 46560
rect 21876 46520 21882 46532
rect 21913 46529 21925 46532
rect 21959 46529 21971 46563
rect 22020 46546 22048 46600
rect 22094 46588 22100 46600
rect 22152 46588 22158 46640
rect 23860 46569 23888 46668
rect 24394 46656 24400 46668
rect 24452 46656 24458 46708
rect 30469 46699 30527 46705
rect 30469 46696 30481 46699
rect 27540 46668 30481 46696
rect 25958 46628 25964 46640
rect 24504 46600 25964 46628
rect 23845 46563 23903 46569
rect 21913 46523 21971 46529
rect 23845 46529 23857 46563
rect 23891 46529 23903 46563
rect 23845 46523 23903 46529
rect 24305 46563 24363 46569
rect 24305 46529 24317 46563
rect 24351 46560 24363 46563
rect 24394 46560 24400 46572
rect 24351 46532 24400 46560
rect 24351 46529 24363 46532
rect 24305 46523 24363 46529
rect 24394 46520 24400 46532
rect 24452 46520 24458 46572
rect 24504 46569 24532 46600
rect 25958 46588 25964 46600
rect 26016 46588 26022 46640
rect 24489 46563 24547 46569
rect 24489 46529 24501 46563
rect 24535 46529 24547 46563
rect 24946 46560 24952 46572
rect 24907 46532 24952 46560
rect 24489 46523 24547 46529
rect 24946 46520 24952 46532
rect 25004 46520 25010 46572
rect 25222 46569 25228 46572
rect 25216 46523 25228 46569
rect 25280 46560 25286 46572
rect 25280 46532 25316 46560
rect 25222 46520 25228 46523
rect 25280 46520 25286 46532
rect 25498 46520 25504 46572
rect 25556 46560 25562 46572
rect 25556 46532 26556 46560
rect 25556 46520 25562 46532
rect 18785 46495 18843 46501
rect 18785 46492 18797 46495
rect 18564 46464 18797 46492
rect 18564 46452 18570 46464
rect 18785 46461 18797 46464
rect 18831 46461 18843 46495
rect 18785 46455 18843 46461
rect 19245 46495 19303 46501
rect 19245 46461 19257 46495
rect 19291 46461 19303 46495
rect 22922 46492 22928 46504
rect 22835 46464 22928 46492
rect 19245 46455 19303 46461
rect 22922 46452 22928 46464
rect 22980 46492 22986 46504
rect 23566 46492 23572 46504
rect 22980 46464 23572 46492
rect 22980 46452 22986 46464
rect 23566 46452 23572 46464
rect 23624 46452 23630 46504
rect 26528 46492 26556 46532
rect 26602 46520 26608 46572
rect 26660 46560 26666 46572
rect 27249 46563 27307 46569
rect 27249 46560 27261 46563
rect 26660 46532 27261 46560
rect 26660 46520 26666 46532
rect 27249 46529 27261 46532
rect 27295 46529 27307 46563
rect 27249 46523 27307 46529
rect 26973 46495 27031 46501
rect 26973 46492 26985 46495
rect 26528 46464 26985 46492
rect 26973 46461 26985 46464
rect 27019 46492 27031 46495
rect 27540 46492 27568 46668
rect 30469 46665 30481 46668
rect 30515 46665 30527 46699
rect 30469 46659 30527 46665
rect 32858 46656 32864 46708
rect 32916 46696 32922 46708
rect 34241 46699 34299 46705
rect 34241 46696 34253 46699
rect 32916 46668 34253 46696
rect 32916 46656 32922 46668
rect 34241 46665 34253 46668
rect 34287 46665 34299 46699
rect 42426 46696 42432 46708
rect 42387 46668 42432 46696
rect 34241 46659 34299 46665
rect 42426 46656 42432 46668
rect 42484 46656 42490 46708
rect 45186 46696 45192 46708
rect 45147 46668 45192 46696
rect 45186 46656 45192 46668
rect 45244 46656 45250 46708
rect 27019 46464 27568 46492
rect 27908 46600 28488 46628
rect 27019 46461 27031 46464
rect 26973 46455 27031 46461
rect 17221 46427 17279 46433
rect 17221 46393 17233 46427
rect 17267 46424 17279 46427
rect 18230 46424 18236 46436
rect 17267 46396 18236 46424
rect 17267 46393 17279 46396
rect 17221 46387 17279 46393
rect 18230 46384 18236 46396
rect 18288 46384 18294 46436
rect 19978 46424 19984 46436
rect 19939 46396 19984 46424
rect 19978 46384 19984 46396
rect 20036 46384 20042 46436
rect 22186 46384 22192 46436
rect 22244 46424 22250 46436
rect 23385 46427 23443 46433
rect 23385 46424 23397 46427
rect 22244 46396 23397 46424
rect 22244 46384 22250 46396
rect 23385 46393 23397 46396
rect 23431 46393 23443 46427
rect 27908 46424 27936 46600
rect 28350 46560 28356 46572
rect 28311 46532 28356 46560
rect 28350 46520 28356 46532
rect 28408 46520 28414 46572
rect 28460 46560 28488 46600
rect 29288 46600 34100 46628
rect 29288 46560 29316 46600
rect 34072 46572 34100 46600
rect 34790 46588 34796 46640
rect 34848 46628 34854 46640
rect 35253 46631 35311 46637
rect 35253 46628 35265 46631
rect 34848 46600 35265 46628
rect 34848 46588 34854 46600
rect 35253 46597 35265 46600
rect 35299 46597 35311 46631
rect 35253 46591 35311 46597
rect 46937 46631 46995 46637
rect 46937 46597 46949 46631
rect 46983 46628 46995 46631
rect 47210 46628 47216 46640
rect 46983 46600 47216 46628
rect 46983 46597 46995 46600
rect 46937 46591 46995 46597
rect 47210 46588 47216 46600
rect 47268 46628 47274 46640
rect 49602 46628 49608 46640
rect 47268 46600 49608 46628
rect 47268 46588 47274 46600
rect 49602 46588 49608 46600
rect 49660 46588 49666 46640
rect 28460 46532 29316 46560
rect 30926 46520 30932 46572
rect 30984 46560 30990 46572
rect 31389 46563 31447 46569
rect 31389 46560 31401 46563
rect 30984 46532 31401 46560
rect 30984 46520 30990 46532
rect 31389 46529 31401 46532
rect 31435 46560 31447 46563
rect 31478 46560 31484 46572
rect 31435 46532 31484 46560
rect 31435 46529 31447 46532
rect 31389 46523 31447 46529
rect 31478 46520 31484 46532
rect 31536 46520 31542 46572
rect 32122 46560 32128 46572
rect 32083 46532 32128 46560
rect 32122 46520 32128 46532
rect 32180 46520 32186 46572
rect 32392 46563 32450 46569
rect 32392 46529 32404 46563
rect 32438 46560 32450 46563
rect 33962 46560 33968 46572
rect 32438 46532 33968 46560
rect 32438 46529 32450 46532
rect 32392 46523 32450 46529
rect 33962 46520 33968 46532
rect 34020 46520 34026 46572
rect 34054 46520 34060 46572
rect 34112 46560 34118 46572
rect 48041 46563 48099 46569
rect 34112 46532 34205 46560
rect 34112 46520 34118 46532
rect 48041 46529 48053 46563
rect 48087 46560 48099 46563
rect 48130 46560 48136 46572
rect 48087 46532 48136 46560
rect 48087 46529 48099 46532
rect 48041 46523 48099 46529
rect 48130 46520 48136 46532
rect 48188 46520 48194 46572
rect 27982 46452 27988 46504
rect 28040 46492 28046 46504
rect 28629 46495 28687 46501
rect 28629 46492 28641 46495
rect 28040 46464 28641 46492
rect 28040 46452 28046 46464
rect 28629 46461 28641 46464
rect 28675 46461 28687 46495
rect 28629 46455 28687 46461
rect 43254 46452 43260 46504
rect 43312 46492 43318 46504
rect 47857 46495 47915 46501
rect 47857 46492 47869 46495
rect 43312 46464 47869 46492
rect 43312 46452 43318 46464
rect 47857 46461 47869 46464
rect 47903 46461 47915 46495
rect 47857 46455 47915 46461
rect 31018 46424 31024 46436
rect 23385 46387 23443 46393
rect 26436 46396 27936 46424
rect 29288 46396 31024 46424
rect 26436 46368 26464 46396
rect 14047 46328 15148 46356
rect 14047 46325 14059 46328
rect 14001 46319 14059 46325
rect 18414 46316 18420 46368
rect 18472 46356 18478 46368
rect 20990 46356 20996 46368
rect 18472 46328 20996 46356
rect 18472 46316 18478 46328
rect 20990 46316 20996 46328
rect 21048 46316 21054 46368
rect 23753 46359 23811 46365
rect 23753 46325 23765 46359
rect 23799 46356 23811 46359
rect 24578 46356 24584 46368
rect 23799 46328 24584 46356
rect 23799 46325 23811 46328
rect 23753 46319 23811 46325
rect 24578 46316 24584 46328
rect 24636 46316 24642 46368
rect 26329 46359 26387 46365
rect 26329 46325 26341 46359
rect 26375 46356 26387 46359
rect 26418 46356 26424 46368
rect 26375 46328 26424 46356
rect 26375 46325 26387 46328
rect 26329 46319 26387 46325
rect 26418 46316 26424 46328
rect 26476 46316 26482 46368
rect 27430 46316 27436 46368
rect 27488 46356 27494 46368
rect 29288 46356 29316 46396
rect 31018 46384 31024 46396
rect 31076 46384 31082 46436
rect 34698 46384 34704 46436
rect 34756 46424 34762 46436
rect 35069 46427 35127 46433
rect 35069 46424 35081 46427
rect 34756 46396 35081 46424
rect 34756 46384 34762 46396
rect 35069 46393 35081 46396
rect 35115 46393 35127 46427
rect 46750 46424 46756 46436
rect 46711 46396 46756 46424
rect 35069 46387 35127 46393
rect 46750 46384 46756 46396
rect 46808 46384 46814 46436
rect 27488 46328 29316 46356
rect 29917 46359 29975 46365
rect 27488 46316 27494 46328
rect 29917 46325 29929 46359
rect 29963 46356 29975 46359
rect 31294 46356 31300 46368
rect 29963 46328 31300 46356
rect 29963 46325 29975 46328
rect 29917 46319 29975 46325
rect 31294 46316 31300 46328
rect 31352 46316 31358 46368
rect 31570 46356 31576 46368
rect 31531 46328 31576 46356
rect 31570 46316 31576 46328
rect 31628 46316 31634 46368
rect 33505 46359 33563 46365
rect 33505 46325 33517 46359
rect 33551 46356 33563 46359
rect 34422 46356 34428 46368
rect 33551 46328 34428 46356
rect 33551 46325 33563 46328
rect 33505 46319 33563 46325
rect 34422 46316 34428 46328
rect 34480 46316 34486 46368
rect 35894 46316 35900 46368
rect 35952 46356 35958 46368
rect 36814 46356 36820 46368
rect 35952 46328 36820 46356
rect 35952 46316 35958 46328
rect 36814 46316 36820 46328
rect 36872 46316 36878 46368
rect 46198 46356 46204 46368
rect 46159 46328 46204 46356
rect 46198 46316 46204 46328
rect 46256 46316 46262 46368
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 1394 46112 1400 46164
rect 1452 46152 1458 46164
rect 2501 46155 2559 46161
rect 2501 46152 2513 46155
rect 1452 46124 2513 46152
rect 1452 46112 1458 46124
rect 2501 46121 2513 46124
rect 2547 46121 2559 46155
rect 2501 46115 2559 46121
rect 9125 46155 9183 46161
rect 9125 46121 9137 46155
rect 9171 46152 9183 46155
rect 11606 46152 11612 46164
rect 9171 46124 11612 46152
rect 9171 46121 9183 46124
rect 9125 46115 9183 46121
rect 11606 46112 11612 46124
rect 11664 46112 11670 46164
rect 12710 46112 12716 46164
rect 12768 46152 12774 46164
rect 12897 46155 12955 46161
rect 12897 46152 12909 46155
rect 12768 46124 12909 46152
rect 12768 46112 12774 46124
rect 12897 46121 12909 46124
rect 12943 46121 12955 46155
rect 13446 46152 13452 46164
rect 13407 46124 13452 46152
rect 12897 46115 12955 46121
rect 13446 46112 13452 46124
rect 13504 46112 13510 46164
rect 14182 46152 14188 46164
rect 13556 46124 14188 46152
rect 9306 46044 9312 46096
rect 9364 46084 9370 46096
rect 13556 46084 13584 46124
rect 14182 46112 14188 46124
rect 14240 46112 14246 46164
rect 16301 46155 16359 46161
rect 16301 46121 16313 46155
rect 16347 46152 16359 46155
rect 18506 46152 18512 46164
rect 16347 46124 18512 46152
rect 16347 46121 16359 46124
rect 16301 46115 16359 46121
rect 18506 46112 18512 46124
rect 18564 46112 18570 46164
rect 18690 46152 18696 46164
rect 18651 46124 18696 46152
rect 18690 46112 18696 46124
rect 18748 46112 18754 46164
rect 19889 46155 19947 46161
rect 19889 46121 19901 46155
rect 19935 46152 19947 46155
rect 23382 46152 23388 46164
rect 19935 46124 23388 46152
rect 19935 46121 19947 46124
rect 19889 46115 19947 46121
rect 23382 46112 23388 46124
rect 23440 46112 23446 46164
rect 25958 46112 25964 46164
rect 26016 46152 26022 46164
rect 31662 46152 31668 46164
rect 26016 46124 31668 46152
rect 26016 46112 26022 46124
rect 31662 46112 31668 46124
rect 31720 46112 31726 46164
rect 33505 46155 33563 46161
rect 33505 46152 33517 46155
rect 32140 46124 33517 46152
rect 18414 46084 18420 46096
rect 9364 46056 13584 46084
rect 13648 46056 18420 46084
rect 9364 46044 9370 46056
rect 12437 46019 12495 46025
rect 12437 45985 12449 46019
rect 12483 46016 12495 46019
rect 13648 46016 13676 46056
rect 18414 46044 18420 46056
rect 18472 46044 18478 46096
rect 12483 45988 13676 46016
rect 12483 45985 12495 45988
rect 12437 45979 12495 45985
rect 13722 45976 13728 46028
rect 13780 46016 13786 46028
rect 18524 46016 18552 46112
rect 18708 46016 18736 46112
rect 21729 46087 21787 46093
rect 21729 46053 21741 46087
rect 21775 46084 21787 46087
rect 21775 46056 24716 46084
rect 21775 46053 21787 46056
rect 21729 46047 21787 46053
rect 19613 46019 19671 46025
rect 19613 46016 19625 46019
rect 13780 45988 14596 46016
rect 13780 45976 13786 45988
rect 1670 45908 1676 45960
rect 1728 45948 1734 45960
rect 1857 45951 1915 45957
rect 1857 45948 1869 45951
rect 1728 45920 1869 45948
rect 1728 45908 1734 45920
rect 1857 45917 1869 45920
rect 1903 45948 1915 45951
rect 2774 45948 2780 45960
rect 1903 45920 2780 45948
rect 1903 45917 1915 45920
rect 1857 45911 1915 45917
rect 2774 45908 2780 45920
rect 2832 45908 2838 45960
rect 14090 45948 14096 45960
rect 14051 45920 14096 45948
rect 14090 45908 14096 45920
rect 14148 45908 14154 45960
rect 14274 45948 14280 45960
rect 14235 45920 14280 45948
rect 14274 45908 14280 45920
rect 14332 45908 14338 45960
rect 14568 45957 14596 45988
rect 17696 45988 18460 46016
rect 18524 45988 18644 46016
rect 18708 45988 19625 46016
rect 14553 45951 14611 45957
rect 14553 45917 14565 45951
rect 14599 45917 14611 45951
rect 16482 45948 16488 45960
rect 16443 45920 16488 45948
rect 14553 45911 14611 45917
rect 16482 45908 16488 45920
rect 16540 45908 16546 45960
rect 16758 45948 16764 45960
rect 16719 45920 16764 45948
rect 16758 45908 16764 45920
rect 16816 45908 16822 45960
rect 17696 45957 17724 45988
rect 17681 45951 17739 45957
rect 17681 45917 17693 45951
rect 17727 45917 17739 45951
rect 17681 45911 17739 45917
rect 17865 45951 17923 45957
rect 17865 45917 17877 45951
rect 17911 45948 17923 45951
rect 18432 45948 18460 45988
rect 18616 45948 18644 45988
rect 19613 45985 19625 45988
rect 19659 45985 19671 46019
rect 20898 46016 20904 46028
rect 20859 45988 20904 46016
rect 19613 45979 19671 45985
rect 20898 45976 20904 45988
rect 20956 45976 20962 46028
rect 22002 46016 22008 46028
rect 21100 45988 22008 46016
rect 21100 45957 21128 45988
rect 22002 45976 22008 45988
rect 22060 45976 22066 46028
rect 22186 45976 22192 46028
rect 22244 46016 22250 46028
rect 22281 46019 22339 46025
rect 22281 46016 22293 46019
rect 22244 45988 22293 46016
rect 22244 45976 22250 45988
rect 22281 45985 22293 45988
rect 22327 45985 22339 46019
rect 22281 45979 22339 45985
rect 23293 46019 23351 46025
rect 23293 45985 23305 46019
rect 23339 46016 23351 46019
rect 23339 45988 24624 46016
rect 23339 45985 23351 45988
rect 23293 45979 23351 45985
rect 19705 45951 19763 45957
rect 19705 45948 19717 45951
rect 17911 45920 18368 45948
rect 18432 45920 18552 45948
rect 18616 45920 19717 45948
rect 17911 45917 17923 45920
rect 17865 45911 17923 45917
rect 13906 45840 13912 45892
rect 13964 45880 13970 45892
rect 14369 45883 14427 45889
rect 14369 45880 14381 45883
rect 13964 45852 14381 45880
rect 13964 45840 13970 45852
rect 14369 45849 14381 45852
rect 14415 45849 14427 45883
rect 14369 45843 14427 45849
rect 14458 45840 14464 45892
rect 14516 45880 14522 45892
rect 14737 45883 14795 45889
rect 14516 45852 14561 45880
rect 14516 45840 14522 45852
rect 14737 45849 14749 45883
rect 14783 45880 14795 45883
rect 16666 45880 16672 45892
rect 14783 45852 16528 45880
rect 16627 45852 16672 45880
rect 14783 45849 14795 45852
rect 14737 45843 14795 45849
rect 1946 45812 1952 45824
rect 1907 45784 1952 45812
rect 1946 45772 1952 45784
rect 2004 45772 2010 45824
rect 9677 45815 9735 45821
rect 9677 45781 9689 45815
rect 9723 45812 9735 45815
rect 10226 45812 10232 45824
rect 9723 45784 10232 45812
rect 9723 45781 9735 45784
rect 9677 45775 9735 45781
rect 10226 45772 10232 45784
rect 10284 45772 10290 45824
rect 10781 45815 10839 45821
rect 10781 45781 10793 45815
rect 10827 45812 10839 45815
rect 11241 45815 11299 45821
rect 11241 45812 11253 45815
rect 10827 45784 11253 45812
rect 10827 45781 10839 45784
rect 10781 45775 10839 45781
rect 11241 45781 11253 45784
rect 11287 45812 11299 45815
rect 11698 45812 11704 45824
rect 11287 45784 11704 45812
rect 11287 45781 11299 45784
rect 11241 45775 11299 45781
rect 11698 45772 11704 45784
rect 11756 45772 11762 45824
rect 11882 45812 11888 45824
rect 11843 45784 11888 45812
rect 11882 45772 11888 45784
rect 11940 45772 11946 45824
rect 15841 45815 15899 45821
rect 15841 45781 15853 45815
rect 15887 45812 15899 45815
rect 16022 45812 16028 45824
rect 15887 45784 16028 45812
rect 15887 45781 15899 45784
rect 15841 45775 15899 45781
rect 16022 45772 16028 45784
rect 16080 45772 16086 45824
rect 16500 45812 16528 45852
rect 16666 45840 16672 45852
rect 16724 45840 16730 45892
rect 18340 45889 18368 45920
rect 18325 45883 18383 45889
rect 18325 45849 18337 45883
rect 18371 45880 18383 45883
rect 18414 45880 18420 45892
rect 18371 45852 18420 45880
rect 18371 45849 18383 45852
rect 18325 45843 18383 45849
rect 18414 45840 18420 45852
rect 18472 45840 18478 45892
rect 18524 45889 18552 45920
rect 19705 45917 19717 45920
rect 19751 45917 19763 45951
rect 19705 45911 19763 45917
rect 21085 45951 21143 45957
rect 21085 45917 21097 45951
rect 21131 45917 21143 45951
rect 21910 45948 21916 45960
rect 21871 45920 21916 45948
rect 21085 45911 21143 45917
rect 21910 45908 21916 45920
rect 21968 45908 21974 45960
rect 22094 45908 22100 45960
rect 22152 45948 22158 45960
rect 22373 45951 22431 45957
rect 22373 45948 22385 45951
rect 22152 45920 22385 45948
rect 22152 45908 22158 45920
rect 22373 45917 22385 45920
rect 22419 45948 22431 45951
rect 23661 45951 23719 45957
rect 23661 45948 23673 45951
rect 22419 45920 23673 45948
rect 22419 45917 22431 45920
rect 22373 45911 22431 45917
rect 23661 45917 23673 45920
rect 23707 45917 23719 45951
rect 24486 45948 24492 45960
rect 24447 45920 24492 45948
rect 23661 45911 23719 45917
rect 24486 45908 24492 45920
rect 24544 45908 24550 45960
rect 18509 45883 18567 45889
rect 18509 45849 18521 45883
rect 18555 45880 18567 45883
rect 18874 45880 18880 45892
rect 18555 45852 18880 45880
rect 18555 45849 18567 45852
rect 18509 45843 18567 45849
rect 18874 45840 18880 45852
rect 18932 45880 18938 45892
rect 20162 45880 20168 45892
rect 18932 45852 20168 45880
rect 18932 45840 18938 45852
rect 20162 45840 20168 45852
rect 20220 45840 20226 45892
rect 21269 45883 21327 45889
rect 21269 45849 21281 45883
rect 21315 45880 21327 45883
rect 23566 45880 23572 45892
rect 21315 45852 23244 45880
rect 23527 45852 23572 45880
rect 21315 45849 21327 45852
rect 21269 45843 21327 45849
rect 17678 45812 17684 45824
rect 16500 45784 17684 45812
rect 17678 45772 17684 45784
rect 17736 45772 17742 45824
rect 17773 45815 17831 45821
rect 17773 45781 17785 45815
rect 17819 45812 17831 45815
rect 18046 45812 18052 45824
rect 17819 45784 18052 45812
rect 17819 45781 17831 45784
rect 17773 45775 17831 45781
rect 18046 45772 18052 45784
rect 18104 45812 18110 45824
rect 19245 45815 19303 45821
rect 19245 45812 19257 45815
rect 18104 45784 19257 45812
rect 18104 45772 18110 45784
rect 19245 45781 19257 45784
rect 19291 45781 19303 45815
rect 19245 45775 19303 45781
rect 20441 45815 20499 45821
rect 20441 45781 20453 45815
rect 20487 45812 20499 45815
rect 21450 45812 21456 45824
rect 20487 45784 21456 45812
rect 20487 45781 20499 45784
rect 20441 45775 20499 45781
rect 21450 45772 21456 45784
rect 21508 45772 21514 45824
rect 22186 45812 22192 45824
rect 22147 45784 22192 45812
rect 22186 45772 22192 45784
rect 22244 45772 22250 45824
rect 23216 45812 23244 45852
rect 23566 45840 23572 45852
rect 23624 45840 23630 45892
rect 23845 45883 23903 45889
rect 23845 45849 23857 45883
rect 23891 45880 23903 45883
rect 24397 45883 24455 45889
rect 24397 45880 24409 45883
rect 23891 45852 24409 45880
rect 23891 45849 23903 45852
rect 23845 45843 23903 45849
rect 24397 45849 24409 45852
rect 24443 45849 24455 45883
rect 24397 45843 24455 45849
rect 23477 45815 23535 45821
rect 23477 45812 23489 45815
rect 23216 45784 23489 45812
rect 23477 45781 23489 45784
rect 23523 45812 23535 45815
rect 24486 45812 24492 45824
rect 23523 45784 24492 45812
rect 23523 45781 23535 45784
rect 23477 45775 23535 45781
rect 24486 45772 24492 45784
rect 24544 45772 24550 45824
rect 24596 45812 24624 45988
rect 24688 45957 24716 46056
rect 31018 46044 31024 46096
rect 31076 46084 31082 46096
rect 31076 46056 31754 46084
rect 31076 46044 31082 46056
rect 24946 45976 24952 46028
rect 25004 46016 25010 46028
rect 25593 46019 25651 46025
rect 25593 46016 25605 46019
rect 25004 45988 25605 46016
rect 25004 45976 25010 45988
rect 25593 45985 25605 45988
rect 25639 45985 25651 46019
rect 25593 45979 25651 45985
rect 28626 45976 28632 46028
rect 28684 46016 28690 46028
rect 31389 46019 31447 46025
rect 31389 46016 31401 46019
rect 28684 45988 31401 46016
rect 28684 45976 28690 45988
rect 31389 45985 31401 45988
rect 31435 45985 31447 46019
rect 31726 46016 31754 46056
rect 32140 46016 32168 46124
rect 33505 46121 33517 46124
rect 33551 46121 33563 46155
rect 34054 46152 34060 46164
rect 34015 46124 34060 46152
rect 33505 46115 33563 46121
rect 31726 45988 32168 46016
rect 31389 45979 31447 45985
rect 24673 45951 24731 45957
rect 24673 45917 24685 45951
rect 24719 45917 24731 45951
rect 24673 45911 24731 45917
rect 24762 45908 24768 45960
rect 24820 45948 24826 45960
rect 25849 45951 25907 45957
rect 25849 45948 25861 45951
rect 24820 45920 25861 45948
rect 24820 45908 24826 45920
rect 25849 45917 25861 45920
rect 25895 45917 25907 45951
rect 25849 45911 25907 45917
rect 27062 45908 27068 45960
rect 27120 45948 27126 45960
rect 27525 45951 27583 45957
rect 27525 45948 27537 45951
rect 27120 45920 27537 45948
rect 27120 45908 27126 45920
rect 27525 45917 27537 45920
rect 27571 45948 27583 45951
rect 29086 45948 29092 45960
rect 27571 45920 29092 45948
rect 27571 45917 27583 45920
rect 27525 45911 27583 45917
rect 29086 45908 29092 45920
rect 29144 45948 29150 45960
rect 30009 45951 30067 45957
rect 30009 45948 30021 45951
rect 29144 45920 30021 45948
rect 29144 45908 29150 45920
rect 30009 45917 30021 45920
rect 30055 45917 30067 45951
rect 30282 45948 30288 45960
rect 30243 45920 30288 45948
rect 30009 45911 30067 45917
rect 30282 45908 30288 45920
rect 30340 45908 30346 45960
rect 32122 45948 32128 45960
rect 32083 45920 32128 45948
rect 32122 45908 32128 45920
rect 32180 45908 32186 45960
rect 24857 45883 24915 45889
rect 24857 45849 24869 45883
rect 24903 45880 24915 45883
rect 25130 45880 25136 45892
rect 24903 45852 25136 45880
rect 24903 45849 24915 45852
rect 24857 45843 24915 45849
rect 25130 45840 25136 45852
rect 25188 45840 25194 45892
rect 27792 45883 27850 45889
rect 27792 45849 27804 45883
rect 27838 45880 27850 45883
rect 27838 45852 30052 45880
rect 27838 45849 27850 45852
rect 27792 45843 27850 45849
rect 30024 45824 30052 45852
rect 31754 45840 31760 45892
rect 31812 45880 31818 45892
rect 32370 45883 32428 45889
rect 32370 45880 32382 45883
rect 31812 45852 32382 45880
rect 31812 45840 31818 45852
rect 32370 45849 32382 45852
rect 32416 45849 32428 45883
rect 33520 45880 33548 46115
rect 34054 46112 34060 46124
rect 34112 46112 34118 46164
rect 34790 46112 34796 46164
rect 34848 46152 34854 46164
rect 34885 46155 34943 46161
rect 34885 46152 34897 46155
rect 34848 46124 34897 46152
rect 34848 46112 34854 46124
rect 34885 46121 34897 46124
rect 34931 46121 34943 46155
rect 34885 46115 34943 46121
rect 46661 46155 46719 46161
rect 46661 46121 46673 46155
rect 46707 46152 46719 46155
rect 48130 46152 48136 46164
rect 46707 46124 48136 46152
rect 46707 46121 46719 46124
rect 46661 46115 46719 46121
rect 48130 46112 48136 46124
rect 48188 46112 48194 46164
rect 47210 46084 47216 46096
rect 47171 46056 47216 46084
rect 47210 46044 47216 46056
rect 47268 46044 47274 46096
rect 48038 45948 48044 45960
rect 47999 45920 48044 45948
rect 48038 45908 48044 45920
rect 48096 45908 48102 45960
rect 33520 45852 35894 45880
rect 32370 45843 32428 45849
rect 26142 45812 26148 45824
rect 24596 45784 26148 45812
rect 26142 45772 26148 45784
rect 26200 45772 26206 45824
rect 26970 45812 26976 45824
rect 26931 45784 26976 45812
rect 26970 45772 26976 45784
rect 27028 45772 27034 45824
rect 28534 45772 28540 45824
rect 28592 45812 28598 45824
rect 28905 45815 28963 45821
rect 28905 45812 28917 45815
rect 28592 45784 28917 45812
rect 28592 45772 28598 45784
rect 28905 45781 28917 45784
rect 28951 45781 28963 45815
rect 28905 45775 28963 45781
rect 30006 45772 30012 45824
rect 30064 45772 30070 45824
rect 35866 45812 35894 45852
rect 47026 45840 47032 45892
rect 47084 45880 47090 45892
rect 47857 45883 47915 45889
rect 47857 45880 47869 45883
rect 47084 45852 47869 45880
rect 47084 45840 47090 45852
rect 47857 45849 47869 45852
rect 47903 45849 47915 45883
rect 47857 45843 47915 45849
rect 46198 45812 46204 45824
rect 35866 45784 46204 45812
rect 46198 45772 46204 45784
rect 46256 45772 46262 45824
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 1670 45608 1676 45620
rect 1631 45580 1676 45608
rect 1670 45568 1676 45580
rect 1728 45568 1734 45620
rect 1946 45568 1952 45620
rect 2004 45608 2010 45620
rect 11146 45608 11152 45620
rect 2004 45580 11152 45608
rect 2004 45568 2010 45580
rect 11146 45568 11152 45580
rect 11204 45568 11210 45620
rect 13906 45608 13912 45620
rect 13740 45580 13912 45608
rect 9674 45540 9680 45552
rect 9635 45512 9680 45540
rect 9674 45500 9680 45512
rect 9732 45500 9738 45552
rect 11882 45540 11888 45552
rect 11843 45512 11888 45540
rect 11882 45500 11888 45512
rect 11940 45500 11946 45552
rect 12526 45540 12532 45552
rect 12487 45512 12532 45540
rect 12526 45500 12532 45512
rect 12584 45500 12590 45552
rect 13173 45543 13231 45549
rect 13173 45509 13185 45543
rect 13219 45540 13231 45543
rect 13740 45540 13768 45580
rect 13906 45568 13912 45580
rect 13964 45568 13970 45620
rect 16758 45568 16764 45620
rect 16816 45608 16822 45620
rect 16945 45611 17003 45617
rect 16945 45608 16957 45611
rect 16816 45580 16957 45608
rect 16816 45568 16822 45580
rect 16945 45577 16957 45580
rect 16991 45577 17003 45611
rect 16945 45571 17003 45577
rect 17678 45568 17684 45620
rect 17736 45608 17742 45620
rect 21726 45608 21732 45620
rect 17736 45580 21732 45608
rect 17736 45568 17742 45580
rect 14458 45540 14464 45552
rect 13219 45512 13768 45540
rect 13832 45512 14464 45540
rect 13219 45509 13231 45512
rect 13173 45503 13231 45509
rect 12544 45404 12572 45500
rect 12802 45432 12808 45484
rect 12860 45472 12866 45484
rect 12989 45475 13047 45481
rect 12989 45472 13001 45475
rect 12860 45444 13001 45472
rect 12860 45432 12866 45444
rect 12989 45441 13001 45444
rect 13035 45441 13047 45475
rect 12989 45435 13047 45441
rect 13262 45432 13268 45484
rect 13320 45472 13326 45484
rect 13832 45472 13860 45512
rect 14458 45500 14464 45512
rect 14516 45500 14522 45552
rect 15488 45512 17632 45540
rect 13320 45444 13860 45472
rect 13320 45432 13326 45444
rect 13832 45413 13860 45444
rect 13906 45432 13912 45484
rect 13964 45472 13970 45484
rect 15488 45481 15516 45512
rect 17604 45484 17632 45512
rect 15473 45475 15531 45481
rect 13964 45444 14009 45472
rect 13964 45432 13970 45444
rect 15473 45441 15485 45475
rect 15519 45441 15531 45475
rect 15473 45435 15531 45441
rect 16482 45432 16488 45484
rect 16540 45472 16546 45484
rect 16669 45475 16727 45481
rect 16669 45472 16681 45475
rect 16540 45444 16681 45472
rect 16540 45432 16546 45444
rect 16669 45441 16681 45444
rect 16715 45441 16727 45475
rect 17405 45475 17463 45481
rect 17405 45472 17417 45475
rect 16669 45435 16727 45441
rect 16776 45444 17417 45472
rect 13817 45407 13875 45413
rect 12544 45376 13768 45404
rect 12986 45336 12992 45348
rect 12947 45308 12992 45336
rect 12986 45296 12992 45308
rect 13044 45296 13050 45348
rect 13740 45336 13768 45376
rect 13817 45373 13829 45407
rect 13863 45373 13875 45407
rect 13817 45367 13875 45373
rect 14277 45407 14335 45413
rect 14277 45373 14289 45407
rect 14323 45404 14335 45407
rect 15565 45407 15623 45413
rect 15565 45404 15577 45407
rect 14323 45376 15577 45404
rect 14323 45373 14335 45376
rect 14277 45367 14335 45373
rect 15565 45373 15577 45376
rect 15611 45404 15623 45407
rect 16776 45404 16804 45444
rect 17405 45441 17417 45444
rect 17451 45441 17463 45475
rect 17586 45472 17592 45484
rect 17547 45444 17592 45472
rect 17405 45435 17463 45441
rect 17586 45432 17592 45444
rect 17644 45432 17650 45484
rect 18230 45472 18236 45484
rect 18191 45444 18236 45472
rect 18230 45432 18236 45444
rect 18288 45432 18294 45484
rect 18322 45432 18328 45484
rect 18380 45472 18386 45484
rect 18509 45475 18567 45481
rect 18380 45444 18425 45472
rect 18380 45432 18386 45444
rect 18509 45441 18521 45475
rect 18555 45472 18567 45475
rect 18598 45472 18604 45484
rect 18555 45444 18604 45472
rect 18555 45441 18567 45444
rect 18509 45435 18567 45441
rect 18598 45432 18604 45444
rect 18656 45432 18662 45484
rect 15611 45376 16804 45404
rect 16945 45407 17003 45413
rect 15611 45373 15623 45376
rect 15565 45367 15623 45373
rect 16945 45373 16957 45407
rect 16991 45404 17003 45407
rect 17497 45407 17555 45413
rect 17497 45404 17509 45407
rect 16991 45376 17509 45404
rect 16991 45373 17003 45376
rect 16945 45367 17003 45373
rect 17497 45373 17509 45376
rect 17543 45373 17555 45407
rect 17497 45367 17555 45373
rect 18414 45364 18420 45416
rect 18472 45404 18478 45416
rect 18969 45407 19027 45413
rect 18969 45404 18981 45407
rect 18472 45376 18981 45404
rect 18472 45364 18478 45376
rect 18969 45373 18981 45376
rect 19015 45373 19027 45407
rect 19261 45404 19289 45580
rect 21726 45568 21732 45580
rect 21784 45568 21790 45620
rect 22094 45568 22100 45620
rect 22152 45608 22158 45620
rect 26142 45608 26148 45620
rect 22152 45580 23152 45608
rect 26103 45580 26148 45608
rect 22152 45568 22158 45580
rect 20714 45500 20720 45552
rect 20772 45540 20778 45552
rect 20901 45543 20959 45549
rect 20901 45540 20913 45543
rect 20772 45512 20913 45540
rect 20772 45500 20778 45512
rect 20901 45509 20913 45512
rect 20947 45509 20959 45543
rect 20901 45503 20959 45509
rect 20990 45500 20996 45552
rect 21048 45540 21054 45552
rect 21634 45540 21640 45552
rect 21048 45512 21640 45540
rect 21048 45500 21054 45512
rect 21634 45500 21640 45512
rect 21692 45540 21698 45552
rect 21959 45543 22017 45549
rect 21959 45540 21971 45543
rect 21692 45512 21971 45540
rect 21692 45500 21698 45512
rect 21959 45509 21971 45512
rect 22005 45509 22017 45543
rect 21959 45503 22017 45509
rect 22186 45500 22192 45552
rect 22244 45540 22250 45552
rect 22922 45540 22928 45552
rect 22244 45512 22928 45540
rect 22244 45500 22250 45512
rect 22922 45500 22928 45512
rect 22980 45500 22986 45552
rect 19337 45475 19395 45481
rect 19337 45441 19349 45475
rect 19383 45472 19395 45475
rect 20806 45472 20812 45484
rect 19383 45444 20812 45472
rect 19383 45441 19395 45444
rect 19337 45435 19395 45441
rect 20806 45432 20812 45444
rect 20864 45432 20870 45484
rect 21082 45472 21088 45484
rect 21043 45444 21088 45472
rect 21082 45432 21088 45444
rect 21140 45432 21146 45484
rect 21269 45475 21327 45481
rect 21269 45441 21281 45475
rect 21315 45472 21327 45475
rect 22097 45475 22155 45481
rect 22097 45472 22109 45475
rect 21315 45444 22109 45472
rect 21315 45441 21327 45444
rect 21269 45435 21327 45441
rect 22020 45416 22048 45444
rect 22097 45441 22109 45444
rect 22143 45441 22155 45475
rect 22097 45435 22155 45441
rect 22278 45432 22284 45484
rect 22336 45472 22342 45484
rect 23124 45481 23152 45580
rect 26142 45568 26148 45580
rect 26200 45568 26206 45620
rect 26786 45568 26792 45620
rect 26844 45608 26850 45620
rect 28626 45608 28632 45620
rect 26844 45580 28632 45608
rect 26844 45568 26850 45580
rect 28626 45568 28632 45580
rect 28684 45568 28690 45620
rect 28994 45568 29000 45620
rect 29052 45608 29058 45620
rect 30374 45608 30380 45620
rect 29052 45580 30380 45608
rect 29052 45568 29058 45580
rect 30374 45568 30380 45580
rect 30432 45608 30438 45620
rect 31478 45608 31484 45620
rect 30432 45580 30972 45608
rect 31439 45580 31484 45608
rect 30432 45568 30438 45580
rect 23198 45500 23204 45552
rect 23256 45540 23262 45552
rect 30944 45549 30972 45580
rect 31478 45568 31484 45580
rect 31536 45568 31542 45620
rect 31662 45568 31668 45620
rect 31720 45608 31726 45620
rect 38746 45608 38752 45620
rect 31720 45580 38752 45608
rect 31720 45568 31726 45580
rect 38746 45568 38752 45580
rect 38804 45568 38810 45620
rect 48038 45608 48044 45620
rect 47999 45580 48044 45608
rect 48038 45568 48044 45580
rect 48096 45568 48102 45620
rect 30929 45543 30987 45549
rect 23256 45512 25544 45540
rect 23256 45500 23262 45512
rect 23109 45475 23167 45481
rect 22336 45444 22381 45472
rect 22336 45432 22342 45444
rect 23109 45441 23121 45475
rect 23155 45441 23167 45475
rect 23109 45435 23167 45441
rect 23566 45432 23572 45484
rect 23624 45472 23630 45484
rect 24121 45475 24179 45481
rect 24121 45472 24133 45475
rect 23624 45444 24133 45472
rect 23624 45432 23630 45444
rect 24121 45441 24133 45444
rect 24167 45441 24179 45475
rect 24121 45435 24179 45441
rect 24486 45432 24492 45484
rect 24544 45472 24550 45484
rect 25239 45475 25297 45481
rect 25239 45472 25251 45475
rect 24544 45444 25251 45472
rect 24544 45432 24550 45444
rect 25239 45441 25251 45444
rect 25285 45441 25297 45475
rect 25239 45435 25297 45441
rect 19429 45407 19487 45413
rect 19429 45404 19441 45407
rect 19261 45376 19441 45404
rect 18969 45367 19027 45373
rect 19429 45373 19441 45376
rect 19475 45373 19487 45407
rect 19429 45367 19487 45373
rect 20990 45364 20996 45416
rect 21048 45404 21054 45416
rect 21818 45404 21824 45416
rect 21048 45376 21824 45404
rect 21048 45364 21054 45376
rect 21818 45364 21824 45376
rect 21876 45364 21882 45416
rect 22002 45364 22008 45416
rect 22060 45364 22066 45416
rect 22465 45407 22523 45413
rect 22465 45373 22477 45407
rect 22511 45404 22523 45407
rect 23017 45407 23075 45413
rect 23017 45404 23029 45407
rect 22511 45376 23029 45404
rect 22511 45373 22523 45376
rect 22465 45367 22523 45373
rect 23017 45373 23029 45376
rect 23063 45373 23075 45407
rect 24026 45404 24032 45416
rect 23987 45376 24032 45404
rect 23017 45367 23075 45373
rect 24026 45364 24032 45376
rect 24084 45364 24090 45416
rect 24394 45364 24400 45416
rect 24452 45404 24458 45416
rect 25038 45404 25044 45416
rect 24452 45376 25044 45404
rect 24452 45364 24458 45376
rect 25038 45364 25044 45376
rect 25096 45404 25102 45416
rect 25409 45407 25467 45413
rect 25096 45376 25268 45404
rect 25096 45364 25102 45376
rect 14458 45336 14464 45348
rect 13740 45308 14464 45336
rect 14458 45296 14464 45308
rect 14516 45296 14522 45348
rect 15841 45339 15899 45345
rect 15841 45305 15853 45339
rect 15887 45336 15899 45339
rect 16574 45336 16580 45348
rect 15887 45308 16580 45336
rect 15887 45305 15899 45308
rect 15841 45299 15899 45305
rect 16574 45296 16580 45308
rect 16632 45336 16638 45348
rect 16761 45339 16819 45345
rect 16761 45336 16773 45339
rect 16632 45308 16773 45336
rect 16632 45296 16638 45308
rect 16761 45305 16773 45308
rect 16807 45305 16819 45339
rect 16761 45299 16819 45305
rect 18509 45339 18567 45345
rect 18509 45305 18521 45339
rect 18555 45336 18567 45339
rect 19150 45336 19156 45348
rect 18555 45308 19156 45336
rect 18555 45305 18567 45308
rect 18509 45299 18567 45305
rect 19150 45296 19156 45308
rect 19208 45296 19214 45348
rect 19334 45296 19340 45348
rect 19392 45336 19398 45348
rect 19392 45308 20852 45336
rect 19392 45296 19398 45308
rect 10410 45268 10416 45280
rect 10323 45240 10416 45268
rect 10410 45228 10416 45240
rect 10468 45268 10474 45280
rect 10965 45271 11023 45277
rect 10965 45268 10977 45271
rect 10468 45240 10977 45268
rect 10468 45228 10474 45240
rect 10965 45237 10977 45240
rect 11011 45268 11023 45271
rect 12158 45268 12164 45280
rect 11011 45240 12164 45268
rect 11011 45237 11023 45240
rect 10965 45231 11023 45237
rect 12158 45228 12164 45240
rect 12216 45228 12222 45280
rect 12618 45228 12624 45280
rect 12676 45268 12682 45280
rect 14737 45271 14795 45277
rect 14737 45268 14749 45271
rect 12676 45240 14749 45268
rect 12676 45228 12682 45240
rect 14737 45237 14749 45240
rect 14783 45237 14795 45271
rect 14737 45231 14795 45237
rect 16022 45228 16028 45280
rect 16080 45268 16086 45280
rect 20438 45268 20444 45280
rect 16080 45240 20444 45268
rect 16080 45228 16086 45240
rect 20438 45228 20444 45240
rect 20496 45228 20502 45280
rect 20824 45268 20852 45308
rect 21174 45296 21180 45348
rect 21232 45336 21238 45348
rect 24412 45336 24440 45364
rect 21232 45308 24440 45336
rect 24489 45339 24547 45345
rect 21232 45296 21238 45308
rect 24489 45305 24501 45339
rect 24535 45336 24547 45339
rect 24854 45336 24860 45348
rect 24535 45308 24860 45336
rect 24535 45305 24547 45308
rect 24489 45299 24547 45305
rect 24854 45296 24860 45308
rect 24912 45296 24918 45348
rect 23198 45268 23204 45280
rect 20824 45240 23204 45268
rect 23198 45228 23204 45240
rect 23256 45228 23262 45280
rect 23474 45268 23480 45280
rect 23435 45240 23480 45268
rect 23474 45228 23480 45240
rect 23532 45228 23538 45280
rect 23934 45228 23940 45280
rect 23992 45268 23998 45280
rect 25041 45271 25099 45277
rect 25041 45268 25053 45271
rect 23992 45240 25053 45268
rect 23992 45228 23998 45240
rect 25041 45237 25053 45240
rect 25087 45237 25099 45271
rect 25240 45268 25268 45376
rect 25409 45373 25421 45407
rect 25455 45373 25467 45407
rect 25516 45404 25544 45512
rect 30929 45509 30941 45543
rect 30975 45509 30987 45543
rect 30929 45503 30987 45509
rect 32140 45512 33548 45540
rect 32140 45484 32168 45512
rect 25958 45472 25964 45484
rect 25919 45444 25964 45472
rect 25958 45432 25964 45444
rect 26016 45432 26022 45484
rect 26234 45472 26240 45484
rect 26195 45444 26240 45472
rect 26234 45432 26240 45444
rect 26292 45432 26298 45484
rect 26970 45432 26976 45484
rect 27028 45472 27034 45484
rect 27157 45475 27215 45481
rect 27157 45472 27169 45475
rect 27028 45444 27169 45472
rect 27028 45432 27034 45444
rect 27157 45441 27169 45444
rect 27203 45441 27215 45475
rect 29638 45472 29644 45484
rect 29599 45444 29644 45472
rect 27157 45435 27215 45441
rect 29638 45432 29644 45444
rect 29696 45432 29702 45484
rect 29917 45475 29975 45481
rect 29917 45441 29929 45475
rect 29963 45472 29975 45475
rect 32122 45472 32128 45484
rect 29963 45444 32128 45472
rect 29963 45441 29975 45444
rect 29917 45435 29975 45441
rect 32122 45432 32128 45444
rect 32180 45432 32186 45484
rect 33226 45472 33232 45484
rect 33284 45481 33290 45484
rect 33520 45481 33548 45512
rect 33870 45500 33876 45552
rect 33928 45540 33934 45552
rect 33928 45512 34836 45540
rect 33928 45500 33934 45512
rect 33196 45444 33232 45472
rect 33226 45432 33232 45444
rect 33284 45435 33296 45481
rect 33505 45475 33563 45481
rect 33505 45441 33517 45475
rect 33551 45441 33563 45475
rect 34606 45472 34612 45484
rect 34567 45444 34612 45472
rect 33505 45435 33563 45441
rect 33284 45432 33290 45435
rect 34606 45432 34612 45444
rect 34664 45432 34670 45484
rect 34808 45481 34836 45512
rect 34793 45475 34851 45481
rect 34793 45441 34805 45475
rect 34839 45472 34851 45475
rect 35253 45475 35311 45481
rect 35253 45472 35265 45475
rect 34839 45444 35265 45472
rect 34839 45441 34851 45444
rect 34793 45435 34851 45441
rect 35253 45441 35265 45444
rect 35299 45441 35311 45475
rect 35253 45435 35311 45441
rect 31018 45404 31024 45416
rect 25516 45376 31024 45404
rect 25409 45367 25467 45373
rect 25424 45336 25452 45367
rect 31018 45364 31024 45376
rect 31076 45364 31082 45416
rect 34701 45407 34759 45413
rect 34701 45373 34713 45407
rect 34747 45404 34759 45407
rect 35526 45404 35532 45416
rect 34747 45376 35532 45404
rect 34747 45373 34759 45376
rect 34701 45367 34759 45373
rect 35526 45364 35532 45376
rect 35584 45364 35590 45416
rect 25961 45339 26019 45345
rect 25961 45336 25973 45339
rect 25424 45308 25973 45336
rect 25961 45305 25973 45308
rect 26007 45305 26019 45339
rect 25961 45299 26019 45305
rect 27154 45296 27160 45348
rect 27212 45336 27218 45348
rect 27341 45339 27399 45345
rect 27341 45336 27353 45339
rect 27212 45308 27353 45336
rect 27212 45296 27218 45308
rect 27341 45305 27353 45308
rect 27387 45305 27399 45339
rect 27341 45299 27399 45305
rect 27448 45308 28488 45336
rect 27448 45268 27476 45308
rect 28350 45268 28356 45280
rect 25240 45240 27476 45268
rect 28311 45240 28356 45268
rect 25041 45231 25099 45237
rect 28350 45228 28356 45240
rect 28408 45228 28414 45280
rect 28460 45268 28488 45308
rect 32030 45296 32036 45348
rect 32088 45336 32094 45348
rect 32125 45339 32183 45345
rect 32125 45336 32137 45339
rect 32088 45308 32137 45336
rect 32088 45296 32094 45308
rect 32125 45305 32137 45308
rect 32171 45305 32183 45339
rect 43254 45336 43260 45348
rect 32125 45299 32183 45305
rect 33520 45308 43260 45336
rect 30469 45271 30527 45277
rect 30469 45268 30481 45271
rect 28460 45240 30481 45268
rect 30469 45237 30481 45240
rect 30515 45268 30527 45271
rect 33520 45268 33548 45308
rect 43254 45296 43260 45308
rect 43312 45296 43318 45348
rect 30515 45240 33548 45268
rect 30515 45237 30527 45240
rect 30469 45231 30527 45237
rect 33870 45228 33876 45280
rect 33928 45268 33934 45280
rect 34054 45268 34060 45280
rect 33928 45240 34060 45268
rect 33928 45228 33934 45240
rect 34054 45228 34060 45240
rect 34112 45228 34118 45280
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 12989 45067 13047 45073
rect 12989 45033 13001 45067
rect 13035 45064 13047 45067
rect 13262 45064 13268 45076
rect 13035 45036 13268 45064
rect 13035 45033 13047 45036
rect 12989 45027 13047 45033
rect 13262 45024 13268 45036
rect 13320 45024 13326 45076
rect 14274 45024 14280 45076
rect 14332 45064 14338 45076
rect 14737 45067 14795 45073
rect 14737 45064 14749 45067
rect 14332 45036 14749 45064
rect 14332 45024 14338 45036
rect 14737 45033 14749 45036
rect 14783 45033 14795 45067
rect 14737 45027 14795 45033
rect 16025 45067 16083 45073
rect 16025 45033 16037 45067
rect 16071 45064 16083 45067
rect 17034 45064 17040 45076
rect 16071 45036 17040 45064
rect 16071 45033 16083 45036
rect 16025 45027 16083 45033
rect 17034 45024 17040 45036
rect 17092 45064 17098 45076
rect 17497 45067 17555 45073
rect 17497 45064 17509 45067
rect 17092 45036 17509 45064
rect 17092 45024 17098 45036
rect 17497 45033 17509 45036
rect 17543 45064 17555 45067
rect 20530 45064 20536 45076
rect 17543 45036 20536 45064
rect 17543 45033 17555 45036
rect 17497 45027 17555 45033
rect 20530 45024 20536 45036
rect 20588 45064 20594 45076
rect 21634 45064 21640 45076
rect 20588 45036 21640 45064
rect 20588 45024 20594 45036
rect 21634 45024 21640 45036
rect 21692 45024 21698 45076
rect 22094 45024 22100 45076
rect 22152 45064 22158 45076
rect 22649 45067 22707 45073
rect 22152 45036 22197 45064
rect 22152 45024 22158 45036
rect 22649 45033 22661 45067
rect 22695 45064 22707 45067
rect 24026 45064 24032 45076
rect 22695 45036 24032 45064
rect 22695 45033 22707 45036
rect 22649 45027 22707 45033
rect 24026 45024 24032 45036
rect 24084 45024 24090 45076
rect 24578 45024 24584 45076
rect 24636 45064 24642 45076
rect 24765 45067 24823 45073
rect 24765 45064 24777 45067
rect 24636 45036 24777 45064
rect 24636 45024 24642 45036
rect 24765 45033 24777 45036
rect 24811 45064 24823 45067
rect 25958 45064 25964 45076
rect 24811 45036 25964 45064
rect 24811 45033 24823 45036
rect 24765 45027 24823 45033
rect 25958 45024 25964 45036
rect 26016 45024 26022 45076
rect 26237 45067 26295 45073
rect 26237 45033 26249 45067
rect 26283 45064 26295 45067
rect 28445 45067 28503 45073
rect 26283 45036 28120 45064
rect 26283 45033 26295 45036
rect 26237 45027 26295 45033
rect 18049 44999 18107 45005
rect 18049 44996 18061 44999
rect 6886 44968 18061 44996
rect 6886 44804 6914 44968
rect 18049 44965 18061 44968
rect 18095 44996 18107 44999
rect 19981 44999 20039 45005
rect 19981 44996 19993 44999
rect 18095 44968 19993 44996
rect 18095 44965 18107 44968
rect 18049 44959 18107 44965
rect 19981 44965 19993 44968
rect 20027 44996 20039 44999
rect 22186 44996 22192 45008
rect 20027 44968 22192 44996
rect 20027 44965 20039 44968
rect 19981 44959 20039 44965
rect 22186 44956 22192 44968
rect 22244 44956 22250 45008
rect 23474 44956 23480 45008
rect 23532 44996 23538 45008
rect 23532 44968 25728 44996
rect 23532 44956 23538 44968
rect 13998 44888 14004 44940
rect 14056 44928 14062 44940
rect 16574 44928 16580 44940
rect 14056 44900 14320 44928
rect 16535 44900 16580 44928
rect 14056 44888 14062 44900
rect 10226 44820 10232 44872
rect 10284 44860 10290 44872
rect 10597 44863 10655 44869
rect 10597 44860 10609 44863
rect 10284 44832 10609 44860
rect 10284 44820 10290 44832
rect 10597 44829 10609 44832
rect 10643 44860 10655 44863
rect 12802 44860 12808 44872
rect 10643 44832 12572 44860
rect 12763 44832 12808 44860
rect 10643 44829 10655 44832
rect 10597 44823 10655 44829
rect 6822 44752 6828 44804
rect 6880 44764 6914 44804
rect 6880 44752 6886 44764
rect 10870 44752 10876 44804
rect 10928 44792 10934 44804
rect 11701 44795 11759 44801
rect 11701 44792 11713 44795
rect 10928 44764 11713 44792
rect 10928 44752 10934 44764
rect 11701 44761 11713 44764
rect 11747 44761 11759 44795
rect 11701 44755 11759 44761
rect 12345 44795 12403 44801
rect 12345 44761 12357 44795
rect 12391 44792 12403 44795
rect 12434 44792 12440 44804
rect 12391 44764 12440 44792
rect 12391 44761 12403 44764
rect 12345 44755 12403 44761
rect 12434 44752 12440 44764
rect 12492 44752 12498 44804
rect 12544 44792 12572 44832
rect 12802 44820 12808 44832
rect 12860 44820 12866 44872
rect 12989 44863 13047 44869
rect 12989 44829 13001 44863
rect 13035 44860 13047 44863
rect 13262 44860 13268 44872
rect 13035 44832 13268 44860
rect 13035 44829 13047 44832
rect 12989 44823 13047 44829
rect 13262 44820 13268 44832
rect 13320 44820 13326 44872
rect 13354 44820 13360 44872
rect 13412 44860 13418 44872
rect 14292 44869 14320 44900
rect 16574 44888 16580 44900
rect 16632 44888 16638 44940
rect 17034 44928 17040 44940
rect 16995 44900 17040 44928
rect 17034 44888 17040 44900
rect 17092 44888 17098 44940
rect 20438 44888 20444 44940
rect 20496 44928 20502 44940
rect 21634 44928 21640 44940
rect 20496 44900 21128 44928
rect 21595 44900 21640 44928
rect 20496 44888 20502 44900
rect 14117 44863 14175 44869
rect 14117 44860 14129 44863
rect 13412 44850 13952 44860
rect 14108 44850 14129 44860
rect 13412 44832 14129 44850
rect 13412 44820 13418 44832
rect 13924 44829 14129 44832
rect 14163 44829 14175 44863
rect 13924 44823 14175 44829
rect 14277 44863 14335 44869
rect 14277 44829 14289 44863
rect 14323 44829 14335 44863
rect 14277 44823 14335 44829
rect 14388 44860 14446 44866
rect 14388 44826 14400 44860
rect 14434 44826 14446 44860
rect 13924 44822 14136 44823
rect 14388 44820 14446 44826
rect 14507 44863 14565 44869
rect 14507 44829 14519 44863
rect 14553 44860 14565 44863
rect 14734 44860 14740 44872
rect 14553 44832 14740 44860
rect 14553 44829 14565 44832
rect 14507 44823 14565 44829
rect 14734 44820 14740 44832
rect 14792 44820 14798 44872
rect 15102 44820 15108 44872
rect 15160 44860 15166 44872
rect 15289 44863 15347 44869
rect 15289 44860 15301 44863
rect 15160 44832 15301 44860
rect 15160 44820 15166 44832
rect 15289 44829 15301 44832
rect 15335 44829 15347 44863
rect 15470 44860 15476 44872
rect 15431 44832 15476 44860
rect 15289 44823 15347 44829
rect 15470 44820 15476 44832
rect 15528 44820 15534 44872
rect 16482 44860 16488 44872
rect 16395 44832 16488 44860
rect 13814 44792 13820 44804
rect 12544 44764 13820 44792
rect 13814 44752 13820 44764
rect 13872 44752 13878 44804
rect 14403 44792 14431 44820
rect 14642 44792 14648 44804
rect 14403 44764 14648 44792
rect 14642 44752 14648 44764
rect 14700 44752 14706 44804
rect 15381 44795 15439 44801
rect 15381 44761 15393 44795
rect 15427 44792 15439 44795
rect 16408 44792 16436 44832
rect 16482 44820 16488 44832
rect 16540 44860 16546 44872
rect 16662 44863 16720 44869
rect 16662 44860 16674 44863
rect 16540 44832 16674 44860
rect 16540 44820 16546 44832
rect 16662 44829 16674 44832
rect 16708 44829 16720 44863
rect 19242 44860 19248 44872
rect 19203 44832 19248 44860
rect 16662 44823 16720 44829
rect 19242 44820 19248 44832
rect 19300 44820 19306 44872
rect 19429 44863 19487 44869
rect 19429 44829 19441 44863
rect 19475 44829 19487 44863
rect 20530 44860 20536 44872
rect 20491 44832 20536 44860
rect 19429 44823 19487 44829
rect 15427 44764 16436 44792
rect 19444 44792 19472 44823
rect 20530 44820 20536 44832
rect 20588 44820 20594 44872
rect 20732 44869 20760 44900
rect 20717 44863 20775 44869
rect 20717 44829 20729 44863
rect 20763 44829 20775 44863
rect 20898 44860 20904 44872
rect 20859 44832 20904 44860
rect 20717 44823 20775 44829
rect 20898 44820 20904 44832
rect 20956 44820 20962 44872
rect 21100 44860 21128 44900
rect 21634 44888 21640 44900
rect 21692 44888 21698 44940
rect 22002 44888 22008 44940
rect 22060 44928 22066 44940
rect 25700 44928 25728 44968
rect 25774 44956 25780 45008
rect 25832 44996 25838 45008
rect 26252 44996 26280 45027
rect 25832 44968 26280 44996
rect 25832 44956 25838 44968
rect 27062 44928 27068 44940
rect 22060 44900 22784 44928
rect 25700 44900 26924 44928
rect 27023 44900 27068 44928
rect 22060 44888 22066 44900
rect 21726 44860 21732 44872
rect 21100 44832 21732 44860
rect 21726 44820 21732 44832
rect 21784 44820 21790 44872
rect 22278 44820 22284 44872
rect 22336 44860 22342 44872
rect 22756 44869 22784 44900
rect 22557 44863 22615 44869
rect 22557 44860 22569 44863
rect 22336 44832 22569 44860
rect 22336 44820 22342 44832
rect 22557 44829 22569 44832
rect 22603 44829 22615 44863
rect 22557 44823 22615 44829
rect 22741 44863 22799 44869
rect 22741 44829 22753 44863
rect 22787 44829 22799 44863
rect 22741 44823 22799 44829
rect 24949 44863 25007 44869
rect 24949 44829 24961 44863
rect 24995 44829 25007 44863
rect 24949 44823 25007 44829
rect 20809 44795 20867 44801
rect 19444 44764 20760 44792
rect 15427 44761 15439 44764
rect 15381 44755 15439 44761
rect 20732 44736 20760 44764
rect 20809 44761 20821 44795
rect 20855 44761 20867 44795
rect 20809 44755 20867 44761
rect 9858 44684 9864 44736
rect 9916 44724 9922 44736
rect 10045 44727 10103 44733
rect 10045 44724 10057 44727
rect 9916 44696 10057 44724
rect 9916 44684 9922 44696
rect 10045 44693 10057 44696
rect 10091 44693 10103 44727
rect 11238 44724 11244 44736
rect 11199 44696 11244 44724
rect 10045 44687 10103 44693
rect 11238 44684 11244 44696
rect 11296 44684 11302 44736
rect 13541 44727 13599 44733
rect 13541 44693 13553 44727
rect 13587 44724 13599 44727
rect 16022 44724 16028 44736
rect 13587 44696 16028 44724
rect 13587 44693 13599 44696
rect 13541 44687 13599 44693
rect 16022 44684 16028 44696
rect 16080 44684 16086 44736
rect 17954 44684 17960 44736
rect 18012 44724 18018 44736
rect 18601 44727 18659 44733
rect 18601 44724 18613 44727
rect 18012 44696 18613 44724
rect 18012 44684 18018 44696
rect 18601 44693 18613 44696
rect 18647 44724 18659 44727
rect 19150 44724 19156 44736
rect 18647 44696 19156 44724
rect 18647 44693 18659 44696
rect 18601 44687 18659 44693
rect 19150 44684 19156 44696
rect 19208 44684 19214 44736
rect 19334 44724 19340 44736
rect 19295 44696 19340 44724
rect 19334 44684 19340 44696
rect 19392 44684 19398 44736
rect 20714 44684 20720 44736
rect 20772 44684 20778 44736
rect 20824 44724 20852 44755
rect 23198 44752 23204 44804
rect 23256 44792 23262 44804
rect 24964 44792 24992 44823
rect 25038 44820 25044 44872
rect 25096 44860 25102 44872
rect 26050 44860 26056 44872
rect 25096 44832 25141 44860
rect 25240 44832 26056 44860
rect 25096 44820 25102 44832
rect 25240 44792 25268 44832
rect 26050 44820 26056 44832
rect 26108 44820 26114 44872
rect 26896 44860 26924 44900
rect 27062 44888 27068 44900
rect 27120 44888 27126 44940
rect 28092 44928 28120 45036
rect 28445 45033 28457 45067
rect 28491 45064 28503 45067
rect 30926 45064 30932 45076
rect 28491 45036 30932 45064
rect 28491 45033 28503 45036
rect 28445 45027 28503 45033
rect 30926 45024 30932 45036
rect 30984 45024 30990 45076
rect 31018 45024 31024 45076
rect 31076 45064 31082 45076
rect 47946 45064 47952 45076
rect 31076 45036 47952 45064
rect 31076 45024 31082 45036
rect 47946 45024 47952 45036
rect 48004 45024 48010 45076
rect 48130 45064 48136 45076
rect 48091 45036 48136 45064
rect 48130 45024 48136 45036
rect 48188 45024 48194 45076
rect 31205 44931 31263 44937
rect 28092 44900 31156 44928
rect 26896 44832 28212 44860
rect 23256 44764 24900 44792
rect 24964 44764 25268 44792
rect 25685 44795 25743 44801
rect 23256 44752 23262 44764
rect 20990 44724 20996 44736
rect 20824 44696 20996 44724
rect 20990 44684 20996 44696
rect 21048 44684 21054 44736
rect 21085 44727 21143 44733
rect 21085 44693 21097 44727
rect 21131 44724 21143 44727
rect 22002 44724 22008 44736
rect 21131 44696 22008 44724
rect 21131 44693 21143 44696
rect 21085 44687 21143 44693
rect 22002 44684 22008 44696
rect 22060 44684 22066 44736
rect 23293 44727 23351 44733
rect 23293 44693 23305 44727
rect 23339 44724 23351 44727
rect 23474 44724 23480 44736
rect 23339 44696 23480 44724
rect 23339 44693 23351 44696
rect 23293 44687 23351 44693
rect 23474 44684 23480 44696
rect 23532 44684 23538 44736
rect 23750 44724 23756 44736
rect 23711 44696 23756 44724
rect 23750 44684 23756 44696
rect 23808 44684 23814 44736
rect 24872 44724 24900 44764
rect 25685 44761 25697 44795
rect 25731 44792 25743 44795
rect 27332 44795 27390 44801
rect 25731 44764 27200 44792
rect 25731 44761 25743 44764
rect 25685 44755 25743 44761
rect 25774 44724 25780 44736
rect 24872 44696 25780 44724
rect 25774 44684 25780 44696
rect 25832 44684 25838 44736
rect 27172 44724 27200 44764
rect 27332 44761 27344 44795
rect 27378 44792 27390 44795
rect 27522 44792 27528 44804
rect 27378 44764 27528 44792
rect 27378 44761 27390 44764
rect 27332 44755 27390 44761
rect 27522 44752 27528 44764
rect 27580 44752 27586 44804
rect 28074 44724 28080 44736
rect 27172 44696 28080 44724
rect 28074 44684 28080 44696
rect 28132 44684 28138 44736
rect 28184 44724 28212 44832
rect 30650 44820 30656 44872
rect 30708 44860 30714 44872
rect 30929 44863 30987 44869
rect 30929 44860 30941 44863
rect 30708 44832 30941 44860
rect 30708 44820 30714 44832
rect 30929 44829 30941 44832
rect 30975 44829 30987 44863
rect 31128 44860 31156 44900
rect 31205 44897 31217 44931
rect 31251 44928 31263 44931
rect 32030 44928 32036 44940
rect 31251 44900 32036 44928
rect 31251 44897 31263 44900
rect 31205 44891 31263 44897
rect 32030 44888 32036 44900
rect 32088 44888 32094 44940
rect 34698 44888 34704 44940
rect 34756 44928 34762 44940
rect 35529 44931 35587 44937
rect 35529 44928 35541 44931
rect 34756 44900 35541 44928
rect 34756 44888 34762 44900
rect 35529 44897 35541 44900
rect 35575 44897 35587 44931
rect 35529 44891 35587 44897
rect 33689 44863 33747 44869
rect 33689 44860 33701 44863
rect 31128 44832 33701 44860
rect 30929 44823 30987 44829
rect 33689 44829 33701 44832
rect 33735 44860 33747 44863
rect 33778 44860 33784 44872
rect 33735 44832 33784 44860
rect 33735 44829 33747 44832
rect 33689 44823 33747 44829
rect 33778 44820 33784 44832
rect 33836 44820 33842 44872
rect 34054 44820 34060 44872
rect 34112 44860 34118 44872
rect 34885 44863 34943 44869
rect 34885 44860 34897 44863
rect 34112 44832 34897 44860
rect 34112 44820 34118 44832
rect 34885 44829 34897 44832
rect 34931 44829 34943 44863
rect 34885 44823 34943 44829
rect 29270 44752 29276 44804
rect 29328 44792 29334 44804
rect 29549 44795 29607 44801
rect 29549 44792 29561 44795
rect 29328 44764 29561 44792
rect 29328 44752 29334 44764
rect 29549 44761 29561 44764
rect 29595 44761 29607 44795
rect 34606 44792 34612 44804
rect 29549 44755 29607 44761
rect 31864 44764 34612 44792
rect 31864 44724 31892 44764
rect 34606 44752 34612 44764
rect 34664 44792 34670 44804
rect 34701 44795 34759 44801
rect 34701 44792 34713 44795
rect 34664 44764 34713 44792
rect 34664 44752 34670 44764
rect 34701 44761 34713 44764
rect 34747 44761 34759 44795
rect 34701 44755 34759 44761
rect 28184 44696 31892 44724
rect 32125 44727 32183 44733
rect 32125 44693 32137 44727
rect 32171 44724 32183 44727
rect 32306 44724 32312 44736
rect 32171 44696 32312 44724
rect 32171 44693 32183 44696
rect 32125 44687 32183 44693
rect 32306 44684 32312 44696
rect 32364 44684 32370 44736
rect 33229 44727 33287 44733
rect 33229 44693 33241 44727
rect 33275 44724 33287 44727
rect 33870 44724 33876 44736
rect 33275 44696 33876 44724
rect 33275 44693 33287 44696
rect 33229 44687 33287 44693
rect 33870 44684 33876 44696
rect 33928 44684 33934 44736
rect 35069 44727 35127 44733
rect 35069 44693 35081 44727
rect 35115 44724 35127 44727
rect 35434 44724 35440 44736
rect 35115 44696 35440 44724
rect 35115 44693 35127 44696
rect 35069 44687 35127 44693
rect 35434 44684 35440 44696
rect 35492 44684 35498 44736
rect 36078 44724 36084 44736
rect 36039 44696 36084 44724
rect 36078 44684 36084 44696
rect 36136 44684 36142 44736
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 9861 44523 9919 44529
rect 9861 44489 9873 44523
rect 9907 44520 9919 44523
rect 10410 44520 10416 44532
rect 9907 44492 10416 44520
rect 9907 44489 9919 44492
rect 9861 44483 9919 44489
rect 10410 44480 10416 44492
rect 10468 44480 10474 44532
rect 11885 44523 11943 44529
rect 11885 44489 11897 44523
rect 11931 44520 11943 44523
rect 12618 44520 12624 44532
rect 11931 44492 12624 44520
rect 11931 44489 11943 44492
rect 11885 44483 11943 44489
rect 12618 44480 12624 44492
rect 12676 44480 12682 44532
rect 12713 44523 12771 44529
rect 12713 44489 12725 44523
rect 12759 44520 12771 44523
rect 12802 44520 12808 44532
rect 12759 44492 12808 44520
rect 12759 44489 12771 44492
rect 12713 44483 12771 44489
rect 12802 44480 12808 44492
rect 12860 44480 12866 44532
rect 13262 44520 13268 44532
rect 13223 44492 13268 44520
rect 13262 44480 13268 44492
rect 13320 44480 13326 44532
rect 16022 44520 16028 44532
rect 15983 44492 16028 44520
rect 16022 44480 16028 44492
rect 16080 44480 16086 44532
rect 16224 44492 18460 44520
rect 12636 44452 12664 44480
rect 16224 44452 16252 44492
rect 12636 44424 16252 44452
rect 16298 44412 16304 44464
rect 16356 44452 16362 44464
rect 18432 44452 18460 44492
rect 19242 44480 19248 44532
rect 19300 44520 19306 44532
rect 19889 44523 19947 44529
rect 19889 44520 19901 44523
rect 19300 44492 19901 44520
rect 19300 44480 19306 44492
rect 19889 44489 19901 44492
rect 19935 44489 19947 44523
rect 19889 44483 19947 44489
rect 21726 44480 21732 44532
rect 21784 44520 21790 44532
rect 22278 44520 22284 44532
rect 21784 44492 22284 44520
rect 21784 44480 21790 44492
rect 22278 44480 22284 44492
rect 22336 44480 22342 44532
rect 23750 44480 23756 44532
rect 23808 44520 23814 44532
rect 32217 44523 32275 44529
rect 32217 44520 32229 44523
rect 23808 44492 32229 44520
rect 23808 44480 23814 44492
rect 32217 44489 32229 44492
rect 32263 44489 32275 44523
rect 32217 44483 32275 44489
rect 33962 44480 33968 44532
rect 34020 44520 34026 44532
rect 34333 44523 34391 44529
rect 34333 44520 34345 44523
rect 34020 44492 34345 44520
rect 34020 44480 34026 44492
rect 34333 44489 34345 44492
rect 34379 44489 34391 44523
rect 34333 44483 34391 44489
rect 34422 44480 34428 44532
rect 34480 44520 34486 44532
rect 47946 44520 47952 44532
rect 34480 44492 36216 44520
rect 47907 44492 47952 44520
rect 34480 44480 34486 44492
rect 19429 44455 19487 44461
rect 16356 44424 18368 44452
rect 18432 44424 19380 44452
rect 16356 44412 16362 44424
rect 1394 44384 1400 44396
rect 1355 44356 1400 44384
rect 1394 44344 1400 44356
rect 1452 44344 1458 44396
rect 9858 44344 9864 44396
rect 9916 44384 9922 44396
rect 12529 44387 12587 44393
rect 12529 44384 12541 44387
rect 9916 44356 12541 44384
rect 9916 44344 9922 44356
rect 12529 44353 12541 44356
rect 12575 44384 12587 44387
rect 13173 44387 13231 44393
rect 13173 44384 13185 44387
rect 12575 44356 13185 44384
rect 12575 44353 12587 44356
rect 12529 44347 12587 44353
rect 13173 44353 13185 44356
rect 13219 44384 13231 44387
rect 13262 44384 13268 44396
rect 13219 44356 13268 44384
rect 13219 44353 13231 44356
rect 13173 44347 13231 44353
rect 13262 44344 13268 44356
rect 13320 44344 13326 44396
rect 13357 44387 13415 44393
rect 13357 44353 13369 44387
rect 13403 44384 13415 44387
rect 13998 44384 14004 44396
rect 13403 44356 14004 44384
rect 13403 44353 13415 44356
rect 13357 44347 13415 44353
rect 12158 44276 12164 44328
rect 12216 44316 12222 44328
rect 12345 44319 12403 44325
rect 12345 44316 12357 44319
rect 12216 44288 12357 44316
rect 12216 44276 12222 44288
rect 12345 44285 12357 44288
rect 12391 44316 12403 44319
rect 13372 44316 13400 44347
rect 13998 44344 14004 44356
rect 14056 44344 14062 44396
rect 15102 44344 15108 44396
rect 15160 44384 15166 44396
rect 15197 44387 15255 44393
rect 15197 44384 15209 44387
rect 15160 44356 15209 44384
rect 15160 44344 15166 44356
rect 15197 44353 15209 44356
rect 15243 44353 15255 44387
rect 15197 44347 15255 44353
rect 15286 44344 15292 44396
rect 15344 44384 15350 44396
rect 15381 44387 15439 44393
rect 15381 44384 15393 44387
rect 15344 44356 15393 44384
rect 15344 44344 15350 44356
rect 15381 44353 15393 44356
rect 15427 44384 15439 44387
rect 15470 44384 15476 44396
rect 15427 44356 15476 44384
rect 15427 44353 15439 44356
rect 15381 44347 15439 44353
rect 15470 44344 15476 44356
rect 15528 44344 15534 44396
rect 15565 44387 15623 44393
rect 15565 44353 15577 44387
rect 15611 44384 15623 44387
rect 16853 44387 16911 44393
rect 16853 44384 16865 44387
rect 15611 44356 16865 44384
rect 15611 44353 15623 44356
rect 15565 44347 15623 44353
rect 16853 44353 16865 44356
rect 16899 44353 16911 44387
rect 17494 44384 17500 44396
rect 17455 44356 17500 44384
rect 16853 44347 16911 44353
rect 17494 44344 17500 44356
rect 17552 44344 17558 44396
rect 18046 44384 18052 44396
rect 18007 44356 18052 44384
rect 18046 44344 18052 44356
rect 18104 44344 18110 44396
rect 18138 44344 18144 44396
rect 18196 44384 18202 44396
rect 18340 44393 18368 44424
rect 18325 44387 18383 44393
rect 18196 44356 18241 44384
rect 18196 44344 18202 44356
rect 18325 44353 18337 44387
rect 18371 44384 18383 44387
rect 19242 44384 19248 44396
rect 18371 44356 19104 44384
rect 19203 44356 19248 44384
rect 18371 44353 18383 44356
rect 18325 44347 18383 44353
rect 12391 44288 13400 44316
rect 12391 44285 12403 44288
rect 12345 44279 12403 44285
rect 13446 44276 13452 44328
rect 13504 44316 13510 44328
rect 15010 44316 15016 44328
rect 13504 44288 15016 44316
rect 13504 44276 13510 44288
rect 15010 44276 15016 44288
rect 15068 44276 15074 44328
rect 16482 44276 16488 44328
rect 16540 44316 16546 44328
rect 16669 44319 16727 44325
rect 16669 44316 16681 44319
rect 16540 44288 16681 44316
rect 16540 44276 16546 44288
rect 16669 44285 16681 44288
rect 16715 44285 16727 44319
rect 18966 44316 18972 44328
rect 18927 44288 18972 44316
rect 16669 44279 16727 44285
rect 18966 44276 18972 44288
rect 19024 44276 19030 44328
rect 19076 44316 19104 44356
rect 19242 44344 19248 44356
rect 19300 44344 19306 44396
rect 19352 44384 19380 44424
rect 19429 44421 19441 44455
rect 19475 44452 19487 44455
rect 24762 44452 24768 44464
rect 19475 44424 24768 44452
rect 19475 44421 19487 44424
rect 19429 44415 19487 44421
rect 24762 44412 24768 44424
rect 24820 44412 24826 44464
rect 25314 44412 25320 44464
rect 25372 44452 25378 44464
rect 25372 44424 29132 44452
rect 25372 44412 25378 44424
rect 20073 44387 20131 44393
rect 20073 44384 20085 44387
rect 19352 44356 20085 44384
rect 20073 44353 20085 44356
rect 20119 44353 20131 44387
rect 20073 44347 20131 44353
rect 20088 44316 20116 44347
rect 20162 44344 20168 44396
rect 20220 44384 20226 44396
rect 20257 44387 20315 44393
rect 20257 44384 20269 44387
rect 20220 44356 20269 44384
rect 20220 44344 20226 44356
rect 20257 44353 20269 44356
rect 20303 44384 20315 44387
rect 20714 44384 20720 44396
rect 20303 44356 20720 44384
rect 20303 44353 20315 44356
rect 20257 44347 20315 44353
rect 20714 44344 20720 44356
rect 20772 44344 20778 44396
rect 20901 44387 20959 44393
rect 20901 44353 20913 44387
rect 20947 44384 20959 44387
rect 21174 44384 21180 44396
rect 20947 44356 21180 44384
rect 20947 44353 20959 44356
rect 20901 44347 20959 44353
rect 20346 44316 20352 44328
rect 19076 44288 19196 44316
rect 20088 44288 20352 44316
rect 10413 44251 10471 44257
rect 10413 44217 10425 44251
rect 10459 44248 10471 44251
rect 12434 44248 12440 44260
rect 10459 44220 12440 44248
rect 10459 44217 10471 44220
rect 10413 44211 10471 44217
rect 12434 44208 12440 44220
rect 12492 44248 12498 44260
rect 14645 44251 14703 44257
rect 14645 44248 14657 44251
rect 12492 44220 14657 44248
rect 12492 44208 12498 44220
rect 14645 44217 14657 44220
rect 14691 44217 14703 44251
rect 14645 44211 14703 44217
rect 17037 44251 17095 44257
rect 17037 44217 17049 44251
rect 17083 44248 17095 44251
rect 19061 44251 19119 44257
rect 19061 44248 19073 44251
rect 17083 44220 19073 44248
rect 17083 44217 17095 44220
rect 17037 44211 17095 44217
rect 19061 44217 19073 44220
rect 19107 44217 19119 44251
rect 19168 44248 19196 44288
rect 20346 44276 20352 44288
rect 20404 44316 20410 44328
rect 20916 44316 20944 44347
rect 21174 44344 21180 44356
rect 21232 44344 21238 44396
rect 21818 44384 21824 44396
rect 21779 44356 21824 44384
rect 21818 44344 21824 44356
rect 21876 44344 21882 44396
rect 22002 44384 22008 44396
rect 21963 44356 22008 44384
rect 22002 44344 22008 44356
rect 22060 44344 22066 44396
rect 23750 44384 23756 44396
rect 23711 44356 23756 44384
rect 23750 44344 23756 44356
rect 23808 44344 23814 44396
rect 23934 44384 23940 44396
rect 23895 44356 23940 44384
rect 23934 44344 23940 44356
rect 23992 44344 23998 44396
rect 24581 44387 24639 44393
rect 24581 44353 24593 44387
rect 24627 44384 24639 44387
rect 24854 44384 24860 44396
rect 24627 44356 24860 44384
rect 24627 44353 24639 44356
rect 24581 44347 24639 44353
rect 24854 44344 24860 44356
rect 24912 44344 24918 44396
rect 27890 44344 27896 44396
rect 27948 44384 27954 44396
rect 28270 44387 28328 44393
rect 28270 44384 28282 44387
rect 27948 44356 28282 44384
rect 27948 44344 27954 44356
rect 28270 44353 28282 44356
rect 28316 44353 28328 44387
rect 28270 44347 28328 44353
rect 28537 44387 28595 44393
rect 28537 44353 28549 44387
rect 28583 44353 28595 44387
rect 29104 44384 29132 44424
rect 32030 44412 32036 44464
rect 32088 44452 32094 44464
rect 32088 44424 33640 44452
rect 32088 44412 32094 44424
rect 29273 44387 29331 44393
rect 29273 44384 29285 44387
rect 29104 44356 29285 44384
rect 28537 44347 28595 44353
rect 29273 44353 29285 44356
rect 29319 44353 29331 44387
rect 33318 44384 33324 44396
rect 33376 44393 33382 44396
rect 33612 44393 33640 44424
rect 33288 44356 33324 44384
rect 29273 44347 29331 44353
rect 20404 44288 20944 44316
rect 20404 44276 20410 44288
rect 22278 44276 22284 44328
rect 22336 44316 22342 44328
rect 23106 44316 23112 44328
rect 22336 44288 23112 44316
rect 22336 44276 22342 44288
rect 23106 44276 23112 44288
rect 23164 44276 23170 44328
rect 23293 44319 23351 44325
rect 23293 44285 23305 44319
rect 23339 44316 23351 44319
rect 23474 44316 23480 44328
rect 23339 44288 23480 44316
rect 23339 44285 23351 44288
rect 23293 44279 23351 44285
rect 23474 44276 23480 44288
rect 23532 44316 23538 44328
rect 24762 44316 24768 44328
rect 23532 44288 24768 44316
rect 23532 44276 23538 44288
rect 24762 44276 24768 44288
rect 24820 44276 24826 44328
rect 25498 44248 25504 44260
rect 19168 44220 25504 44248
rect 19061 44211 19119 44217
rect 25498 44208 25504 44220
rect 25556 44208 25562 44260
rect 25590 44208 25596 44260
rect 25648 44248 25654 44260
rect 27157 44251 27215 44257
rect 27157 44248 27169 44251
rect 25648 44220 27169 44248
rect 25648 44208 25654 44220
rect 27157 44217 27169 44220
rect 27203 44217 27215 44251
rect 27157 44211 27215 44217
rect 1581 44183 1639 44189
rect 1581 44149 1593 44183
rect 1627 44180 1639 44183
rect 1670 44180 1676 44192
rect 1627 44152 1676 44180
rect 1627 44149 1639 44152
rect 1581 44143 1639 44149
rect 1670 44140 1676 44152
rect 1728 44140 1734 44192
rect 9309 44183 9367 44189
rect 9309 44149 9321 44183
rect 9355 44180 9367 44183
rect 9858 44180 9864 44192
rect 9355 44152 9864 44180
rect 9355 44149 9367 44152
rect 9309 44143 9367 44149
rect 9858 44140 9864 44152
rect 9916 44140 9922 44192
rect 10962 44180 10968 44192
rect 10923 44152 10968 44180
rect 10962 44140 10968 44152
rect 11020 44140 11026 44192
rect 14090 44180 14096 44192
rect 14051 44152 14096 44180
rect 14090 44140 14096 44152
rect 14148 44140 14154 44192
rect 18230 44140 18236 44192
rect 18288 44180 18294 44192
rect 18509 44183 18567 44189
rect 18509 44180 18521 44183
rect 18288 44152 18521 44180
rect 18288 44140 18294 44152
rect 18509 44149 18521 44152
rect 18555 44149 18567 44183
rect 20806 44180 20812 44192
rect 20767 44152 20812 44180
rect 18509 44143 18567 44149
rect 20806 44140 20812 44152
rect 20864 44140 20870 44192
rect 21634 44140 21640 44192
rect 21692 44180 21698 44192
rect 22189 44183 22247 44189
rect 22189 44180 22201 44183
rect 21692 44152 22201 44180
rect 21692 44140 21698 44152
rect 22189 44149 22201 44152
rect 22235 44180 22247 44183
rect 22922 44180 22928 44192
rect 22235 44152 22928 44180
rect 22235 44149 22247 44152
rect 22189 44143 22247 44149
rect 22922 44140 22928 44152
rect 22980 44140 22986 44192
rect 23934 44180 23940 44192
rect 23895 44152 23940 44180
rect 23934 44140 23940 44152
rect 23992 44140 23998 44192
rect 24394 44180 24400 44192
rect 24355 44152 24400 44180
rect 24394 44140 24400 44152
rect 24452 44140 24458 44192
rect 25038 44140 25044 44192
rect 25096 44180 25102 44192
rect 25409 44183 25467 44189
rect 25409 44180 25421 44183
rect 25096 44152 25421 44180
rect 25096 44140 25102 44152
rect 25409 44149 25421 44152
rect 25455 44149 25467 44183
rect 26050 44180 26056 44192
rect 26011 44152 26056 44180
rect 25409 44143 25467 44149
rect 26050 44140 26056 44152
rect 26108 44140 26114 44192
rect 28552 44180 28580 44347
rect 33318 44344 33324 44356
rect 33376 44347 33388 44393
rect 33597 44387 33655 44393
rect 33597 44353 33609 44387
rect 33643 44353 33655 44387
rect 33597 44347 33655 44353
rect 34517 44387 34575 44393
rect 34517 44353 34529 44387
rect 34563 44384 34575 44387
rect 34698 44384 34704 44396
rect 34563 44356 34704 44384
rect 34563 44353 34575 44356
rect 34517 44347 34575 44353
rect 33376 44344 33382 44347
rect 34698 44344 34704 44356
rect 34756 44344 34762 44396
rect 35434 44384 35440 44396
rect 35395 44356 35440 44384
rect 35434 44344 35440 44356
rect 35492 44344 35498 44396
rect 35526 44344 35532 44396
rect 35584 44384 35590 44396
rect 35584 44356 35629 44384
rect 35584 44344 35590 44356
rect 28994 44316 29000 44328
rect 28955 44288 29000 44316
rect 28994 44276 29000 44288
rect 29052 44276 29058 44328
rect 30653 44319 30711 44325
rect 30653 44285 30665 44319
rect 30699 44316 30711 44319
rect 31478 44316 31484 44328
rect 30699 44288 31484 44316
rect 30699 44285 30711 44288
rect 30653 44279 30711 44285
rect 31478 44276 31484 44288
rect 31536 44276 31542 44328
rect 34790 44316 34796 44328
rect 34751 44288 34796 44316
rect 34790 44276 34796 44288
rect 34848 44276 34854 44328
rect 34701 44251 34759 44257
rect 34701 44217 34713 44251
rect 34747 44248 34759 44251
rect 35894 44248 35900 44260
rect 34747 44220 35900 44248
rect 34747 44217 34759 44220
rect 34701 44211 34759 44217
rect 35894 44208 35900 44220
rect 35952 44208 35958 44260
rect 36188 44257 36216 44492
rect 47946 44480 47952 44492
rect 48004 44480 48010 44532
rect 48038 44384 48044 44396
rect 47999 44356 48044 44384
rect 48038 44344 48044 44356
rect 48096 44344 48102 44396
rect 36173 44251 36231 44257
rect 36173 44217 36185 44251
rect 36219 44248 36231 44251
rect 36219 44220 37964 44248
rect 36219 44217 36231 44220
rect 36173 44211 36231 44217
rect 37936 44192 37964 44220
rect 28994 44180 29000 44192
rect 28552 44152 29000 44180
rect 28994 44140 29000 44152
rect 29052 44140 29058 44192
rect 30466 44140 30472 44192
rect 30524 44180 30530 44192
rect 31481 44183 31539 44189
rect 31481 44180 31493 44183
rect 30524 44152 31493 44180
rect 30524 44140 30530 44152
rect 31481 44149 31493 44152
rect 31527 44180 31539 44183
rect 33594 44180 33600 44192
rect 31527 44152 33600 44180
rect 31527 44149 31539 44152
rect 31481 44143 31539 44149
rect 33594 44140 33600 44152
rect 33652 44140 33658 44192
rect 35253 44183 35311 44189
rect 35253 44149 35265 44183
rect 35299 44180 35311 44183
rect 35342 44180 35348 44192
rect 35299 44152 35348 44180
rect 35299 44149 35311 44152
rect 35253 44143 35311 44149
rect 35342 44140 35348 44152
rect 35400 44140 35406 44192
rect 36722 44180 36728 44192
rect 36683 44152 36728 44180
rect 36722 44140 36728 44152
rect 36780 44140 36786 44192
rect 37274 44140 37280 44192
rect 37332 44180 37338 44192
rect 37369 44183 37427 44189
rect 37369 44180 37381 44183
rect 37332 44152 37381 44180
rect 37332 44140 37338 44152
rect 37369 44149 37381 44152
rect 37415 44180 37427 44183
rect 37734 44180 37740 44192
rect 37415 44152 37740 44180
rect 37415 44149 37427 44152
rect 37369 44143 37427 44149
rect 37734 44140 37740 44152
rect 37792 44140 37798 44192
rect 37918 44180 37924 44192
rect 37879 44152 37924 44180
rect 37918 44140 37924 44152
rect 37976 44140 37982 44192
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 1394 43976 1400 43988
rect 1355 43948 1400 43976
rect 1394 43936 1400 43948
rect 1452 43936 1458 43988
rect 11698 43936 11704 43988
rect 11756 43976 11762 43988
rect 12437 43979 12495 43985
rect 12437 43976 12449 43979
rect 11756 43948 12449 43976
rect 11756 43936 11762 43948
rect 12437 43945 12449 43948
rect 12483 43976 12495 43979
rect 14090 43976 14096 43988
rect 12483 43948 14096 43976
rect 12483 43945 12495 43948
rect 12437 43939 12495 43945
rect 14090 43936 14096 43948
rect 14148 43936 14154 43988
rect 14458 43936 14464 43988
rect 14516 43976 14522 43988
rect 14516 43948 14561 43976
rect 14516 43936 14522 43948
rect 16022 43936 16028 43988
rect 16080 43976 16086 43988
rect 16945 43979 17003 43985
rect 16945 43976 16957 43979
rect 16080 43948 16957 43976
rect 16080 43936 16086 43948
rect 16945 43945 16957 43948
rect 16991 43945 17003 43979
rect 17954 43976 17960 43988
rect 17867 43948 17960 43976
rect 16945 43939 17003 43945
rect 17926 43936 17960 43948
rect 18012 43976 18018 43988
rect 18966 43976 18972 43988
rect 18012 43948 18972 43976
rect 18012 43936 18018 43948
rect 18966 43936 18972 43948
rect 19024 43936 19030 43988
rect 20530 43976 20536 43988
rect 19536 43948 20536 43976
rect 13541 43911 13599 43917
rect 13541 43877 13553 43911
rect 13587 43908 13599 43911
rect 15102 43908 15108 43920
rect 13587 43880 15108 43908
rect 13587 43877 13599 43880
rect 13541 43871 13599 43877
rect 15102 43868 15108 43880
rect 15160 43868 15166 43920
rect 17589 43911 17647 43917
rect 17589 43877 17601 43911
rect 17635 43908 17647 43911
rect 17926 43908 17954 43936
rect 17635 43880 17954 43908
rect 17635 43877 17647 43880
rect 17589 43871 17647 43877
rect 13078 43840 13084 43852
rect 13039 43812 13084 43840
rect 13078 43800 13084 43812
rect 13136 43800 13142 43852
rect 14826 43800 14832 43852
rect 14884 43840 14890 43852
rect 15749 43843 15807 43849
rect 15749 43840 15761 43843
rect 14884 43812 15761 43840
rect 14884 43800 14890 43812
rect 15749 43809 15761 43812
rect 15795 43840 15807 43843
rect 17862 43840 17868 43852
rect 15795 43812 17868 43840
rect 15795 43809 15807 43812
rect 15749 43803 15807 43809
rect 17862 43800 17868 43812
rect 17920 43800 17926 43852
rect 19536 43840 19564 43948
rect 20530 43936 20536 43948
rect 20588 43936 20594 43988
rect 20622 43936 20628 43988
rect 20680 43976 20686 43988
rect 20680 43948 25452 43976
rect 20680 43936 20686 43948
rect 20806 43908 20812 43920
rect 18340 43812 19564 43840
rect 19628 43880 20812 43908
rect 10870 43772 10876 43784
rect 10783 43744 10876 43772
rect 10870 43732 10876 43744
rect 10928 43772 10934 43784
rect 11425 43775 11483 43781
rect 10928 43744 11100 43772
rect 10928 43732 10934 43744
rect 10321 43707 10379 43713
rect 10321 43673 10333 43707
rect 10367 43704 10379 43707
rect 10962 43704 10968 43716
rect 10367 43676 10968 43704
rect 10367 43673 10379 43676
rect 10321 43667 10379 43673
rect 10962 43664 10968 43676
rect 11020 43664 11026 43716
rect 11072 43704 11100 43744
rect 11425 43741 11437 43775
rect 11471 43772 11483 43775
rect 12802 43772 12808 43784
rect 11471 43744 12808 43772
rect 11471 43741 11483 43744
rect 11425 43735 11483 43741
rect 12802 43732 12808 43744
rect 12860 43732 12866 43784
rect 12894 43732 12900 43784
rect 12952 43772 12958 43784
rect 13173 43775 13231 43781
rect 13173 43772 13185 43775
rect 12952 43744 13185 43772
rect 12952 43732 12958 43744
rect 13173 43741 13185 43744
rect 13219 43741 13231 43775
rect 14918 43772 14924 43784
rect 14879 43744 14924 43772
rect 13173 43735 13231 43741
rect 14918 43732 14924 43744
rect 14976 43732 14982 43784
rect 15105 43775 15163 43781
rect 15105 43741 15117 43775
rect 15151 43772 15163 43775
rect 15194 43772 15200 43784
rect 15151 43744 15200 43772
rect 15151 43741 15163 43744
rect 15105 43735 15163 43741
rect 15194 43732 15200 43744
rect 15252 43732 15258 43784
rect 16298 43772 16304 43784
rect 15580 43744 16304 43772
rect 15580 43704 15608 43744
rect 16298 43732 16304 43744
rect 16356 43732 16362 43784
rect 16482 43772 16488 43784
rect 16443 43744 16488 43772
rect 16482 43732 16488 43744
rect 16540 43732 16546 43784
rect 16574 43732 16580 43784
rect 16632 43772 16638 43784
rect 18049 43775 18107 43781
rect 18049 43772 18061 43775
rect 16632 43744 18061 43772
rect 16632 43732 16638 43744
rect 18049 43741 18061 43744
rect 18095 43741 18107 43775
rect 18230 43772 18236 43784
rect 18191 43744 18236 43772
rect 18049 43735 18107 43741
rect 18230 43732 18236 43744
rect 18288 43732 18294 43784
rect 18340 43781 18368 43812
rect 19628 43781 19656 43880
rect 20806 43868 20812 43880
rect 20864 43868 20870 43920
rect 24762 43908 24768 43920
rect 23584 43880 24768 43908
rect 21174 43840 21180 43852
rect 20548 43812 21180 43840
rect 20548 43781 20576 43812
rect 21174 43800 21180 43812
rect 21232 43840 21238 43852
rect 22002 43840 22008 43852
rect 21232 43812 22008 43840
rect 21232 43800 21238 43812
rect 22002 43800 22008 43812
rect 22060 43800 22066 43852
rect 18325 43775 18383 43781
rect 18325 43741 18337 43775
rect 18371 43741 18383 43775
rect 18325 43735 18383 43741
rect 18417 43775 18475 43781
rect 18417 43741 18429 43775
rect 18463 43741 18475 43775
rect 18417 43735 18475 43741
rect 19613 43775 19671 43781
rect 19613 43741 19625 43775
rect 19659 43741 19671 43775
rect 19613 43735 19671 43741
rect 20533 43775 20591 43781
rect 20533 43741 20545 43775
rect 20579 43741 20591 43775
rect 20533 43735 20591 43741
rect 20717 43775 20775 43781
rect 20717 43741 20729 43775
rect 20763 43772 20775 43775
rect 21542 43772 21548 43784
rect 20763 43744 21548 43772
rect 20763 43741 20775 43744
rect 20717 43735 20775 43741
rect 11072 43676 15608 43704
rect 15654 43664 15660 43716
rect 15712 43704 15718 43716
rect 16393 43707 16451 43713
rect 16393 43704 16405 43707
rect 15712 43676 16405 43704
rect 15712 43664 15718 43676
rect 16393 43673 16405 43676
rect 16439 43704 16451 43707
rect 18432 43704 18460 43735
rect 21542 43732 21548 43744
rect 21600 43732 21606 43784
rect 22097 43775 22155 43781
rect 22097 43741 22109 43775
rect 22143 43741 22155 43775
rect 22278 43772 22284 43784
rect 22239 43744 22284 43772
rect 22097 43735 22155 43741
rect 18690 43704 18696 43716
rect 16439 43676 18460 43704
rect 18651 43676 18696 43704
rect 16439 43673 16451 43676
rect 16393 43667 16451 43673
rect 18690 43664 18696 43676
rect 18748 43664 18754 43716
rect 19426 43664 19432 43716
rect 19484 43704 19490 43716
rect 19705 43707 19763 43713
rect 19705 43704 19717 43707
rect 19484 43676 19717 43704
rect 19484 43664 19490 43676
rect 19705 43673 19717 43676
rect 19751 43673 19763 43707
rect 19705 43667 19763 43673
rect 19889 43707 19947 43713
rect 19889 43673 19901 43707
rect 19935 43704 19947 43707
rect 21177 43707 21235 43713
rect 19935 43676 20668 43704
rect 19935 43673 19947 43676
rect 19889 43667 19947 43673
rect 9769 43639 9827 43645
rect 9769 43605 9781 43639
rect 9815 43636 9827 43639
rect 9858 43636 9864 43648
rect 9815 43608 9864 43636
rect 9815 43605 9827 43608
rect 9769 43599 9827 43605
rect 9858 43596 9864 43608
rect 9916 43596 9922 43648
rect 11790 43596 11796 43648
rect 11848 43636 11854 43648
rect 11885 43639 11943 43645
rect 11885 43636 11897 43639
rect 11848 43608 11897 43636
rect 11848 43596 11854 43608
rect 11885 43605 11897 43608
rect 11931 43605 11943 43639
rect 11885 43599 11943 43605
rect 15105 43639 15163 43645
rect 15105 43605 15117 43639
rect 15151 43636 15163 43639
rect 15562 43636 15568 43648
rect 15151 43608 15568 43636
rect 15151 43605 15163 43608
rect 15105 43599 15163 43605
rect 15562 43596 15568 43608
rect 15620 43596 15626 43648
rect 19797 43639 19855 43645
rect 19797 43605 19809 43639
rect 19843 43636 19855 43639
rect 19978 43636 19984 43648
rect 19843 43608 19984 43636
rect 19843 43605 19855 43608
rect 19797 43599 19855 43605
rect 19978 43596 19984 43608
rect 20036 43596 20042 43648
rect 20640 43645 20668 43676
rect 21177 43673 21189 43707
rect 21223 43673 21235 43707
rect 21177 43667 21235 43673
rect 20625 43639 20683 43645
rect 20625 43605 20637 43639
rect 20671 43636 20683 43639
rect 20714 43636 20720 43648
rect 20671 43608 20720 43636
rect 20671 43605 20683 43608
rect 20625 43599 20683 43605
rect 20714 43596 20720 43608
rect 20772 43596 20778 43648
rect 21192 43636 21220 43667
rect 21266 43664 21272 43716
rect 21324 43704 21330 43716
rect 21361 43707 21419 43713
rect 21361 43704 21373 43707
rect 21324 43676 21373 43704
rect 21324 43664 21330 43676
rect 21361 43673 21373 43676
rect 21407 43673 21419 43707
rect 22112 43704 22140 43735
rect 22278 43732 22284 43744
rect 22336 43772 22342 43784
rect 22738 43772 22744 43784
rect 22336 43744 22744 43772
rect 22336 43732 22342 43744
rect 22738 43732 22744 43744
rect 22796 43732 22802 43784
rect 23382 43732 23388 43784
rect 23440 43772 23446 43784
rect 23584 43781 23612 43880
rect 24762 43868 24768 43880
rect 24820 43868 24826 43920
rect 25424 43908 25452 43948
rect 25498 43936 25504 43988
rect 25556 43976 25562 43988
rect 25593 43979 25651 43985
rect 25593 43976 25605 43979
rect 25556 43948 25605 43976
rect 25556 43936 25562 43948
rect 25593 43945 25605 43948
rect 25639 43976 25651 43979
rect 25639 43948 32076 43976
rect 25639 43945 25651 43948
rect 25593 43939 25651 43945
rect 26970 43908 26976 43920
rect 25424 43880 26976 43908
rect 26970 43868 26976 43880
rect 27028 43868 27034 43920
rect 32048 43908 32076 43948
rect 34790 43936 34796 43988
rect 34848 43976 34854 43988
rect 35897 43979 35955 43985
rect 35897 43976 35909 43979
rect 34848 43948 35909 43976
rect 34848 43936 34854 43948
rect 35897 43945 35909 43948
rect 35943 43945 35955 43979
rect 48038 43976 48044 43988
rect 47999 43948 48044 43976
rect 35897 43939 35955 43945
rect 48038 43936 48044 43948
rect 48096 43936 48102 43988
rect 32048 43880 36308 43908
rect 24486 43840 24492 43852
rect 23676 43812 24492 43840
rect 23676 43781 23704 43812
rect 24486 43800 24492 43812
rect 24544 43840 24550 43852
rect 24857 43843 24915 43849
rect 24857 43840 24869 43843
rect 24544 43812 24869 43840
rect 24544 43800 24550 43812
rect 24857 43809 24869 43812
rect 24903 43809 24915 43843
rect 24857 43803 24915 43809
rect 27062 43800 27068 43852
rect 27120 43840 27126 43852
rect 27341 43843 27399 43849
rect 27341 43840 27353 43843
rect 27120 43812 27353 43840
rect 27120 43800 27126 43812
rect 27341 43809 27353 43812
rect 27387 43809 27399 43843
rect 34054 43840 34060 43852
rect 27341 43803 27399 43809
rect 27448 43812 34060 43840
rect 23569 43775 23627 43781
rect 23569 43772 23581 43775
rect 23440 43744 23581 43772
rect 23440 43732 23446 43744
rect 23569 43741 23581 43744
rect 23615 43741 23627 43775
rect 23569 43735 23627 43741
rect 23661 43775 23719 43781
rect 23661 43741 23673 43775
rect 23707 43741 23719 43775
rect 23661 43735 23719 43741
rect 23772 43775 23830 43781
rect 23772 43741 23784 43775
rect 23818 43772 23830 43775
rect 24581 43775 24639 43781
rect 24581 43772 24593 43775
rect 23818 43744 24593 43772
rect 23818 43741 23830 43744
rect 23772 43735 23830 43741
rect 24581 43741 24593 43744
rect 24627 43741 24639 43775
rect 24581 43735 24639 43741
rect 24946 43732 24952 43784
rect 25004 43772 25010 43784
rect 25317 43775 25375 43781
rect 25317 43772 25329 43775
rect 25004 43744 25329 43772
rect 25004 43732 25010 43744
rect 25317 43741 25329 43744
rect 25363 43741 25375 43775
rect 25317 43735 25375 43741
rect 26881 43775 26939 43781
rect 26881 43741 26893 43775
rect 26927 43772 26939 43775
rect 26970 43772 26976 43784
rect 26927 43744 26976 43772
rect 26927 43741 26939 43744
rect 26881 43735 26939 43741
rect 26970 43732 26976 43744
rect 27028 43772 27034 43784
rect 27448 43772 27476 43812
rect 34054 43800 34060 43812
rect 34112 43800 34118 43852
rect 27028 43744 27476 43772
rect 27617 43775 27675 43781
rect 27028 43732 27034 43744
rect 27617 43741 27629 43775
rect 27663 43772 27675 43775
rect 29362 43772 29368 43784
rect 27663 43744 29368 43772
rect 27663 43741 27675 43744
rect 27617 43735 27675 43741
rect 29362 43732 29368 43744
rect 29420 43732 29426 43784
rect 33965 43775 34023 43781
rect 33965 43741 33977 43775
rect 34011 43772 34023 43775
rect 34606 43772 34612 43784
rect 34011 43744 34612 43772
rect 34011 43741 34023 43744
rect 33965 43735 34023 43741
rect 34606 43732 34612 43744
rect 34664 43732 34670 43784
rect 22186 43704 22192 43716
rect 22099 43676 22192 43704
rect 21361 43667 21419 43673
rect 22186 43664 22192 43676
rect 22244 43704 22250 43716
rect 22830 43704 22836 43716
rect 22244 43676 22836 43704
rect 22244 43664 22250 43676
rect 22830 43664 22836 43676
rect 22888 43664 22894 43716
rect 23855 43707 23913 43713
rect 23855 43673 23867 43707
rect 23901 43704 23913 43707
rect 24118 43704 24124 43716
rect 23901 43676 24124 43704
rect 23901 43673 23913 43676
rect 23855 43667 23913 43673
rect 24118 43664 24124 43676
rect 24176 43664 24182 43716
rect 24854 43664 24860 43716
rect 24912 43704 24918 43716
rect 25501 43707 25559 43713
rect 25501 43704 25513 43707
rect 24912 43676 25513 43704
rect 24912 43664 24918 43676
rect 25501 43673 25513 43676
rect 25547 43704 25559 43707
rect 26237 43707 26295 43713
rect 26237 43704 26249 43707
rect 25547 43676 26249 43704
rect 25547 43673 25559 43676
rect 25501 43667 25559 43673
rect 26237 43673 26249 43676
rect 26283 43704 26295 43707
rect 26283 43676 26924 43704
rect 26283 43673 26295 43676
rect 26237 43667 26295 43673
rect 21450 43636 21456 43648
rect 21192 43608 21456 43636
rect 21450 43596 21456 43608
rect 21508 43636 21514 43648
rect 22094 43636 22100 43648
rect 21508 43608 22100 43636
rect 21508 43596 21514 43608
rect 22094 43596 22100 43608
rect 22152 43596 22158 43648
rect 22281 43639 22339 43645
rect 22281 43605 22293 43639
rect 22327 43636 22339 43639
rect 22462 43636 22468 43648
rect 22327 43608 22468 43636
rect 22327 43605 22339 43608
rect 22281 43599 22339 43605
rect 22462 43596 22468 43608
rect 22520 43596 22526 43648
rect 23109 43639 23167 43645
rect 23109 43605 23121 43639
rect 23155 43636 23167 43639
rect 23198 43636 23204 43648
rect 23155 43608 23204 43636
rect 23155 43605 23167 43608
rect 23109 43599 23167 43605
rect 23198 43596 23204 43608
rect 23256 43596 23262 43648
rect 23750 43596 23756 43648
rect 23808 43636 23814 43648
rect 24397 43639 24455 43645
rect 24397 43636 24409 43639
rect 23808 43608 24409 43636
rect 23808 43596 23814 43608
rect 24397 43605 24409 43608
rect 24443 43605 24455 43639
rect 26896 43636 26924 43676
rect 29178 43664 29184 43716
rect 29236 43704 29242 43716
rect 31205 43707 31263 43713
rect 31205 43704 31217 43707
rect 29236 43676 31217 43704
rect 29236 43664 29242 43676
rect 31205 43673 31217 43676
rect 31251 43673 31263 43707
rect 34716 43704 34744 43880
rect 35342 43840 35348 43852
rect 34900 43812 35348 43840
rect 34900 43781 34928 43812
rect 35342 43800 35348 43812
rect 35400 43840 35406 43852
rect 36170 43840 36176 43852
rect 35400 43812 36176 43840
rect 35400 43800 35406 43812
rect 36170 43800 36176 43812
rect 36228 43800 36234 43852
rect 36280 43784 36308 43880
rect 34885 43775 34943 43781
rect 34885 43741 34897 43775
rect 34931 43741 34943 43775
rect 35158 43772 35164 43784
rect 35119 43744 35164 43772
rect 34885 43735 34943 43741
rect 35158 43732 35164 43744
rect 35216 43732 35222 43784
rect 35618 43772 35624 43784
rect 35579 43744 35624 43772
rect 35618 43732 35624 43744
rect 35676 43772 35682 43784
rect 35676 43744 36124 43772
rect 35676 43732 35682 43744
rect 35069 43707 35127 43713
rect 35069 43704 35081 43707
rect 34716 43676 35081 43704
rect 31205 43667 31263 43673
rect 35069 43673 35081 43676
rect 35115 43673 35127 43707
rect 35069 43667 35127 43673
rect 35526 43664 35532 43716
rect 35584 43704 35590 43716
rect 35713 43707 35771 43713
rect 35713 43704 35725 43707
rect 35584 43676 35725 43704
rect 35584 43664 35590 43676
rect 35713 43673 35725 43676
rect 35759 43673 35771 43707
rect 35713 43667 35771 43673
rect 35897 43707 35955 43713
rect 35897 43673 35909 43707
rect 35943 43704 35955 43707
rect 35986 43704 35992 43716
rect 35943 43676 35992 43704
rect 35943 43673 35955 43676
rect 35897 43667 35955 43673
rect 35986 43664 35992 43676
rect 36044 43664 36050 43716
rect 36096 43704 36124 43744
rect 36262 43732 36268 43784
rect 36320 43772 36326 43784
rect 36357 43775 36415 43781
rect 36357 43772 36369 43775
rect 36320 43744 36369 43772
rect 36320 43732 36326 43744
rect 36357 43741 36369 43744
rect 36403 43741 36415 43775
rect 36357 43735 36415 43741
rect 37553 43775 37611 43781
rect 37553 43741 37565 43775
rect 37599 43772 37611 43775
rect 37918 43772 37924 43784
rect 37599 43744 37924 43772
rect 37599 43741 37611 43744
rect 37553 43735 37611 43741
rect 37918 43732 37924 43744
rect 37976 43772 37982 43784
rect 37976 43744 38608 43772
rect 37976 43732 37982 43744
rect 36096 43676 36400 43704
rect 27614 43636 27620 43648
rect 26896 43608 27620 43636
rect 24397 43599 24455 43605
rect 27614 43596 27620 43608
rect 27672 43596 27678 43648
rect 28718 43636 28724 43648
rect 28679 43608 28724 43636
rect 28718 43596 28724 43608
rect 28776 43596 28782 43648
rect 29641 43639 29699 43645
rect 29641 43605 29653 43639
rect 29687 43636 29699 43639
rect 30285 43639 30343 43645
rect 30285 43636 30297 43639
rect 29687 43608 30297 43636
rect 29687 43605 29699 43608
rect 29641 43599 29699 43605
rect 30285 43605 30297 43608
rect 30331 43636 30343 43639
rect 30558 43636 30564 43648
rect 30331 43608 30564 43636
rect 30331 43605 30343 43608
rect 30285 43599 30343 43605
rect 30558 43596 30564 43608
rect 30616 43596 30622 43648
rect 32030 43596 32036 43648
rect 32088 43636 32094 43648
rect 32493 43639 32551 43645
rect 32493 43636 32505 43639
rect 32088 43608 32505 43636
rect 32088 43596 32094 43608
rect 32493 43605 32505 43608
rect 32539 43605 32551 43639
rect 32493 43599 32551 43605
rect 33134 43596 33140 43648
rect 33192 43636 33198 43648
rect 33413 43639 33471 43645
rect 33413 43636 33425 43639
rect 33192 43608 33425 43636
rect 33192 43596 33198 43608
rect 33413 43605 33425 43608
rect 33459 43605 33471 43639
rect 33413 43599 33471 43605
rect 34054 43596 34060 43648
rect 34112 43636 34118 43648
rect 36372 43645 36400 43676
rect 36446 43664 36452 43716
rect 36504 43704 36510 43716
rect 36630 43704 36636 43716
rect 36504 43676 36549 43704
rect 36591 43676 36636 43704
rect 36504 43664 36510 43676
rect 36630 43664 36636 43676
rect 36688 43664 36694 43716
rect 37734 43664 37740 43716
rect 37792 43704 37798 43716
rect 37792 43676 38424 43704
rect 37792 43664 37798 43676
rect 38396 43648 38424 43676
rect 38580 43648 38608 43744
rect 34701 43639 34759 43645
rect 34701 43636 34713 43639
rect 34112 43608 34713 43636
rect 34112 43596 34118 43608
rect 34701 43605 34713 43608
rect 34747 43605 34759 43639
rect 34701 43599 34759 43605
rect 36357 43639 36415 43645
rect 36357 43605 36369 43639
rect 36403 43605 36415 43639
rect 36357 43599 36415 43605
rect 37826 43596 37832 43648
rect 37884 43636 37890 43648
rect 37921 43639 37979 43645
rect 37921 43636 37933 43639
rect 37884 43608 37933 43636
rect 37884 43596 37890 43608
rect 37921 43605 37933 43608
rect 37967 43605 37979 43639
rect 38378 43636 38384 43648
rect 38339 43608 38384 43636
rect 37921 43599 37979 43605
rect 38378 43596 38384 43608
rect 38436 43596 38442 43648
rect 38562 43596 38568 43648
rect 38620 43636 38626 43648
rect 38933 43639 38991 43645
rect 38933 43636 38945 43639
rect 38620 43608 38945 43636
rect 38620 43596 38626 43608
rect 38933 43605 38945 43608
rect 38979 43605 38991 43639
rect 38933 43599 38991 43605
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 10778 43392 10784 43444
rect 10836 43432 10842 43444
rect 10873 43435 10931 43441
rect 10873 43432 10885 43435
rect 10836 43404 10885 43432
rect 10836 43392 10842 43404
rect 10873 43401 10885 43404
rect 10919 43401 10931 43435
rect 12894 43432 12900 43444
rect 12855 43404 12900 43432
rect 10873 43395 10931 43401
rect 12894 43392 12900 43404
rect 12952 43392 12958 43444
rect 13078 43392 13084 43444
rect 13136 43432 13142 43444
rect 13906 43432 13912 43444
rect 13136 43404 13768 43432
rect 13867 43404 13912 43432
rect 13136 43392 13142 43404
rect 10962 43324 10968 43376
rect 11020 43364 11026 43376
rect 11020 43336 13584 43364
rect 11020 43324 11026 43336
rect 12912 43305 12940 43336
rect 12713 43299 12771 43305
rect 12713 43265 12725 43299
rect 12759 43265 12771 43299
rect 12713 43259 12771 43265
rect 12897 43299 12955 43305
rect 12897 43265 12909 43299
rect 12943 43296 12955 43299
rect 12986 43296 12992 43308
rect 12943 43268 12992 43296
rect 12943 43265 12955 43268
rect 12897 43259 12955 43265
rect 9861 43231 9919 43237
rect 9861 43197 9873 43231
rect 9907 43228 9919 43231
rect 10413 43231 10471 43237
rect 10413 43228 10425 43231
rect 9907 43200 10425 43228
rect 9907 43197 9919 43200
rect 9861 43191 9919 43197
rect 10413 43197 10425 43200
rect 10459 43228 10471 43231
rect 12728 43228 12756 43259
rect 12986 43256 12992 43268
rect 13044 43256 13050 43308
rect 13556 43305 13584 43336
rect 13740 43305 13768 43404
rect 13906 43392 13912 43404
rect 13964 43392 13970 43444
rect 15194 43392 15200 43444
rect 15252 43432 15258 43444
rect 18969 43435 19027 43441
rect 15252 43404 18920 43432
rect 15252 43392 15258 43404
rect 13541 43299 13599 43305
rect 13541 43265 13553 43299
rect 13587 43265 13599 43299
rect 13541 43259 13599 43265
rect 13725 43299 13783 43305
rect 13725 43265 13737 43299
rect 13771 43265 13783 43299
rect 13725 43259 13783 43265
rect 14645 43299 14703 43305
rect 14645 43265 14657 43299
rect 14691 43296 14703 43299
rect 15212 43296 15240 43392
rect 17954 43364 17960 43376
rect 17512 43336 17960 43364
rect 14691 43268 15240 43296
rect 15749 43299 15807 43305
rect 14691 43265 14703 43268
rect 14645 43259 14703 43265
rect 15749 43265 15761 43299
rect 15795 43265 15807 43299
rect 15749 43259 15807 43265
rect 16669 43299 16727 43305
rect 16669 43265 16681 43299
rect 16715 43296 16727 43299
rect 16758 43296 16764 43308
rect 16715 43268 16764 43296
rect 16715 43265 16727 43268
rect 16669 43259 16727 43265
rect 13446 43228 13452 43240
rect 10459 43200 12756 43228
rect 13407 43200 13452 43228
rect 10459 43197 10471 43200
rect 10413 43191 10471 43197
rect 11701 43163 11759 43169
rect 11701 43129 11713 43163
rect 11747 43160 11759 43163
rect 12618 43160 12624 43172
rect 11747 43132 12624 43160
rect 11747 43129 11759 43132
rect 11701 43123 11759 43129
rect 12618 43120 12624 43132
rect 12676 43120 12682 43172
rect 12728 43160 12756 43200
rect 13446 43188 13452 43200
rect 13504 43188 13510 43240
rect 13633 43231 13691 43237
rect 13633 43197 13645 43231
rect 13679 43197 13691 43231
rect 13633 43191 13691 43197
rect 14737 43231 14795 43237
rect 14737 43197 14749 43231
rect 14783 43228 14795 43231
rect 14918 43228 14924 43240
rect 14783 43200 14924 43228
rect 14783 43197 14795 43200
rect 14737 43191 14795 43197
rect 13354 43160 13360 43172
rect 12728 43132 13360 43160
rect 13354 43120 13360 43132
rect 13412 43160 13418 43172
rect 13648 43160 13676 43191
rect 14918 43188 14924 43200
rect 14976 43188 14982 43240
rect 15654 43228 15660 43240
rect 15615 43200 15660 43228
rect 15654 43188 15660 43200
rect 15712 43188 15718 43240
rect 13412 43132 13676 43160
rect 15013 43163 15071 43169
rect 13412 43120 13418 43132
rect 15013 43129 15025 43163
rect 15059 43160 15071 43163
rect 15764 43160 15792 43259
rect 16758 43256 16764 43268
rect 16816 43256 16822 43308
rect 16853 43299 16911 43305
rect 16853 43265 16865 43299
rect 16899 43296 16911 43299
rect 16942 43296 16948 43308
rect 16899 43268 16948 43296
rect 16899 43265 16911 43268
rect 16853 43259 16911 43265
rect 16942 43256 16948 43268
rect 17000 43256 17006 43308
rect 17034 43256 17040 43308
rect 17092 43296 17098 43308
rect 17512 43305 17540 43336
rect 17954 43324 17960 43336
rect 18012 43324 18018 43376
rect 18892 43364 18920 43404
rect 18969 43401 18981 43435
rect 19015 43432 19027 43435
rect 19242 43432 19248 43444
rect 19015 43404 19248 43432
rect 19015 43401 19027 43404
rect 18969 43395 19027 43401
rect 19242 43392 19248 43404
rect 19300 43392 19306 43444
rect 21542 43392 21548 43444
rect 21600 43432 21606 43444
rect 22465 43435 22523 43441
rect 22465 43432 22477 43435
rect 21600 43404 22477 43432
rect 21600 43392 21606 43404
rect 22465 43401 22477 43404
rect 22511 43401 22523 43435
rect 22465 43395 22523 43401
rect 23569 43435 23627 43441
rect 23569 43401 23581 43435
rect 23615 43432 23627 43435
rect 28074 43432 28080 43444
rect 23615 43404 27660 43432
rect 28035 43404 28080 43432
rect 23615 43401 23627 43404
rect 23569 43395 23627 43401
rect 20622 43364 20628 43376
rect 18892 43336 20628 43364
rect 17405 43299 17463 43305
rect 17405 43296 17417 43299
rect 17092 43268 17417 43296
rect 17092 43256 17098 43268
rect 17405 43265 17417 43268
rect 17451 43265 17463 43299
rect 17405 43259 17463 43265
rect 17497 43299 17555 43305
rect 17497 43265 17509 43299
rect 17543 43265 17555 43299
rect 17678 43296 17684 43308
rect 17639 43268 17684 43296
rect 17497 43259 17555 43265
rect 17678 43256 17684 43268
rect 17736 43256 17742 43308
rect 18322 43296 18328 43308
rect 18283 43268 18328 43296
rect 18322 43256 18328 43268
rect 18380 43256 18386 43308
rect 18506 43296 18512 43308
rect 18467 43268 18512 43296
rect 18506 43256 18512 43268
rect 18564 43256 18570 43308
rect 18620 43299 18678 43305
rect 18620 43296 18632 43299
rect 18616 43265 18632 43296
rect 18666 43265 18678 43299
rect 18713 43299 18771 43305
rect 18713 43296 18725 43299
rect 18616 43259 18678 43265
rect 18708 43265 18725 43296
rect 18759 43286 18771 43299
rect 18759 43265 18782 43286
rect 17862 43228 17868 43240
rect 17823 43200 17868 43228
rect 17862 43188 17868 43200
rect 17920 43188 17926 43240
rect 18616 43172 18644 43259
rect 18708 43258 18782 43265
rect 18754 43228 18782 43258
rect 18892 43228 18920 43336
rect 20622 43324 20628 43336
rect 20680 43324 20686 43376
rect 20806 43324 20812 43376
rect 20864 43364 20870 43376
rect 20901 43367 20959 43373
rect 20901 43364 20913 43367
rect 20864 43336 20913 43364
rect 20864 43324 20870 43336
rect 20901 43333 20913 43336
rect 20947 43364 20959 43367
rect 23750 43364 23756 43376
rect 20947 43336 22140 43364
rect 20947 43333 20959 43336
rect 20901 43327 20959 43333
rect 19797 43299 19855 43305
rect 19797 43265 19809 43299
rect 19843 43296 19855 43299
rect 20533 43299 20591 43305
rect 20533 43296 20545 43299
rect 19843 43268 20545 43296
rect 19843 43265 19855 43268
rect 19797 43259 19855 43265
rect 20533 43265 20545 43268
rect 20579 43265 20591 43299
rect 20714 43296 20720 43308
rect 20675 43268 20720 43296
rect 20533 43259 20591 43265
rect 20714 43256 20720 43268
rect 20772 43256 20778 43308
rect 20993 43299 21051 43305
rect 20993 43265 21005 43299
rect 21039 43265 21051 43299
rect 22002 43296 22008 43308
rect 21963 43268 22008 43296
rect 20993 43259 21051 43265
rect 18754 43200 18920 43228
rect 19426 43188 19432 43240
rect 19484 43228 19490 43240
rect 19613 43231 19671 43237
rect 19613 43228 19625 43231
rect 19484 43200 19625 43228
rect 19484 43188 19490 43200
rect 19613 43197 19625 43200
rect 19659 43197 19671 43231
rect 19613 43191 19671 43197
rect 19705 43231 19763 43237
rect 19705 43197 19717 43231
rect 19751 43197 19763 43231
rect 19705 43191 19763 43197
rect 19889 43231 19947 43237
rect 19889 43197 19901 43231
rect 19935 43228 19947 43231
rect 19978 43228 19984 43240
rect 19935 43200 19984 43228
rect 19935 43197 19947 43200
rect 19889 43191 19947 43197
rect 15838 43160 15844 43172
rect 15059 43132 15844 43160
rect 15059 43129 15071 43132
rect 15013 43123 15071 43129
rect 15838 43120 15844 43132
rect 15896 43120 15902 43172
rect 16117 43163 16175 43169
rect 16117 43129 16129 43163
rect 16163 43160 16175 43163
rect 17954 43160 17960 43172
rect 16163 43132 17960 43160
rect 16163 43129 16175 43132
rect 16117 43123 16175 43129
rect 17954 43120 17960 43132
rect 18012 43120 18018 43172
rect 18598 43120 18604 43172
rect 18656 43120 18662 43172
rect 19720 43160 19748 43191
rect 19978 43188 19984 43200
rect 20036 43188 20042 43240
rect 20346 43188 20352 43240
rect 20404 43228 20410 43240
rect 21008 43228 21036 43259
rect 22002 43256 22008 43268
rect 22060 43256 22066 43308
rect 22112 43305 22140 43336
rect 23124 43336 23756 43364
rect 23124 43305 23152 43336
rect 23750 43324 23756 43336
rect 23808 43324 23814 43376
rect 24762 43364 24768 43376
rect 24412 43336 24768 43364
rect 22097 43299 22155 43305
rect 22097 43265 22109 43299
rect 22143 43265 22155 43299
rect 22097 43259 22155 43265
rect 23109 43299 23167 43305
rect 23109 43265 23121 43299
rect 23155 43265 23167 43299
rect 23382 43296 23388 43308
rect 23343 43268 23388 43296
rect 23109 43259 23167 43265
rect 23382 43256 23388 43268
rect 23440 43256 23446 43308
rect 24026 43296 24032 43308
rect 23987 43268 24032 43296
rect 24026 43256 24032 43268
rect 24084 43256 24090 43308
rect 24412 43305 24440 43336
rect 24762 43324 24768 43336
rect 24820 43324 24826 43376
rect 26176 43367 26234 43373
rect 26176 43333 26188 43367
rect 26222 43364 26234 43367
rect 27246 43364 27252 43376
rect 26222 43336 27252 43364
rect 26222 43333 26234 43336
rect 26176 43327 26234 43333
rect 27246 43324 27252 43336
rect 27304 43324 27310 43376
rect 27632 43364 27660 43404
rect 28074 43392 28080 43404
rect 28132 43392 28138 43444
rect 28994 43392 29000 43444
rect 29052 43432 29058 43444
rect 29089 43435 29147 43441
rect 29089 43432 29101 43435
rect 29052 43404 29101 43432
rect 29052 43392 29058 43404
rect 29089 43401 29101 43404
rect 29135 43432 29147 43435
rect 29178 43432 29184 43444
rect 29135 43404 29184 43432
rect 29135 43401 29147 43404
rect 29089 43395 29147 43401
rect 29178 43392 29184 43404
rect 29236 43392 29242 43444
rect 33318 43432 33324 43444
rect 29288 43404 33324 43432
rect 29288 43364 29316 43404
rect 33318 43392 33324 43404
rect 33376 43392 33382 43444
rect 34514 43392 34520 43444
rect 34572 43432 34578 43444
rect 35437 43435 35495 43441
rect 35437 43432 35449 43435
rect 34572 43404 35449 43432
rect 34572 43392 34578 43404
rect 35437 43401 35449 43404
rect 35483 43401 35495 43435
rect 35437 43395 35495 43401
rect 35894 43392 35900 43444
rect 35952 43432 35958 43444
rect 35989 43435 36047 43441
rect 35989 43432 36001 43435
rect 35952 43404 36001 43432
rect 35952 43392 35958 43404
rect 35989 43401 36001 43404
rect 36035 43401 36047 43435
rect 35989 43395 36047 43401
rect 30374 43364 30380 43376
rect 27632 43336 29316 43364
rect 30335 43336 30380 43364
rect 30374 43324 30380 43336
rect 30432 43324 30438 43376
rect 32030 43324 32036 43376
rect 32088 43364 32094 43376
rect 32088 43336 33640 43364
rect 32088 43324 32094 43336
rect 24121 43299 24179 43305
rect 24121 43265 24133 43299
rect 24167 43265 24179 43299
rect 24232 43299 24290 43305
rect 24232 43296 24244 43299
rect 24121 43259 24179 43265
rect 24228 43265 24244 43296
rect 24278 43265 24290 43299
rect 24228 43259 24290 43265
rect 24397 43299 24455 43305
rect 24397 43265 24409 43299
rect 24443 43265 24455 43299
rect 24397 43259 24455 43265
rect 20404 43200 21036 43228
rect 20404 43188 20410 43200
rect 20073 43163 20131 43169
rect 19720 43132 20024 43160
rect 19996 43104 20024 43132
rect 20073 43129 20085 43163
rect 20119 43160 20131 43163
rect 23201 43163 23259 43169
rect 23201 43160 23213 43163
rect 20119 43132 23213 43160
rect 20119 43129 20131 43132
rect 20073 43123 20131 43129
rect 23201 43129 23213 43132
rect 23247 43129 23259 43163
rect 24136 43160 24164 43259
rect 24228 43228 24256 43259
rect 26326 43256 26332 43308
rect 26384 43256 26390 43308
rect 26421 43299 26479 43305
rect 26421 43265 26433 43299
rect 26467 43296 26479 43299
rect 27062 43296 27068 43308
rect 26467 43268 27068 43296
rect 26467 43265 26479 43268
rect 26421 43259 26479 43265
rect 27062 43256 27068 43268
rect 27120 43256 27126 43308
rect 33318 43296 33324 43308
rect 33376 43305 33382 43308
rect 33612 43305 33640 43336
rect 33686 43324 33692 43376
rect 33744 43364 33750 43376
rect 34302 43367 34360 43373
rect 34302 43364 34314 43367
rect 33744 43336 34314 43364
rect 33744 43324 33750 43336
rect 34302 43333 34314 43336
rect 34348 43333 34360 43367
rect 34302 43327 34360 43333
rect 35526 43324 35532 43376
rect 35584 43364 35590 43376
rect 35584 43336 36400 43364
rect 35584 43324 35590 43336
rect 33288 43268 33324 43296
rect 33318 43256 33324 43268
rect 33376 43259 33388 43305
rect 33597 43299 33655 43305
rect 33597 43265 33609 43299
rect 33643 43296 33655 43299
rect 34057 43299 34115 43305
rect 34057 43296 34069 43299
rect 33643 43268 34069 43296
rect 33643 43265 33655 43268
rect 33597 43259 33655 43265
rect 34057 43265 34069 43268
rect 34103 43265 34115 43299
rect 34057 43259 34115 43265
rect 33376 43256 33382 43259
rect 35618 43256 35624 43308
rect 35676 43296 35682 43308
rect 36372 43305 36400 43336
rect 36265 43299 36323 43305
rect 36265 43296 36277 43299
rect 35676 43268 36277 43296
rect 35676 43256 35682 43268
rect 36265 43265 36277 43268
rect 36311 43265 36323 43299
rect 36265 43259 36323 43265
rect 36357 43299 36415 43305
rect 36357 43265 36369 43299
rect 36403 43265 36415 43299
rect 36357 43259 36415 43265
rect 37737 43299 37795 43305
rect 37737 43265 37749 43299
rect 37783 43296 37795 43299
rect 37826 43296 37832 43308
rect 37783 43268 37832 43296
rect 37783 43265 37795 43268
rect 37737 43259 37795 43265
rect 37826 43256 37832 43268
rect 37884 43256 37890 43308
rect 37921 43299 37979 43305
rect 37921 43265 37933 43299
rect 37967 43296 37979 43299
rect 38286 43296 38292 43308
rect 37967 43268 38292 43296
rect 37967 43265 37979 43268
rect 37921 43259 37979 43265
rect 38286 43256 38292 43268
rect 38344 43256 38350 43308
rect 38378 43256 38384 43308
rect 38436 43296 38442 43308
rect 38436 43268 38481 43296
rect 38436 43256 38442 43268
rect 38562 43256 38568 43308
rect 38620 43296 38626 43308
rect 38620 43268 38665 43296
rect 38620 43256 38626 43268
rect 24486 43228 24492 43240
rect 24228 43200 24492 43228
rect 24486 43188 24492 43200
rect 24544 43188 24550 43240
rect 26344 43228 26372 43256
rect 26970 43228 26976 43240
rect 26344 43200 26976 43228
rect 26970 43188 26976 43200
rect 27028 43188 27034 43240
rect 35986 43188 35992 43240
rect 36044 43228 36050 43240
rect 36173 43231 36231 43237
rect 36173 43228 36185 43231
rect 36044 43200 36185 43228
rect 36044 43188 36050 43200
rect 36173 43197 36185 43200
rect 36219 43197 36231 43231
rect 36173 43191 36231 43197
rect 36449 43231 36507 43237
rect 36449 43197 36461 43231
rect 36495 43228 36507 43231
rect 36722 43228 36728 43240
rect 36495 43200 36728 43228
rect 36495 43197 36507 43200
rect 36449 43191 36507 43197
rect 36722 43188 36728 43200
rect 36780 43188 36786 43240
rect 24394 43160 24400 43172
rect 24136 43132 24400 43160
rect 23201 43123 23259 43129
rect 24394 43120 24400 43132
rect 24452 43120 24458 43172
rect 24581 43163 24639 43169
rect 24581 43129 24593 43163
rect 24627 43160 24639 43163
rect 35894 43160 35900 43172
rect 24627 43132 25544 43160
rect 24627 43129 24639 43132
rect 24581 43123 24639 43129
rect 12253 43095 12311 43101
rect 12253 43061 12265 43095
rect 12299 43092 12311 43095
rect 14182 43092 14188 43104
rect 12299 43064 14188 43092
rect 12299 43061 12311 43064
rect 12253 43055 12311 43061
rect 14182 43052 14188 43064
rect 14240 43052 14246 43104
rect 16666 43052 16672 43104
rect 16724 43092 16730 43104
rect 16761 43095 16819 43101
rect 16761 43092 16773 43095
rect 16724 43064 16773 43092
rect 16724 43052 16730 43064
rect 16761 43061 16773 43064
rect 16807 43061 16819 43095
rect 16761 43055 16819 43061
rect 19978 43052 19984 43104
rect 20036 43052 20042 43104
rect 21821 43095 21879 43101
rect 21821 43061 21833 43095
rect 21867 43092 21879 43095
rect 21910 43092 21916 43104
rect 21867 43064 21916 43092
rect 21867 43061 21879 43064
rect 21821 43055 21879 43061
rect 21910 43052 21916 43064
rect 21968 43052 21974 43104
rect 25041 43095 25099 43101
rect 25041 43061 25053 43095
rect 25087 43092 25099 43095
rect 25406 43092 25412 43104
rect 25087 43064 25412 43092
rect 25087 43061 25099 43064
rect 25041 43055 25099 43061
rect 25406 43052 25412 43064
rect 25464 43052 25470 43104
rect 25516 43092 25544 43132
rect 26896 43132 32720 43160
rect 26896 43092 26924 43132
rect 27614 43092 27620 43104
rect 25516 43064 26924 43092
rect 27575 43064 27620 43092
rect 27614 43052 27620 43064
rect 27672 43052 27678 43104
rect 30834 43092 30840 43104
rect 30795 43064 30840 43092
rect 30834 43052 30840 43064
rect 30892 43092 30898 43104
rect 31389 43095 31447 43101
rect 31389 43092 31401 43095
rect 30892 43064 31401 43092
rect 30892 43052 30898 43064
rect 31389 43061 31401 43064
rect 31435 43061 31447 43095
rect 32214 43092 32220 43104
rect 32175 43064 32220 43092
rect 31389 43055 31447 43061
rect 32214 43052 32220 43064
rect 32272 43052 32278 43104
rect 32692 43092 32720 43132
rect 35360 43132 35900 43160
rect 35158 43092 35164 43104
rect 32692 43064 35164 43092
rect 35158 43052 35164 43064
rect 35216 43092 35222 43104
rect 35360 43092 35388 43132
rect 35894 43120 35900 43132
rect 35952 43160 35958 43172
rect 36630 43160 36636 43172
rect 35952 43132 36636 43160
rect 35952 43120 35958 43132
rect 36630 43120 36636 43132
rect 36688 43120 36694 43172
rect 39942 43160 39948 43172
rect 39132 43132 39948 43160
rect 39132 43104 39160 43132
rect 39942 43120 39948 43132
rect 40000 43160 40006 43172
rect 40129 43163 40187 43169
rect 40129 43160 40141 43163
rect 40000 43132 40141 43160
rect 40000 43120 40006 43132
rect 40129 43129 40141 43132
rect 40175 43129 40187 43163
rect 40129 43123 40187 43129
rect 35216 43064 35388 43092
rect 37829 43095 37887 43101
rect 35216 43052 35222 43064
rect 37829 43061 37841 43095
rect 37875 43092 37887 43095
rect 38010 43092 38016 43104
rect 37875 43064 38016 43092
rect 37875 43061 37887 43064
rect 37829 43055 37887 43061
rect 38010 43052 38016 43064
rect 38068 43052 38074 43104
rect 38286 43052 38292 43104
rect 38344 43092 38350 43104
rect 38473 43095 38531 43101
rect 38473 43092 38485 43095
rect 38344 43064 38485 43092
rect 38344 43052 38350 43064
rect 38473 43061 38485 43064
rect 38519 43061 38531 43095
rect 39114 43092 39120 43104
rect 39075 43064 39120 43092
rect 38473 43055 38531 43061
rect 39114 43052 39120 43064
rect 39172 43052 39178 43104
rect 39669 43095 39727 43101
rect 39669 43061 39681 43095
rect 39715 43092 39727 43095
rect 40218 43092 40224 43104
rect 39715 43064 40224 43092
rect 39715 43061 39727 43064
rect 39669 43055 39727 43061
rect 40218 43052 40224 43064
rect 40276 43052 40282 43104
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 10137 42891 10195 42897
rect 10137 42857 10149 42891
rect 10183 42888 10195 42891
rect 10689 42891 10747 42897
rect 10689 42888 10701 42891
rect 10183 42860 10701 42888
rect 10183 42857 10195 42860
rect 10137 42851 10195 42857
rect 10689 42857 10701 42860
rect 10735 42888 10747 42891
rect 10962 42888 10968 42900
rect 10735 42860 10968 42888
rect 10735 42857 10747 42860
rect 10689 42851 10747 42857
rect 10962 42848 10968 42860
rect 11020 42848 11026 42900
rect 12805 42891 12863 42897
rect 12805 42857 12817 42891
rect 12851 42888 12863 42891
rect 13078 42888 13084 42900
rect 12851 42860 13084 42888
rect 12851 42857 12863 42860
rect 12805 42851 12863 42857
rect 13078 42848 13084 42860
rect 13136 42848 13142 42900
rect 15654 42848 15660 42900
rect 15712 42888 15718 42900
rect 15749 42891 15807 42897
rect 15749 42888 15761 42891
rect 15712 42860 15761 42888
rect 15712 42848 15718 42860
rect 15749 42857 15761 42860
rect 15795 42857 15807 42891
rect 15749 42851 15807 42857
rect 18049 42891 18107 42897
rect 18049 42857 18061 42891
rect 18095 42888 18107 42891
rect 18506 42888 18512 42900
rect 18095 42860 18512 42888
rect 18095 42857 18107 42860
rect 18049 42851 18107 42857
rect 18506 42848 18512 42860
rect 18564 42848 18570 42900
rect 19518 42848 19524 42900
rect 19576 42888 19582 42900
rect 19705 42891 19763 42897
rect 19705 42888 19717 42891
rect 19576 42860 19717 42888
rect 19576 42848 19582 42860
rect 19705 42857 19717 42860
rect 19751 42857 19763 42891
rect 19705 42851 19763 42857
rect 20441 42891 20499 42897
rect 20441 42857 20453 42891
rect 20487 42888 20499 42891
rect 20714 42888 20720 42900
rect 20487 42860 20720 42888
rect 20487 42857 20499 42860
rect 20441 42851 20499 42857
rect 12618 42780 12624 42832
rect 12676 42820 12682 42832
rect 16574 42820 16580 42832
rect 12676 42792 16580 42820
rect 12676 42780 12682 42792
rect 16574 42780 16580 42792
rect 16632 42780 16638 42832
rect 9582 42712 9588 42764
rect 9640 42752 9646 42764
rect 12345 42755 12403 42761
rect 12345 42752 12357 42755
rect 9640 42724 12357 42752
rect 9640 42712 9646 42724
rect 12345 42721 12357 42724
rect 12391 42752 12403 42755
rect 12391 42724 12756 42752
rect 12391 42721 12403 42724
rect 12345 42715 12403 42721
rect 1673 42687 1731 42693
rect 1673 42653 1685 42687
rect 1719 42684 1731 42687
rect 2225 42687 2283 42693
rect 2225 42684 2237 42687
rect 1719 42656 2237 42684
rect 1719 42653 1731 42656
rect 1673 42647 1731 42653
rect 2225 42653 2237 42656
rect 2271 42684 2283 42687
rect 2271 42656 6914 42684
rect 2271 42653 2283 42656
rect 2225 42647 2283 42653
rect 6886 42616 6914 42656
rect 10778 42644 10784 42696
rect 10836 42684 10842 42696
rect 11238 42684 11244 42696
rect 10836 42656 11244 42684
rect 10836 42644 10842 42656
rect 11238 42644 11244 42656
rect 11296 42684 11302 42696
rect 12250 42684 12256 42696
rect 11296 42656 12256 42684
rect 11296 42644 11302 42656
rect 12250 42644 12256 42656
rect 12308 42684 12314 42696
rect 12437 42687 12495 42693
rect 12437 42684 12449 42687
rect 12308 42656 12449 42684
rect 12308 42644 12314 42656
rect 12437 42653 12449 42656
rect 12483 42684 12495 42687
rect 12728 42684 12756 42724
rect 12894 42712 12900 42764
rect 12952 42752 12958 42764
rect 12952 42724 13492 42752
rect 12952 42712 12958 42724
rect 12986 42684 12992 42696
rect 12483 42656 12664 42684
rect 12728 42656 12992 42684
rect 12483 42653 12495 42656
rect 12437 42647 12495 42653
rect 12636 42616 12664 42656
rect 12986 42644 12992 42656
rect 13044 42644 13050 42696
rect 13464 42684 13492 42724
rect 13538 42712 13544 42764
rect 13596 42752 13602 42764
rect 15838 42752 15844 42764
rect 13596 42724 15700 42752
rect 15799 42724 15844 42752
rect 13596 42712 13602 42724
rect 14826 42684 14832 42696
rect 13464 42656 14832 42684
rect 14826 42644 14832 42656
rect 14884 42644 14890 42696
rect 15562 42684 15568 42696
rect 15523 42656 15568 42684
rect 15562 42644 15568 42656
rect 15620 42644 15626 42696
rect 15672 42684 15700 42724
rect 15838 42712 15844 42724
rect 15896 42712 15902 42764
rect 16758 42712 16764 42764
rect 16816 42712 16822 42764
rect 19720 42752 19748 42851
rect 20714 42848 20720 42860
rect 20772 42888 20778 42900
rect 21453 42891 21511 42897
rect 21453 42888 21465 42891
rect 20772 42860 21465 42888
rect 20772 42848 20778 42860
rect 21453 42857 21465 42860
rect 21499 42857 21511 42891
rect 21634 42888 21640 42900
rect 21595 42860 21640 42888
rect 21453 42851 21511 42857
rect 21634 42848 21640 42860
rect 21692 42848 21698 42900
rect 23198 42848 23204 42900
rect 23256 42888 23262 42900
rect 31478 42888 31484 42900
rect 23256 42860 31484 42888
rect 23256 42848 23262 42860
rect 31478 42848 31484 42860
rect 31536 42848 31542 42900
rect 33965 42891 34023 42897
rect 33965 42857 33977 42891
rect 34011 42888 34023 42891
rect 34054 42888 34060 42900
rect 34011 42860 34060 42888
rect 34011 42857 34023 42860
rect 33965 42851 34023 42857
rect 34054 42848 34060 42860
rect 34112 42848 34118 42900
rect 39942 42848 39948 42900
rect 40000 42888 40006 42900
rect 40405 42891 40463 42897
rect 40405 42888 40417 42891
rect 40000 42860 40417 42888
rect 40000 42848 40006 42860
rect 40405 42857 40417 42860
rect 40451 42857 40463 42891
rect 40405 42851 40463 42857
rect 26326 42820 26332 42832
rect 23584 42792 26332 42820
rect 20346 42752 20352 42764
rect 19720 42724 20352 42752
rect 20346 42712 20352 42724
rect 20404 42712 20410 42764
rect 21910 42752 21916 42764
rect 20640 42724 21916 42752
rect 16776 42684 16804 42712
rect 15672 42656 16804 42684
rect 16850 42644 16856 42696
rect 16908 42684 16914 42696
rect 16945 42687 17003 42693
rect 16945 42684 16957 42687
rect 16908 42656 16957 42684
rect 16908 42644 16914 42656
rect 16945 42653 16957 42656
rect 16991 42653 17003 42687
rect 17954 42684 17960 42696
rect 17915 42656 17960 42684
rect 16945 42647 17003 42653
rect 17954 42644 17960 42656
rect 18012 42644 18018 42696
rect 18138 42684 18144 42696
rect 18099 42656 18144 42684
rect 18138 42644 18144 42656
rect 18196 42644 18202 42696
rect 19334 42684 19340 42696
rect 19295 42656 19340 42684
rect 19334 42644 19340 42656
rect 19392 42644 19398 42696
rect 19429 42687 19487 42693
rect 19429 42653 19441 42687
rect 19475 42653 19487 42687
rect 19429 42647 19487 42653
rect 19521 42687 19579 42693
rect 19521 42653 19533 42687
rect 19567 42653 19579 42687
rect 19521 42647 19579 42653
rect 14918 42616 14924 42628
rect 6886 42588 12434 42616
rect 12636 42588 14924 42616
rect 1486 42548 1492 42560
rect 1447 42520 1492 42548
rect 1486 42508 1492 42520
rect 1544 42508 1550 42560
rect 9582 42548 9588 42560
rect 9543 42520 9588 42548
rect 9582 42508 9588 42520
rect 9640 42508 9646 42560
rect 10778 42508 10784 42560
rect 10836 42548 10842 42560
rect 11149 42551 11207 42557
rect 11149 42548 11161 42551
rect 10836 42520 11161 42548
rect 10836 42508 10842 42520
rect 11149 42517 11161 42520
rect 11195 42517 11207 42551
rect 11790 42548 11796 42560
rect 11751 42520 11796 42548
rect 11149 42511 11207 42517
rect 11790 42508 11796 42520
rect 11848 42508 11854 42560
rect 12406 42548 12434 42588
rect 14918 42576 14924 42588
rect 14976 42576 14982 42628
rect 16761 42619 16819 42625
rect 16761 42616 16773 42619
rect 15304 42588 16773 42616
rect 12894 42548 12900 42560
rect 12406 42520 12900 42548
rect 12894 42508 12900 42520
rect 12952 42508 12958 42560
rect 13814 42508 13820 42560
rect 13872 42548 13878 42560
rect 14369 42551 14427 42557
rect 14369 42548 14381 42551
rect 13872 42520 14381 42548
rect 13872 42508 13878 42520
rect 14369 42517 14381 42520
rect 14415 42548 14427 42551
rect 15304 42548 15332 42588
rect 16761 42585 16773 42588
rect 16807 42616 16819 42619
rect 16807 42588 16988 42616
rect 16807 42585 16819 42588
rect 16761 42579 16819 42585
rect 16960 42560 16988 42588
rect 17126 42576 17132 42628
rect 17184 42616 17190 42628
rect 18506 42616 18512 42628
rect 17184 42588 18512 42616
rect 17184 42576 17190 42588
rect 18506 42576 18512 42588
rect 18564 42616 18570 42628
rect 19444 42616 19472 42647
rect 18564 42588 19472 42616
rect 18564 42576 18570 42588
rect 14415 42520 15332 42548
rect 15381 42551 15439 42557
rect 14415 42517 14427 42520
rect 14369 42511 14427 42517
rect 15381 42517 15393 42551
rect 15427 42548 15439 42551
rect 15654 42548 15660 42560
rect 15427 42520 15660 42548
rect 15427 42517 15439 42520
rect 15381 42511 15439 42517
rect 15654 42508 15660 42520
rect 15712 42508 15718 42560
rect 16942 42508 16948 42560
rect 17000 42508 17006 42560
rect 17954 42508 17960 42560
rect 18012 42548 18018 42560
rect 18601 42551 18659 42557
rect 18601 42548 18613 42551
rect 18012 42520 18613 42548
rect 18012 42508 18018 42520
rect 18601 42517 18613 42520
rect 18647 42517 18659 42551
rect 18601 42511 18659 42517
rect 18782 42508 18788 42560
rect 18840 42548 18846 42560
rect 19536 42548 19564 42647
rect 20364 42616 20392 42712
rect 20640 42693 20668 42724
rect 21910 42712 21916 42724
rect 21968 42712 21974 42764
rect 22094 42712 22100 42764
rect 22152 42752 22158 42764
rect 23474 42752 23480 42764
rect 22152 42724 23480 42752
rect 22152 42712 22158 42724
rect 23474 42712 23480 42724
rect 23532 42712 23538 42764
rect 20625 42687 20683 42693
rect 20625 42653 20637 42687
rect 20671 42653 20683 42687
rect 20625 42647 20683 42653
rect 21269 42687 21327 42693
rect 21269 42653 21281 42687
rect 21315 42653 21327 42687
rect 21542 42684 21548 42696
rect 21503 42656 21548 42684
rect 21269 42647 21327 42653
rect 21284 42616 21312 42647
rect 21542 42644 21548 42656
rect 21600 42644 21606 42696
rect 21729 42687 21787 42693
rect 21729 42653 21741 42687
rect 21775 42684 21787 42687
rect 21818 42684 21824 42696
rect 21775 42656 21824 42684
rect 21775 42653 21787 42656
rect 21729 42647 21787 42653
rect 21818 42644 21824 42656
rect 21876 42644 21882 42696
rect 22002 42616 22008 42628
rect 20364 42588 21312 42616
rect 21963 42588 22008 42616
rect 22002 42576 22008 42588
rect 22060 42576 22066 42628
rect 22738 42616 22744 42628
rect 22699 42588 22744 42616
rect 22738 42576 22744 42588
rect 22796 42576 22802 42628
rect 22830 42576 22836 42628
rect 22888 42616 22894 42628
rect 22925 42619 22983 42625
rect 22925 42616 22937 42619
rect 22888 42588 22937 42616
rect 22888 42576 22894 42588
rect 22925 42585 22937 42588
rect 22971 42616 22983 42619
rect 23584 42616 23612 42792
rect 26326 42780 26332 42792
rect 26384 42780 26390 42832
rect 34606 42780 34612 42832
rect 34664 42820 34670 42832
rect 34664 42792 35020 42820
rect 34664 42780 34670 42792
rect 24026 42712 24032 42764
rect 24084 42712 24090 42764
rect 24486 42712 24492 42764
rect 24544 42752 24550 42764
rect 25501 42755 25559 42761
rect 24544 42724 24808 42752
rect 24544 42712 24550 42724
rect 23661 42687 23719 42693
rect 23661 42653 23673 42687
rect 23707 42684 23719 42687
rect 23750 42684 23756 42696
rect 23707 42656 23756 42684
rect 23707 42653 23719 42656
rect 23661 42647 23719 42653
rect 23750 42644 23756 42656
rect 23808 42644 23814 42696
rect 23845 42687 23903 42693
rect 23845 42653 23857 42687
rect 23891 42684 23903 42687
rect 24044 42684 24072 42712
rect 24581 42687 24639 42693
rect 24581 42684 24593 42687
rect 23891 42656 24593 42684
rect 23891 42653 23903 42656
rect 23845 42647 23903 42653
rect 24581 42653 24593 42656
rect 24627 42684 24639 42687
rect 24670 42684 24676 42696
rect 24627 42656 24676 42684
rect 24627 42653 24639 42656
rect 24581 42647 24639 42653
rect 24670 42644 24676 42656
rect 24728 42644 24734 42696
rect 24780 42693 24808 42724
rect 25501 42721 25513 42755
rect 25547 42752 25559 42755
rect 25774 42752 25780 42764
rect 25547 42724 25780 42752
rect 25547 42721 25559 42724
rect 25501 42715 25559 42721
rect 25774 42712 25780 42724
rect 25832 42712 25838 42764
rect 27062 42712 27068 42764
rect 27120 42752 27126 42764
rect 27341 42755 27399 42761
rect 27341 42752 27353 42755
rect 27120 42724 27353 42752
rect 27120 42712 27126 42724
rect 27341 42721 27353 42724
rect 27387 42721 27399 42755
rect 27341 42715 27399 42721
rect 29549 42755 29607 42761
rect 29549 42721 29561 42755
rect 29595 42752 29607 42755
rect 32030 42752 32036 42764
rect 29595 42724 32036 42752
rect 29595 42721 29607 42724
rect 29549 42715 29607 42721
rect 32030 42712 32036 42724
rect 32088 42752 32094 42764
rect 33321 42755 33379 42761
rect 33321 42752 33333 42755
rect 32088 42724 33333 42752
rect 32088 42712 32094 42724
rect 33321 42721 33333 42724
rect 33367 42721 33379 42755
rect 34422 42752 34428 42764
rect 33321 42715 33379 42721
rect 33796 42724 34428 42752
rect 33796 42696 33824 42724
rect 34422 42712 34428 42724
rect 34480 42712 34486 42764
rect 34698 42752 34704 42764
rect 34659 42724 34704 42752
rect 34698 42712 34704 42724
rect 34756 42712 34762 42764
rect 24765 42687 24823 42693
rect 24765 42653 24777 42687
rect 24811 42653 24823 42687
rect 24765 42647 24823 42653
rect 24854 42644 24860 42696
rect 24912 42684 24918 42696
rect 25317 42687 25375 42693
rect 24912 42656 24957 42684
rect 24912 42644 24918 42656
rect 25317 42653 25329 42687
rect 25363 42653 25375 42687
rect 25682 42684 25688 42696
rect 25643 42656 25688 42684
rect 25317 42647 25375 42653
rect 22971 42588 23612 42616
rect 22971 42585 22983 42588
rect 22925 42579 22983 42585
rect 24026 42576 24032 42628
rect 24084 42616 24090 42628
rect 25332 42616 25360 42647
rect 25682 42644 25688 42656
rect 25740 42644 25746 42696
rect 27617 42687 27675 42693
rect 27617 42684 27629 42687
rect 26620 42656 27629 42684
rect 26620 42616 26648 42656
rect 27617 42653 27629 42656
rect 27663 42653 27675 42687
rect 29822 42684 29828 42696
rect 29783 42656 29828 42684
rect 27617 42647 27675 42653
rect 29822 42644 29828 42656
rect 29880 42644 29886 42696
rect 33045 42687 33103 42693
rect 33045 42684 33057 42687
rect 30484 42656 33057 42684
rect 24084 42588 25360 42616
rect 25608 42588 26648 42616
rect 24084 42576 24090 42588
rect 18840 42520 19564 42548
rect 20809 42551 20867 42557
rect 18840 42508 18846 42520
rect 20809 42517 20821 42551
rect 20855 42548 20867 42551
rect 22186 42548 22192 42560
rect 20855 42520 22192 42548
rect 20855 42517 20867 42520
rect 20809 42511 20867 42517
rect 22186 42508 22192 42520
rect 22244 42508 22250 42560
rect 22554 42508 22560 42560
rect 22612 42548 22618 42560
rect 24397 42551 24455 42557
rect 22612 42520 22657 42548
rect 22612 42508 22618 42520
rect 24397 42517 24409 42551
rect 24443 42548 24455 42551
rect 24578 42548 24584 42560
rect 24443 42520 24584 42548
rect 24443 42517 24455 42520
rect 24397 42511 24455 42517
rect 24578 42508 24584 42520
rect 24636 42508 24642 42560
rect 24854 42508 24860 42560
rect 24912 42548 24918 42560
rect 25608 42557 25636 42588
rect 25409 42551 25467 42557
rect 25409 42548 25421 42551
rect 24912 42520 25421 42548
rect 24912 42508 24918 42520
rect 25409 42517 25421 42520
rect 25455 42517 25467 42551
rect 25409 42511 25467 42517
rect 25593 42551 25651 42557
rect 25593 42517 25605 42551
rect 25639 42517 25651 42551
rect 25593 42511 25651 42517
rect 26050 42508 26056 42560
rect 26108 42548 26114 42560
rect 26145 42551 26203 42557
rect 26145 42548 26157 42551
rect 26108 42520 26157 42548
rect 26108 42508 26114 42520
rect 26145 42517 26157 42520
rect 26191 42517 26203 42551
rect 26694 42548 26700 42560
rect 26655 42520 26700 42548
rect 26145 42511 26203 42517
rect 26694 42508 26700 42520
rect 26752 42508 26758 42560
rect 28626 42508 28632 42560
rect 28684 42548 28690 42560
rect 28721 42551 28779 42557
rect 28721 42548 28733 42551
rect 28684 42520 28733 42548
rect 28684 42508 28690 42520
rect 28721 42517 28733 42520
rect 28767 42517 28779 42551
rect 28721 42511 28779 42517
rect 28902 42508 28908 42560
rect 28960 42548 28966 42560
rect 30484 42548 30512 42656
rect 33045 42653 33057 42656
rect 33091 42653 33103 42687
rect 33045 42647 33103 42653
rect 33778 42644 33784 42696
rect 33836 42644 33842 42696
rect 33870 42644 33876 42696
rect 33928 42684 33934 42696
rect 34885 42687 34943 42693
rect 34885 42684 34897 42687
rect 33928 42656 34897 42684
rect 33928 42644 33934 42656
rect 34885 42653 34897 42656
rect 34931 42653 34943 42687
rect 34992 42684 35020 42792
rect 35069 42755 35127 42761
rect 35069 42721 35081 42755
rect 35115 42752 35127 42755
rect 37001 42755 37059 42761
rect 37001 42752 37013 42755
rect 35115 42724 37013 42752
rect 35115 42721 35127 42724
rect 35069 42715 35127 42721
rect 37001 42721 37013 42724
rect 37047 42721 37059 42755
rect 37274 42752 37280 42764
rect 37235 42724 37280 42752
rect 37001 42715 37059 42721
rect 37274 42712 37280 42724
rect 37332 42752 37338 42764
rect 38105 42755 38163 42761
rect 38105 42752 38117 42755
rect 37332 42724 38117 42752
rect 37332 42712 37338 42724
rect 38105 42721 38117 42724
rect 38151 42721 38163 42755
rect 38286 42752 38292 42764
rect 38247 42724 38292 42752
rect 38105 42715 38163 42721
rect 38286 42712 38292 42724
rect 38344 42712 38350 42764
rect 35158 42684 35164 42696
rect 34992 42656 35164 42684
rect 34885 42647 34943 42653
rect 35158 42644 35164 42656
rect 35216 42644 35222 42696
rect 35253 42687 35311 42693
rect 35253 42653 35265 42687
rect 35299 42653 35311 42687
rect 35434 42684 35440 42696
rect 35395 42656 35440 42684
rect 35253 42647 35311 42653
rect 31386 42576 31392 42628
rect 31444 42616 31450 42628
rect 33796 42616 33824 42644
rect 34149 42619 34207 42625
rect 34149 42616 34161 42619
rect 31444 42588 31892 42616
rect 33796 42588 34161 42616
rect 31444 42576 31450 42588
rect 28960 42520 30512 42548
rect 28960 42508 28966 42520
rect 31018 42508 31024 42560
rect 31076 42548 31082 42560
rect 31113 42551 31171 42557
rect 31113 42548 31125 42551
rect 31076 42520 31125 42548
rect 31076 42508 31082 42520
rect 31113 42517 31125 42520
rect 31159 42517 31171 42551
rect 31754 42548 31760 42560
rect 31715 42520 31760 42548
rect 31113 42511 31171 42517
rect 31754 42508 31760 42520
rect 31812 42508 31818 42560
rect 31864 42548 31892 42588
rect 34149 42585 34161 42588
rect 34195 42585 34207 42619
rect 34149 42579 34207 42585
rect 34238 42576 34244 42628
rect 34296 42616 34302 42628
rect 35268 42616 35296 42647
rect 35434 42644 35440 42656
rect 35492 42644 35498 42696
rect 35897 42687 35955 42693
rect 35897 42653 35909 42687
rect 35943 42684 35955 42687
rect 35986 42684 35992 42696
rect 35943 42656 35992 42684
rect 35943 42653 35955 42656
rect 35897 42647 35955 42653
rect 35986 42644 35992 42656
rect 36044 42644 36050 42696
rect 36262 42684 36268 42696
rect 36223 42656 36268 42684
rect 36262 42644 36268 42656
rect 36320 42644 36326 42696
rect 36357 42687 36415 42693
rect 36357 42653 36369 42687
rect 36403 42653 36415 42687
rect 36357 42647 36415 42653
rect 37369 42687 37427 42693
rect 37369 42653 37381 42687
rect 37415 42684 37427 42687
rect 37458 42684 37464 42696
rect 37415 42656 37464 42684
rect 37415 42653 37427 42656
rect 37369 42647 37427 42653
rect 34296 42588 35296 42616
rect 34296 42576 34302 42588
rect 35342 42576 35348 42628
rect 35400 42616 35406 42628
rect 36372 42616 36400 42647
rect 37458 42644 37464 42656
rect 37516 42684 37522 42696
rect 38010 42684 38016 42696
rect 37516 42656 38016 42684
rect 37516 42644 37522 42656
rect 38010 42644 38016 42656
rect 38068 42644 38074 42696
rect 47489 42687 47547 42693
rect 47489 42653 47501 42687
rect 47535 42684 47547 42687
rect 48130 42684 48136 42696
rect 47535 42656 48136 42684
rect 47535 42653 47547 42656
rect 47489 42647 47547 42653
rect 48130 42644 48136 42656
rect 48188 42644 48194 42696
rect 35400 42588 36400 42616
rect 35400 42576 35406 42588
rect 37182 42576 37188 42628
rect 37240 42616 37246 42628
rect 38749 42619 38807 42625
rect 38749 42616 38761 42619
rect 37240 42588 38761 42616
rect 37240 42576 37246 42588
rect 38749 42585 38761 42588
rect 38795 42585 38807 42619
rect 38749 42579 38807 42585
rect 33781 42551 33839 42557
rect 33781 42548 33793 42551
rect 31864 42520 33793 42548
rect 33781 42517 33793 42520
rect 33827 42517 33839 42551
rect 33781 42511 33839 42517
rect 33949 42551 34007 42557
rect 33949 42517 33961 42551
rect 33995 42548 34007 42551
rect 35618 42548 35624 42560
rect 33995 42520 35624 42548
rect 33995 42517 34007 42520
rect 33949 42511 34007 42517
rect 35618 42508 35624 42520
rect 35676 42508 35682 42560
rect 35894 42508 35900 42560
rect 35952 42548 35958 42560
rect 35989 42551 36047 42557
rect 35989 42548 36001 42551
rect 35952 42520 36001 42548
rect 35952 42508 35958 42520
rect 35989 42517 36001 42520
rect 36035 42517 36047 42551
rect 35989 42511 36047 42517
rect 36173 42551 36231 42557
rect 36173 42517 36185 42551
rect 36219 42548 36231 42551
rect 36446 42548 36452 42560
rect 36219 42520 36452 42548
rect 36219 42517 36231 42520
rect 36173 42511 36231 42517
rect 36446 42508 36452 42520
rect 36504 42508 36510 42560
rect 36538 42508 36544 42560
rect 36596 42548 36602 42560
rect 36596 42520 36641 42548
rect 36596 42508 36602 42520
rect 37734 42508 37740 42560
rect 37792 42548 37798 42560
rect 38289 42551 38347 42557
rect 38289 42548 38301 42551
rect 37792 42520 38301 42548
rect 37792 42508 37798 42520
rect 38289 42517 38301 42520
rect 38335 42517 38347 42551
rect 38289 42511 38347 42517
rect 38562 42508 38568 42560
rect 38620 42548 38626 42560
rect 39945 42551 40003 42557
rect 39945 42548 39957 42551
rect 38620 42520 39957 42548
rect 38620 42508 38626 42520
rect 39945 42517 39957 42520
rect 39991 42548 40003 42551
rect 40034 42548 40040 42560
rect 39991 42520 40040 42548
rect 39991 42517 40003 42520
rect 39945 42511 40003 42517
rect 40034 42508 40040 42520
rect 40092 42508 40098 42560
rect 47946 42548 47952 42560
rect 47907 42520 47952 42548
rect 47946 42508 47952 42520
rect 48004 42508 48010 42560
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 11054 42304 11060 42356
rect 11112 42344 11118 42356
rect 11701 42347 11759 42353
rect 11701 42344 11713 42347
rect 11112 42316 11713 42344
rect 11112 42304 11118 42316
rect 11701 42313 11713 42316
rect 11747 42344 11759 42347
rect 12066 42344 12072 42356
rect 11747 42316 12072 42344
rect 11747 42313 11759 42316
rect 11701 42307 11759 42313
rect 12066 42304 12072 42316
rect 12124 42304 12130 42356
rect 12345 42347 12403 42353
rect 12345 42313 12357 42347
rect 12391 42344 12403 42347
rect 12434 42344 12440 42356
rect 12391 42316 12440 42344
rect 12391 42313 12403 42316
rect 12345 42307 12403 42313
rect 12434 42304 12440 42316
rect 12492 42304 12498 42356
rect 13173 42347 13231 42353
rect 13173 42313 13185 42347
rect 13219 42344 13231 42347
rect 13446 42344 13452 42356
rect 13219 42316 13452 42344
rect 13219 42313 13231 42316
rect 13173 42307 13231 42313
rect 13446 42304 13452 42316
rect 13504 42304 13510 42356
rect 14090 42344 14096 42356
rect 14051 42316 14096 42344
rect 14090 42304 14096 42316
rect 14148 42304 14154 42356
rect 15194 42344 15200 42356
rect 15155 42316 15200 42344
rect 15194 42304 15200 42316
rect 15252 42344 15258 42356
rect 17313 42347 17371 42353
rect 17313 42344 17325 42347
rect 15252 42316 17325 42344
rect 15252 42304 15258 42316
rect 17313 42313 17325 42316
rect 17359 42344 17371 42347
rect 20530 42344 20536 42356
rect 17359 42316 20392 42344
rect 20491 42316 20536 42344
rect 17359 42313 17371 42316
rect 17313 42307 17371 42313
rect 12452 42276 12480 42304
rect 14553 42279 14611 42285
rect 14553 42276 14565 42279
rect 12452 42248 14565 42276
rect 14553 42245 14565 42248
rect 14599 42276 14611 42279
rect 18138 42276 18144 42288
rect 14599 42248 18144 42276
rect 14599 42245 14611 42248
rect 14553 42239 14611 42245
rect 18138 42236 18144 42248
rect 18196 42276 18202 42288
rect 19978 42276 19984 42288
rect 18196 42248 19984 42276
rect 18196 42236 18202 42248
rect 19978 42236 19984 42248
rect 20036 42236 20042 42288
rect 20364 42276 20392 42316
rect 20530 42304 20536 42316
rect 20588 42304 20594 42356
rect 21174 42344 21180 42356
rect 21135 42316 21180 42344
rect 21174 42304 21180 42316
rect 21232 42304 21238 42356
rect 21818 42344 21824 42356
rect 21779 42316 21824 42344
rect 21818 42304 21824 42316
rect 21876 42304 21882 42356
rect 24026 42344 24032 42356
rect 23987 42316 24032 42344
rect 24026 42304 24032 42316
rect 24084 42304 24090 42356
rect 24854 42344 24860 42356
rect 24815 42316 24860 42344
rect 24854 42304 24860 42316
rect 24912 42304 24918 42356
rect 24964 42316 29960 42344
rect 20990 42276 20996 42288
rect 20364 42248 20996 42276
rect 20990 42236 20996 42248
rect 21048 42276 21054 42288
rect 21726 42276 21732 42288
rect 21048 42248 21732 42276
rect 21048 42236 21054 42248
rect 21726 42236 21732 42248
rect 21784 42236 21790 42288
rect 22480 42248 23152 42276
rect 22480 42220 22508 42248
rect 12250 42168 12256 42220
rect 12308 42208 12314 42220
rect 12805 42211 12863 42217
rect 12805 42208 12817 42211
rect 12308 42180 12817 42208
rect 12308 42168 12314 42180
rect 12805 42177 12817 42180
rect 12851 42177 12863 42211
rect 12986 42208 12992 42220
rect 12947 42180 12992 42208
rect 12805 42171 12863 42177
rect 12986 42168 12992 42180
rect 13044 42168 13050 42220
rect 15654 42208 15660 42220
rect 15615 42180 15660 42208
rect 15654 42168 15660 42180
rect 15712 42168 15718 42220
rect 16025 42211 16083 42217
rect 16025 42177 16037 42211
rect 16071 42208 16083 42211
rect 16666 42208 16672 42220
rect 16071 42180 16672 42208
rect 16071 42177 16083 42180
rect 16025 42171 16083 42177
rect 16666 42168 16672 42180
rect 16724 42168 16730 42220
rect 16853 42211 16911 42217
rect 16853 42177 16865 42211
rect 16899 42208 16911 42211
rect 17126 42208 17132 42220
rect 16899 42180 17132 42208
rect 16899 42177 16911 42180
rect 16853 42171 16911 42177
rect 17126 42168 17132 42180
rect 17184 42168 17190 42220
rect 17954 42208 17960 42220
rect 17915 42180 17960 42208
rect 17954 42168 17960 42180
rect 18012 42168 18018 42220
rect 18601 42211 18659 42217
rect 18601 42177 18613 42211
rect 18647 42208 18659 42211
rect 19334 42208 19340 42220
rect 18647 42180 19340 42208
rect 18647 42177 18659 42180
rect 18601 42171 18659 42177
rect 19334 42168 19340 42180
rect 19392 42168 19398 42220
rect 20898 42168 20904 42220
rect 20956 42208 20962 42220
rect 21085 42211 21143 42217
rect 21085 42208 21097 42211
rect 20956 42180 21097 42208
rect 20956 42168 20962 42180
rect 21085 42177 21097 42180
rect 21131 42208 21143 42211
rect 21174 42208 21180 42220
rect 21131 42180 21180 42208
rect 21131 42177 21143 42180
rect 21085 42171 21143 42177
rect 21174 42168 21180 42180
rect 21232 42168 21238 42220
rect 21269 42211 21327 42217
rect 21269 42177 21281 42211
rect 21315 42208 21327 42211
rect 21450 42208 21456 42220
rect 21315 42180 21456 42208
rect 21315 42177 21327 42180
rect 21269 42171 21327 42177
rect 21450 42168 21456 42180
rect 21508 42168 21514 42220
rect 21542 42168 21548 42220
rect 21600 42208 21606 42220
rect 22002 42208 22008 42220
rect 21600 42180 22008 42208
rect 21600 42168 21606 42180
rect 22002 42168 22008 42180
rect 22060 42168 22066 42220
rect 22278 42208 22284 42220
rect 22239 42180 22284 42208
rect 22278 42168 22284 42180
rect 22336 42168 22342 42220
rect 22462 42208 22468 42220
rect 22423 42180 22468 42208
rect 22462 42168 22468 42180
rect 22520 42168 22526 42220
rect 22554 42168 22560 42220
rect 22612 42208 22618 42220
rect 23124 42217 23152 42248
rect 23290 42236 23296 42288
rect 23348 42276 23354 42288
rect 24964 42276 24992 42316
rect 23348 42248 24992 42276
rect 29932 42276 29960 42316
rect 30466 42304 30472 42356
rect 30524 42344 30530 42356
rect 30650 42344 30656 42356
rect 30524 42316 30656 42344
rect 30524 42304 30530 42316
rect 30650 42304 30656 42316
rect 30708 42304 30714 42356
rect 31754 42344 31760 42356
rect 31128 42316 31760 42344
rect 31128 42276 31156 42316
rect 31754 42304 31760 42316
rect 31812 42304 31818 42356
rect 35342 42344 35348 42356
rect 35303 42316 35348 42344
rect 35342 42304 35348 42316
rect 35400 42304 35406 42356
rect 35437 42347 35495 42353
rect 35437 42313 35449 42347
rect 35483 42344 35495 42347
rect 35526 42344 35532 42356
rect 35483 42316 35532 42344
rect 35483 42313 35495 42316
rect 35437 42307 35495 42313
rect 35526 42304 35532 42316
rect 35584 42304 35590 42356
rect 35986 42344 35992 42356
rect 35947 42316 35992 42344
rect 35986 42304 35992 42316
rect 36044 42304 36050 42356
rect 29932 42248 31156 42276
rect 23348 42236 23354 42248
rect 31846 42236 31852 42288
rect 31904 42276 31910 42288
rect 34057 42279 34115 42285
rect 34057 42276 34069 42279
rect 31904 42248 34069 42276
rect 31904 42236 31910 42248
rect 34057 42245 34069 42248
rect 34103 42276 34115 42279
rect 34146 42276 34152 42288
rect 34103 42248 34152 42276
rect 34103 42245 34115 42248
rect 34057 42239 34115 42245
rect 34146 42236 34152 42248
rect 34204 42236 34210 42288
rect 35084 42248 35894 42276
rect 22925 42211 22983 42217
rect 22925 42208 22937 42211
rect 22612 42180 22937 42208
rect 22612 42168 22618 42180
rect 22925 42177 22937 42180
rect 22971 42177 22983 42211
rect 22925 42171 22983 42177
rect 23109 42211 23167 42217
rect 23109 42177 23121 42211
rect 23155 42177 23167 42211
rect 23109 42171 23167 42177
rect 23753 42211 23811 42217
rect 23753 42177 23765 42211
rect 23799 42177 23811 42211
rect 23753 42171 23811 42177
rect 23845 42211 23903 42217
rect 23845 42177 23857 42211
rect 23891 42208 23903 42211
rect 24394 42208 24400 42220
rect 23891 42180 24400 42208
rect 23891 42177 23903 42180
rect 23845 42171 23903 42177
rect 15930 42140 15936 42152
rect 15891 42112 15936 42140
rect 15930 42100 15936 42112
rect 15988 42100 15994 42152
rect 16758 42100 16764 42152
rect 16816 42140 16822 42152
rect 18322 42140 18328 42152
rect 16816 42112 18328 42140
rect 16816 42100 16822 42112
rect 18322 42100 18328 42112
rect 18380 42100 18386 42152
rect 18414 42100 18420 42152
rect 18472 42140 18478 42152
rect 18509 42143 18567 42149
rect 18509 42140 18521 42143
rect 18472 42112 18521 42140
rect 18472 42100 18478 42112
rect 18509 42109 18521 42112
rect 18555 42109 18567 42143
rect 18509 42103 18567 42109
rect 21910 42100 21916 42152
rect 21968 42140 21974 42152
rect 22097 42143 22155 42149
rect 22097 42140 22109 42143
rect 21968 42112 22109 42140
rect 21968 42100 21974 42112
rect 22097 42109 22109 42112
rect 22143 42109 22155 42143
rect 23768 42140 23796 42171
rect 24394 42168 24400 42180
rect 24452 42208 24458 42220
rect 24489 42211 24547 42217
rect 24489 42208 24501 42211
rect 24452 42180 24501 42208
rect 24452 42168 24458 42180
rect 24489 42177 24501 42180
rect 24535 42177 24547 42211
rect 24489 42171 24547 42177
rect 24578 42168 24584 42220
rect 24636 42208 24642 42220
rect 25498 42208 25504 42220
rect 24636 42180 24681 42208
rect 25459 42180 25504 42208
rect 24636 42168 24642 42180
rect 25498 42168 25504 42180
rect 25556 42168 25562 42220
rect 28281 42211 28339 42217
rect 28281 42177 28293 42211
rect 28327 42208 28339 42211
rect 28537 42211 28595 42217
rect 28327 42180 28488 42208
rect 28327 42177 28339 42180
rect 28281 42171 28339 42177
rect 24029 42143 24087 42149
rect 23768 42112 23888 42140
rect 22097 42103 22155 42109
rect 16117 42075 16175 42081
rect 16117 42041 16129 42075
rect 16163 42072 16175 42075
rect 18782 42072 18788 42084
rect 16163 42044 18788 42072
rect 16163 42041 16175 42044
rect 16117 42035 16175 42041
rect 18782 42032 18788 42044
rect 18840 42032 18846 42084
rect 18969 42075 19027 42081
rect 18969 42041 18981 42075
rect 19015 42072 19027 42075
rect 19334 42072 19340 42084
rect 19015 42044 19340 42072
rect 19015 42041 19027 42044
rect 18969 42035 19027 42041
rect 19334 42032 19340 42044
rect 19392 42032 19398 42084
rect 19978 42072 19984 42084
rect 19939 42044 19984 42072
rect 19978 42032 19984 42044
rect 20036 42032 20042 42084
rect 22189 42075 22247 42081
rect 22189 42072 22201 42075
rect 22066 42044 22201 42072
rect 10413 42007 10471 42013
rect 10413 41973 10425 42007
rect 10459 42004 10471 42007
rect 10778 42004 10784 42016
rect 10459 41976 10784 42004
rect 10459 41973 10471 41976
rect 10413 41967 10471 41973
rect 10778 41964 10784 41976
rect 10836 42004 10842 42016
rect 10873 42007 10931 42013
rect 10873 42004 10885 42007
rect 10836 41976 10885 42004
rect 10836 41964 10842 41976
rect 10873 41973 10885 41976
rect 10919 41973 10931 42007
rect 15746 42004 15752 42016
rect 15707 41976 15752 42004
rect 10873 41967 10931 41973
rect 15746 41964 15752 41976
rect 15804 41964 15810 42016
rect 16761 42007 16819 42013
rect 16761 41973 16773 42007
rect 16807 42004 16819 42007
rect 16850 42004 16856 42016
rect 16807 41976 16856 42004
rect 16807 41973 16819 41976
rect 16761 41967 16819 41973
rect 16850 41964 16856 41976
rect 16908 41964 16914 42016
rect 19521 42007 19579 42013
rect 19521 41973 19533 42007
rect 19567 42004 19579 42007
rect 20714 42004 20720 42016
rect 19567 41976 20720 42004
rect 19567 41973 19579 41976
rect 19521 41967 19579 41973
rect 20714 41964 20720 41976
rect 20772 41964 20778 42016
rect 21634 41964 21640 42016
rect 21692 42004 21698 42016
rect 21910 42004 21916 42016
rect 21692 41976 21916 42004
rect 21692 41964 21698 41976
rect 21910 41964 21916 41976
rect 21968 42004 21974 42016
rect 22066 42004 22094 42044
rect 22189 42041 22201 42044
rect 22235 42072 22247 42075
rect 23017 42075 23075 42081
rect 23017 42072 23029 42075
rect 22235 42044 23029 42072
rect 22235 42041 22247 42044
rect 22189 42035 22247 42041
rect 23017 42041 23029 42044
rect 23063 42041 23075 42075
rect 23017 42035 23075 42041
rect 21968 41976 22094 42004
rect 23860 42004 23888 42112
rect 24029 42109 24041 42143
rect 24075 42140 24087 42143
rect 24596 42140 24624 42168
rect 24075 42112 24624 42140
rect 28460 42140 28488 42180
rect 28537 42177 28549 42211
rect 28583 42208 28595 42211
rect 28997 42211 29055 42217
rect 28997 42208 29009 42211
rect 28583 42180 29009 42208
rect 28583 42177 28595 42180
rect 28537 42171 28595 42177
rect 28997 42177 29009 42180
rect 29043 42208 29055 42211
rect 29086 42208 29092 42220
rect 29043 42180 29092 42208
rect 29043 42177 29055 42180
rect 28997 42171 29055 42177
rect 29086 42168 29092 42180
rect 29144 42168 29150 42220
rect 30650 42168 30656 42220
rect 30708 42208 30714 42220
rect 35084 42217 35112 42248
rect 35360 42220 35388 42248
rect 32381 42211 32439 42217
rect 32381 42208 32393 42211
rect 30708 42180 32393 42208
rect 30708 42168 30714 42180
rect 32381 42177 32393 42180
rect 32427 42177 32439 42211
rect 32381 42171 32439 42177
rect 35069 42211 35127 42217
rect 35069 42177 35081 42211
rect 35115 42177 35127 42211
rect 35069 42171 35127 42177
rect 35342 42168 35348 42220
rect 35400 42168 35406 42220
rect 35529 42211 35587 42217
rect 35529 42177 35541 42211
rect 35575 42177 35587 42211
rect 35866 42208 35894 42248
rect 36173 42211 36231 42217
rect 36173 42208 36185 42211
rect 35866 42180 36185 42208
rect 35529 42171 35587 42177
rect 36173 42177 36185 42180
rect 36219 42177 36231 42211
rect 37458 42208 37464 42220
rect 37419 42180 37464 42208
rect 36173 42171 36231 42177
rect 29270 42140 29276 42152
rect 28460 42112 29040 42140
rect 29231 42112 29276 42140
rect 24075 42109 24087 42112
rect 24029 42103 24087 42109
rect 24673 42007 24731 42013
rect 24673 42004 24685 42007
rect 23860 41976 24685 42004
rect 21968 41964 21974 41976
rect 24673 41973 24685 41976
rect 24719 42004 24731 42007
rect 25409 42007 25467 42013
rect 25409 42004 25421 42007
rect 24719 41976 25421 42004
rect 24719 41973 24731 41976
rect 24673 41967 24731 41973
rect 25409 41973 25421 41976
rect 25455 41973 25467 42007
rect 25409 41967 25467 41973
rect 25958 41964 25964 42016
rect 26016 42004 26022 42016
rect 26053 42007 26111 42013
rect 26053 42004 26065 42007
rect 26016 41976 26065 42004
rect 26016 41964 26022 41976
rect 26053 41973 26065 41976
rect 26099 41973 26111 42007
rect 27154 42004 27160 42016
rect 27115 41976 27160 42004
rect 26053 41967 26111 41973
rect 27154 41964 27160 41976
rect 27212 41964 27218 42016
rect 29012 42004 29040 42112
rect 29270 42100 29276 42112
rect 29328 42100 29334 42152
rect 30742 42100 30748 42152
rect 30800 42140 30806 42152
rect 30926 42140 30932 42152
rect 30800 42112 30932 42140
rect 30800 42100 30806 42112
rect 30926 42100 30932 42112
rect 30984 42140 30990 42152
rect 31113 42143 31171 42149
rect 31113 42140 31125 42143
rect 30984 42112 31125 42140
rect 30984 42100 30990 42112
rect 31113 42109 31125 42112
rect 31159 42140 31171 42143
rect 31846 42140 31852 42152
rect 31159 42112 31852 42140
rect 31159 42109 31171 42112
rect 31113 42103 31171 42109
rect 31846 42100 31852 42112
rect 31904 42100 31910 42152
rect 32122 42140 32128 42152
rect 32083 42112 32128 42140
rect 32122 42100 32128 42112
rect 32180 42100 32186 42152
rect 33594 42100 33600 42152
rect 33652 42140 33658 42152
rect 35434 42140 35440 42152
rect 33652 42112 35440 42140
rect 33652 42100 33658 42112
rect 35434 42100 35440 42112
rect 35492 42100 35498 42152
rect 35544 42140 35572 42171
rect 37458 42168 37464 42180
rect 37516 42168 37522 42220
rect 37737 42211 37795 42217
rect 37737 42177 37749 42211
rect 37783 42177 37795 42211
rect 38286 42208 38292 42220
rect 38247 42180 38292 42208
rect 37737 42171 37795 42177
rect 36354 42140 36360 42152
rect 35544 42112 36360 42140
rect 36354 42100 36360 42112
rect 36412 42100 36418 42152
rect 37274 42100 37280 42152
rect 37332 42140 37338 42152
rect 37553 42143 37611 42149
rect 37553 42140 37565 42143
rect 37332 42112 37565 42140
rect 37332 42100 37338 42112
rect 37553 42109 37565 42112
rect 37599 42109 37611 42143
rect 37752 42140 37780 42171
rect 38286 42168 38292 42180
rect 38344 42168 38350 42220
rect 38470 42208 38476 42220
rect 38431 42180 38476 42208
rect 38470 42168 38476 42180
rect 38528 42168 38534 42220
rect 38562 42168 38568 42220
rect 38620 42208 38626 42220
rect 39025 42211 39083 42217
rect 39025 42208 39037 42211
rect 38620 42180 39037 42208
rect 38620 42168 38626 42180
rect 39025 42177 39037 42180
rect 39071 42177 39083 42211
rect 39025 42171 39083 42177
rect 39209 42211 39267 42217
rect 39209 42177 39221 42211
rect 39255 42177 39267 42211
rect 39209 42171 39267 42177
rect 38488 42140 38516 42168
rect 39114 42140 39120 42152
rect 37752 42112 38332 42140
rect 38488 42112 39120 42140
rect 37553 42103 37611 42109
rect 32030 42072 32036 42084
rect 30024 42044 32036 42072
rect 30024 42004 30052 42044
rect 32030 42032 32036 42044
rect 32088 42032 32094 42084
rect 33870 42032 33876 42084
rect 33928 42072 33934 42084
rect 37182 42072 37188 42084
rect 33928 42044 37188 42072
rect 33928 42032 33934 42044
rect 37182 42032 37188 42044
rect 37240 42032 37246 42084
rect 37642 42032 37648 42084
rect 37700 42072 37706 42084
rect 38304 42081 38332 42112
rect 39114 42100 39120 42112
rect 39172 42140 39178 42152
rect 39224 42140 39252 42171
rect 39172 42112 39252 42140
rect 39172 42100 39178 42112
rect 38289 42075 38347 42081
rect 37700 42044 37745 42072
rect 37700 42032 37706 42044
rect 38289 42041 38301 42075
rect 38335 42041 38347 42075
rect 38289 42035 38347 42041
rect 30374 42004 30380 42016
rect 29012 41976 30052 42004
rect 30335 41976 30380 42004
rect 30374 41964 30380 41976
rect 30432 41964 30438 42016
rect 33134 41964 33140 42016
rect 33192 42004 33198 42016
rect 33505 42007 33563 42013
rect 33505 42004 33517 42007
rect 33192 41976 33517 42004
rect 33192 41964 33198 41976
rect 33505 41973 33517 41976
rect 33551 41973 33563 42007
rect 33505 41967 33563 41973
rect 35158 41964 35164 42016
rect 35216 42004 35222 42016
rect 35802 42004 35808 42016
rect 35216 41976 35808 42004
rect 35216 41964 35222 41976
rect 35802 41964 35808 41976
rect 35860 41964 35866 42016
rect 37277 42007 37335 42013
rect 37277 41973 37289 42007
rect 37323 42004 37335 42007
rect 37918 42004 37924 42016
rect 37323 41976 37924 42004
rect 37323 41973 37335 41976
rect 37277 41967 37335 41973
rect 37918 41964 37924 41976
rect 37976 41964 37982 42016
rect 39117 42007 39175 42013
rect 39117 41973 39129 42007
rect 39163 42004 39175 42007
rect 39298 42004 39304 42016
rect 39163 41976 39304 42004
rect 39163 41973 39175 41976
rect 39117 41967 39175 41973
rect 39298 41964 39304 41976
rect 39356 41964 39362 42016
rect 39761 42007 39819 42013
rect 39761 41973 39773 42007
rect 39807 42004 39819 42007
rect 40034 42004 40040 42016
rect 39807 41976 40040 42004
rect 39807 41973 39819 41976
rect 39761 41967 39819 41973
rect 40034 41964 40040 41976
rect 40092 41964 40098 42016
rect 40218 42004 40224 42016
rect 40179 41976 40224 42004
rect 40218 41964 40224 41976
rect 40276 42004 40282 42016
rect 40773 42007 40831 42013
rect 40773 42004 40785 42007
rect 40276 41976 40785 42004
rect 40276 41964 40282 41976
rect 40773 41973 40785 41976
rect 40819 41973 40831 42007
rect 40773 41967 40831 41973
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 12437 41803 12495 41809
rect 12437 41769 12449 41803
rect 12483 41800 12495 41803
rect 13538 41800 13544 41812
rect 12483 41772 13544 41800
rect 12483 41769 12495 41772
rect 12437 41763 12495 41769
rect 13538 41760 13544 41772
rect 13596 41760 13602 41812
rect 14182 41800 14188 41812
rect 14143 41772 14188 41800
rect 14182 41760 14188 41772
rect 14240 41760 14246 41812
rect 15562 41800 15568 41812
rect 15475 41772 15568 41800
rect 15562 41760 15568 41772
rect 15620 41800 15626 41812
rect 15746 41800 15752 41812
rect 15620 41772 15752 41800
rect 15620 41760 15626 41772
rect 15746 41760 15752 41772
rect 15804 41760 15810 41812
rect 17405 41803 17463 41809
rect 16592 41772 17080 41800
rect 15013 41735 15071 41741
rect 15013 41701 15025 41735
rect 15059 41732 15071 41735
rect 16592 41732 16620 41772
rect 15059 41704 16620 41732
rect 15059 41701 15071 41704
rect 15013 41695 15071 41701
rect 17052 41664 17080 41772
rect 17405 41769 17417 41803
rect 17451 41800 17463 41803
rect 17678 41800 17684 41812
rect 17451 41772 17684 41800
rect 17451 41769 17463 41772
rect 17405 41763 17463 41769
rect 17678 41760 17684 41772
rect 17736 41760 17742 41812
rect 18414 41800 18420 41812
rect 18375 41772 18420 41800
rect 18414 41760 18420 41772
rect 18472 41760 18478 41812
rect 19426 41760 19432 41812
rect 19484 41800 19490 41812
rect 19797 41803 19855 41809
rect 19797 41800 19809 41803
rect 19484 41772 19809 41800
rect 19484 41760 19490 41772
rect 19797 41769 19809 41772
rect 19843 41769 19855 41803
rect 20714 41800 20720 41812
rect 20675 41772 20720 41800
rect 19797 41763 19855 41769
rect 20714 41760 20720 41772
rect 20772 41760 20778 41812
rect 22005 41803 22063 41809
rect 22005 41769 22017 41803
rect 22051 41800 22063 41803
rect 22278 41800 22284 41812
rect 22051 41772 22284 41800
rect 22051 41769 22063 41772
rect 22005 41763 22063 41769
rect 22278 41760 22284 41772
rect 22336 41760 22342 41812
rect 23845 41803 23903 41809
rect 23845 41769 23857 41803
rect 23891 41800 23903 41803
rect 25958 41800 25964 41812
rect 23891 41772 25964 41800
rect 23891 41769 23903 41772
rect 23845 41763 23903 41769
rect 25958 41760 25964 41772
rect 26016 41760 26022 41812
rect 26513 41803 26571 41809
rect 26513 41769 26525 41803
rect 26559 41800 26571 41803
rect 27062 41800 27068 41812
rect 26559 41772 27068 41800
rect 26559 41769 26571 41772
rect 26513 41763 26571 41769
rect 27062 41760 27068 41772
rect 27120 41760 27126 41812
rect 27706 41760 27712 41812
rect 27764 41800 27770 41812
rect 28074 41800 28080 41812
rect 27764 41772 28080 41800
rect 27764 41760 27770 41772
rect 28074 41760 28080 41772
rect 28132 41800 28138 41812
rect 28261 41803 28319 41809
rect 28261 41800 28273 41803
rect 28132 41772 28273 41800
rect 28132 41760 28138 41772
rect 28261 41769 28273 41772
rect 28307 41769 28319 41803
rect 32585 41803 32643 41809
rect 28261 41763 28319 41769
rect 28368 41772 31754 41800
rect 20732 41732 20760 41760
rect 22741 41735 22799 41741
rect 20732 41704 22048 41732
rect 18782 41664 18788 41676
rect 17052 41636 17172 41664
rect 14734 41556 14740 41608
rect 14792 41596 14798 41608
rect 15013 41599 15071 41605
rect 14792 41568 14964 41596
rect 14792 41556 14798 41568
rect 11054 41488 11060 41540
rect 11112 41528 11118 41540
rect 11793 41531 11851 41537
rect 11793 41528 11805 41531
rect 11112 41500 11805 41528
rect 11112 41488 11118 41500
rect 11793 41497 11805 41500
rect 11839 41528 11851 41531
rect 12158 41528 12164 41540
rect 11839 41500 12164 41528
rect 11839 41497 11851 41500
rect 11793 41491 11851 41497
rect 12158 41488 12164 41500
rect 12216 41488 12222 41540
rect 14936 41528 14964 41568
rect 15013 41565 15025 41599
rect 15059 41596 15071 41599
rect 15473 41599 15531 41605
rect 15473 41596 15485 41599
rect 15059 41568 15485 41596
rect 15059 41565 15071 41568
rect 15013 41559 15071 41565
rect 15473 41565 15485 41568
rect 15519 41596 15531 41599
rect 15654 41596 15660 41608
rect 15519 41568 15660 41596
rect 15519 41565 15531 41568
rect 15473 41559 15531 41565
rect 15654 41556 15660 41568
rect 15712 41556 15718 41608
rect 15749 41599 15807 41605
rect 15749 41565 15761 41599
rect 15795 41596 15807 41599
rect 15930 41596 15936 41608
rect 15795 41568 15936 41596
rect 15795 41565 15807 41568
rect 15749 41559 15807 41565
rect 15764 41528 15792 41559
rect 15930 41556 15936 41568
rect 15988 41556 15994 41608
rect 16758 41596 16764 41608
rect 16719 41568 16764 41596
rect 16758 41556 16764 41568
rect 16816 41556 16822 41608
rect 16942 41596 16948 41608
rect 16903 41568 16948 41596
rect 16942 41556 16948 41568
rect 17000 41556 17006 41608
rect 17144 41605 17172 41636
rect 18340 41636 18788 41664
rect 18340 41605 18368 41636
rect 18782 41624 18788 41636
rect 18840 41624 18846 41676
rect 19150 41624 19156 41676
rect 19208 41664 19214 41676
rect 19337 41667 19395 41673
rect 19337 41664 19349 41667
rect 19208 41636 19349 41664
rect 19208 41624 19214 41636
rect 19337 41633 19349 41636
rect 19383 41664 19395 41667
rect 20530 41664 20536 41676
rect 19383 41636 20536 41664
rect 19383 41633 19395 41636
rect 19337 41627 19395 41633
rect 20530 41624 20536 41636
rect 20588 41664 20594 41676
rect 21358 41664 21364 41676
rect 20588 41636 21364 41664
rect 20588 41624 20594 41636
rect 21358 41624 21364 41636
rect 21416 41624 21422 41676
rect 17037 41599 17095 41605
rect 17037 41565 17049 41599
rect 17083 41565 17095 41599
rect 17037 41559 17095 41565
rect 17129 41599 17187 41605
rect 17129 41565 17141 41599
rect 17175 41565 17187 41599
rect 17129 41559 17187 41565
rect 18325 41599 18383 41605
rect 18325 41565 18337 41599
rect 18371 41565 18383 41599
rect 18506 41596 18512 41608
rect 18467 41568 18512 41596
rect 18325 41559 18383 41565
rect 14936 41500 15792 41528
rect 16114 41488 16120 41540
rect 16172 41528 16178 41540
rect 17052 41528 17080 41559
rect 18506 41556 18512 41568
rect 18564 41556 18570 41608
rect 19426 41596 19432 41608
rect 19387 41568 19432 41596
rect 19426 41556 19432 41568
rect 19484 41556 19490 41608
rect 19613 41599 19671 41605
rect 19613 41565 19625 41599
rect 19659 41596 19671 41599
rect 20346 41596 20352 41608
rect 19659 41568 20352 41596
rect 19659 41565 19671 41568
rect 19613 41559 19671 41565
rect 20346 41556 20352 41568
rect 20404 41556 20410 41608
rect 21726 41556 21732 41608
rect 21784 41596 21790 41608
rect 21821 41599 21879 41605
rect 21821 41596 21833 41599
rect 21784 41568 21833 41596
rect 21784 41556 21790 41568
rect 21821 41565 21833 41568
rect 21867 41565 21879 41599
rect 21821 41559 21879 41565
rect 16172 41500 17080 41528
rect 16172 41488 16178 41500
rect 17218 41488 17224 41540
rect 17276 41528 17282 41540
rect 18414 41528 18420 41540
rect 17276 41500 18420 41528
rect 17276 41488 17282 41500
rect 18414 41488 18420 41500
rect 18472 41488 18478 41540
rect 21913 41531 21971 41537
rect 21913 41528 21925 41531
rect 21284 41500 21925 41528
rect 9582 41420 9588 41472
rect 9640 41460 9646 41472
rect 11241 41463 11299 41469
rect 11241 41460 11253 41463
rect 9640 41432 11253 41460
rect 9640 41420 9646 41432
rect 11241 41429 11253 41432
rect 11287 41429 11299 41463
rect 11241 41423 11299 41429
rect 12989 41463 13047 41469
rect 12989 41429 13001 41463
rect 13035 41460 13047 41463
rect 13449 41463 13507 41469
rect 13449 41460 13461 41463
rect 13035 41432 13461 41460
rect 13035 41429 13047 41432
rect 12989 41423 13047 41429
rect 13449 41429 13461 41432
rect 13495 41460 13507 41463
rect 13538 41460 13544 41472
rect 13495 41432 13544 41460
rect 13495 41429 13507 41432
rect 13449 41423 13507 41429
rect 13538 41420 13544 41432
rect 13596 41420 13602 41472
rect 14829 41463 14887 41469
rect 14829 41429 14841 41463
rect 14875 41460 14887 41463
rect 15102 41460 15108 41472
rect 14875 41432 15108 41460
rect 14875 41429 14887 41432
rect 14829 41423 14887 41429
rect 15102 41420 15108 41432
rect 15160 41420 15166 41472
rect 15933 41463 15991 41469
rect 15933 41429 15945 41463
rect 15979 41460 15991 41463
rect 16758 41460 16764 41472
rect 15979 41432 16764 41460
rect 15979 41429 15991 41432
rect 15933 41423 15991 41429
rect 16758 41420 16764 41432
rect 16816 41420 16822 41472
rect 17954 41420 17960 41472
rect 18012 41460 18018 41472
rect 21082 41460 21088 41472
rect 18012 41432 21088 41460
rect 18012 41420 18018 41432
rect 21082 41420 21088 41432
rect 21140 41460 21146 41472
rect 21284 41469 21312 41500
rect 21913 41497 21925 41500
rect 21959 41497 21971 41531
rect 21913 41491 21971 41497
rect 21269 41463 21327 41469
rect 21269 41460 21281 41463
rect 21140 41432 21281 41460
rect 21140 41420 21146 41432
rect 21269 41429 21281 41432
rect 21315 41429 21327 41463
rect 22020 41460 22048 41704
rect 22741 41701 22753 41735
rect 22787 41732 22799 41735
rect 23106 41732 23112 41744
rect 22787 41704 23112 41732
rect 22787 41701 22799 41704
rect 22741 41695 22799 41701
rect 23106 41692 23112 41704
rect 23164 41732 23170 41744
rect 23164 41704 24900 41732
rect 23164 41692 23170 41704
rect 24486 41664 24492 41676
rect 24447 41636 24492 41664
rect 24486 41624 24492 41636
rect 24544 41624 24550 41676
rect 24872 41664 24900 41704
rect 25406 41692 25412 41744
rect 25464 41732 25470 41744
rect 25501 41735 25559 41741
rect 25501 41732 25513 41735
rect 25464 41704 25513 41732
rect 25464 41692 25470 41704
rect 25501 41701 25513 41704
rect 25547 41732 25559 41735
rect 27338 41732 27344 41744
rect 25547 41704 27344 41732
rect 25547 41701 25559 41704
rect 25501 41695 25559 41701
rect 27338 41692 27344 41704
rect 27396 41692 27402 41744
rect 28368 41664 28396 41772
rect 31726 41732 31754 41772
rect 32585 41769 32597 41803
rect 32631 41800 32643 41803
rect 34238 41800 34244 41812
rect 32631 41772 34244 41800
rect 32631 41769 32643 41772
rect 32585 41763 32643 41769
rect 34238 41760 34244 41772
rect 34296 41760 34302 41812
rect 35342 41760 35348 41812
rect 35400 41800 35406 41812
rect 35437 41803 35495 41809
rect 35437 41800 35449 41803
rect 35400 41772 35449 41800
rect 35400 41760 35406 41772
rect 35437 41769 35449 41772
rect 35483 41769 35495 41803
rect 36354 41800 36360 41812
rect 36315 41772 36360 41800
rect 35437 41763 35495 41769
rect 36354 41760 36360 41772
rect 36412 41760 36418 41812
rect 38286 41800 38292 41812
rect 38247 41772 38292 41800
rect 38286 41760 38292 41772
rect 38344 41760 38350 41812
rect 38473 41803 38531 41809
rect 38473 41769 38485 41803
rect 38519 41800 38531 41803
rect 40034 41800 40040 41812
rect 38519 41772 40040 41800
rect 38519 41769 38531 41772
rect 38473 41763 38531 41769
rect 34514 41732 34520 41744
rect 31726 41704 34520 41732
rect 34514 41692 34520 41704
rect 34572 41692 34578 41744
rect 34793 41735 34851 41741
rect 34793 41701 34805 41735
rect 34839 41732 34851 41735
rect 34882 41732 34888 41744
rect 34839 41704 34888 41732
rect 34839 41701 34851 41704
rect 34793 41695 34851 41701
rect 34882 41692 34888 41704
rect 34940 41732 34946 41744
rect 36170 41732 36176 41744
rect 34940 41704 36176 41732
rect 34940 41692 34946 41704
rect 36170 41692 36176 41704
rect 36228 41692 36234 41744
rect 38488 41732 38516 41763
rect 40034 41760 40040 41772
rect 40092 41760 40098 41812
rect 37476 41704 38516 41732
rect 24872 41636 28396 41664
rect 29086 41624 29092 41676
rect 29144 41664 29150 41676
rect 29549 41667 29607 41673
rect 29549 41664 29561 41667
rect 29144 41636 29561 41664
rect 29144 41624 29150 41636
rect 29549 41633 29561 41636
rect 29595 41633 29607 41667
rect 31202 41664 31208 41676
rect 31163 41636 31208 41664
rect 29549 41627 29607 41633
rect 31202 41624 31208 41636
rect 31260 41624 31266 41676
rect 33686 41664 33692 41676
rect 31312 41636 33692 41664
rect 22097 41599 22155 41605
rect 22097 41565 22109 41599
rect 22143 41596 22155 41599
rect 22554 41596 22560 41608
rect 22143 41568 22560 41596
rect 22143 41565 22155 41568
rect 22097 41559 22155 41565
rect 22554 41556 22560 41568
rect 22612 41556 22618 41608
rect 23934 41556 23940 41608
rect 23992 41596 23998 41608
rect 24397 41599 24455 41605
rect 24397 41596 24409 41599
rect 23992 41568 24409 41596
rect 23992 41556 23998 41568
rect 24397 41565 24409 41568
rect 24443 41565 24455 41599
rect 24397 41559 24455 41565
rect 24581 41599 24639 41605
rect 24581 41565 24593 41599
rect 24627 41596 24639 41599
rect 24670 41596 24676 41608
rect 24627 41568 24676 41596
rect 24627 41565 24639 41568
rect 24581 41559 24639 41565
rect 24670 41556 24676 41568
rect 24728 41556 24734 41608
rect 27801 41599 27859 41605
rect 27801 41565 27813 41599
rect 27847 41596 27859 41599
rect 28994 41596 29000 41608
rect 27847 41568 29000 41596
rect 27847 41565 27859 41568
rect 27801 41559 27859 41565
rect 28994 41556 29000 41568
rect 29052 41556 29058 41608
rect 29825 41599 29883 41605
rect 29825 41565 29837 41599
rect 29871 41596 29883 41599
rect 29914 41596 29920 41608
rect 29871 41568 29920 41596
rect 29871 41565 29883 41568
rect 29825 41559 29883 41565
rect 29914 41556 29920 41568
rect 29972 41556 29978 41608
rect 30190 41556 30196 41608
rect 30248 41596 30254 41608
rect 31312 41596 31340 41636
rect 33686 41624 33692 41636
rect 33744 41624 33750 41676
rect 33965 41667 34023 41673
rect 33965 41633 33977 41667
rect 34011 41664 34023 41667
rect 36538 41664 36544 41676
rect 34011 41636 36544 41664
rect 34011 41633 34023 41636
rect 33965 41627 34023 41633
rect 36538 41624 36544 41636
rect 36596 41624 36602 41676
rect 32398 41596 32404 41608
rect 30248 41568 31340 41596
rect 32359 41568 32404 41596
rect 30248 41556 30254 41568
rect 32398 41556 32404 41568
rect 32456 41556 32462 41608
rect 32585 41599 32643 41605
rect 32585 41565 32597 41599
rect 32631 41596 32643 41599
rect 33410 41596 33416 41608
rect 32631 41568 33416 41596
rect 32631 41565 32643 41568
rect 32585 41559 32643 41565
rect 33410 41556 33416 41568
rect 33468 41556 33474 41608
rect 33594 41596 33600 41608
rect 33555 41568 33600 41596
rect 33594 41556 33600 41568
rect 33652 41556 33658 41608
rect 33870 41556 33876 41608
rect 33928 41596 33934 41608
rect 34057 41599 34115 41605
rect 34057 41596 34069 41599
rect 33928 41568 34069 41596
rect 33928 41556 33934 41568
rect 34057 41565 34069 41568
rect 34103 41565 34115 41599
rect 34057 41559 34115 41565
rect 35710 41556 35716 41608
rect 35768 41596 35774 41608
rect 35805 41599 35863 41605
rect 35805 41596 35817 41599
rect 35768 41568 35817 41596
rect 35768 41556 35774 41568
rect 35805 41565 35817 41568
rect 35851 41596 35863 41599
rect 36265 41599 36323 41605
rect 36265 41596 36277 41599
rect 35851 41568 36277 41596
rect 35851 41565 35863 41568
rect 35805 41559 35863 41565
rect 36265 41565 36277 41568
rect 36311 41565 36323 41599
rect 36265 41559 36323 41565
rect 36449 41599 36507 41605
rect 36449 41565 36461 41599
rect 36495 41596 36507 41599
rect 37476 41596 37504 41704
rect 38562 41692 38568 41744
rect 38620 41732 38626 41744
rect 39853 41735 39911 41741
rect 39853 41732 39865 41735
rect 38620 41704 39865 41732
rect 38620 41692 38626 41704
rect 39853 41701 39865 41704
rect 39899 41732 39911 41735
rect 40218 41732 40224 41744
rect 39899 41704 40224 41732
rect 39899 41701 39911 41704
rect 39853 41695 39911 41701
rect 40218 41692 40224 41704
rect 40276 41692 40282 41744
rect 37734 41664 37740 41676
rect 37695 41636 37740 41664
rect 37734 41624 37740 41636
rect 37792 41624 37798 41676
rect 39209 41667 39267 41673
rect 39209 41664 39221 41667
rect 38212 41636 39221 41664
rect 37642 41596 37648 41608
rect 36495 41568 37504 41596
rect 37555 41568 37648 41596
rect 36495 41565 36507 41568
rect 36449 41559 36507 41565
rect 33689 41531 33747 41537
rect 25332 41500 29040 41528
rect 25332 41472 25360 41500
rect 23106 41460 23112 41472
rect 22020 41432 23112 41460
rect 21269 41423 21327 41429
rect 23106 41420 23112 41432
rect 23164 41420 23170 41472
rect 23293 41463 23351 41469
rect 23293 41429 23305 41463
rect 23339 41460 23351 41463
rect 23474 41460 23480 41472
rect 23339 41432 23480 41460
rect 23339 41429 23351 41432
rect 23293 41423 23351 41429
rect 23474 41420 23480 41432
rect 23532 41460 23538 41472
rect 24210 41460 24216 41472
rect 23532 41432 24216 41460
rect 23532 41420 23538 41432
rect 24210 41420 24216 41432
rect 24268 41420 24274 41472
rect 25314 41420 25320 41472
rect 25372 41420 25378 41472
rect 25774 41420 25780 41472
rect 25832 41460 25838 41472
rect 27706 41460 27712 41472
rect 25832 41432 27712 41460
rect 25832 41420 25838 41432
rect 27706 41420 27712 41432
rect 27764 41420 27770 41472
rect 28902 41460 28908 41472
rect 28863 41432 28908 41460
rect 28902 41420 28908 41432
rect 28960 41420 28966 41472
rect 29012 41460 29040 41500
rect 33689 41497 33701 41531
rect 33735 41528 33747 41531
rect 33735 41500 34284 41528
rect 33735 41497 33747 41500
rect 33689 41491 33747 41497
rect 30466 41460 30472 41472
rect 29012 41432 30472 41460
rect 30466 41420 30472 41432
rect 30524 41420 30530 41472
rect 31757 41463 31815 41469
rect 31757 41429 31769 41463
rect 31803 41460 31815 41463
rect 32490 41460 32496 41472
rect 31803 41432 32496 41460
rect 31803 41429 31815 41432
rect 31757 41423 31815 41429
rect 32490 41420 32496 41432
rect 32548 41420 32554 41472
rect 33318 41460 33324 41472
rect 33279 41432 33324 41460
rect 33318 41420 33324 41432
rect 33376 41420 33382 41472
rect 33778 41420 33784 41472
rect 33836 41460 33842 41472
rect 34256 41460 34284 41500
rect 34330 41488 34336 41540
rect 34388 41528 34394 41540
rect 35621 41531 35679 41537
rect 35621 41528 35633 41531
rect 34388 41500 35633 41528
rect 34388 41488 34394 41500
rect 35621 41497 35633 41500
rect 35667 41497 35679 41531
rect 35621 41491 35679 41497
rect 34606 41460 34612 41472
rect 33836 41432 33881 41460
rect 34256 41432 34612 41460
rect 33836 41420 33842 41432
rect 34606 41420 34612 41432
rect 34664 41420 34670 41472
rect 35636 41460 35664 41491
rect 36464 41460 36492 41559
rect 37642 41556 37648 41568
rect 37700 41596 37706 41608
rect 38212 41596 38240 41636
rect 39209 41633 39221 41636
rect 39255 41633 39267 41667
rect 39209 41627 39267 41633
rect 38746 41596 38752 41608
rect 37700 41568 38240 41596
rect 38580 41568 38752 41596
rect 37700 41556 37706 41568
rect 38457 41531 38515 41537
rect 38457 41497 38469 41531
rect 38503 41528 38515 41531
rect 38580 41528 38608 41568
rect 38746 41556 38752 41568
rect 38804 41596 38810 41608
rect 39117 41599 39175 41605
rect 39117 41596 39129 41599
rect 38804 41568 39129 41596
rect 38804 41556 38810 41568
rect 39117 41565 39129 41568
rect 39163 41565 39175 41599
rect 39298 41596 39304 41608
rect 39259 41568 39304 41596
rect 39117 41559 39175 41565
rect 39298 41556 39304 41568
rect 39356 41556 39362 41608
rect 38503 41500 38608 41528
rect 38657 41531 38715 41537
rect 38503 41497 38515 41500
rect 38457 41491 38515 41497
rect 38657 41497 38669 41531
rect 38703 41528 38715 41531
rect 40957 41531 41015 41537
rect 40957 41528 40969 41531
rect 38703 41500 40969 41528
rect 38703 41497 38715 41500
rect 38657 41491 38715 41497
rect 40957 41497 40969 41500
rect 41003 41497 41015 41531
rect 40957 41491 41015 41497
rect 35636 41432 36492 41460
rect 36998 41420 37004 41472
rect 37056 41460 37062 41472
rect 37277 41463 37335 41469
rect 37277 41460 37289 41463
rect 37056 41432 37289 41460
rect 37056 41420 37062 41432
rect 37277 41429 37289 41432
rect 37323 41429 37335 41463
rect 37277 41423 37335 41429
rect 38010 41420 38016 41472
rect 38068 41460 38074 41472
rect 38286 41460 38292 41472
rect 38068 41432 38292 41460
rect 38068 41420 38074 41432
rect 38286 41420 38292 41432
rect 38344 41460 38350 41472
rect 38672 41460 38700 41491
rect 40494 41460 40500 41472
rect 38344 41432 38700 41460
rect 40455 41432 40500 41460
rect 38344 41420 38350 41432
rect 40494 41420 40500 41432
rect 40552 41420 40558 41472
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 12529 41259 12587 41265
rect 12529 41225 12541 41259
rect 12575 41256 12587 41259
rect 13538 41256 13544 41268
rect 12575 41228 13544 41256
rect 12575 41225 12587 41228
rect 12529 41219 12587 41225
rect 13538 41216 13544 41228
rect 13596 41216 13602 41268
rect 13633 41259 13691 41265
rect 13633 41225 13645 41259
rect 13679 41256 13691 41259
rect 13814 41256 13820 41268
rect 13679 41228 13820 41256
rect 13679 41225 13691 41228
rect 13633 41219 13691 41225
rect 13814 41216 13820 41228
rect 13872 41216 13878 41268
rect 14185 41259 14243 41265
rect 14185 41225 14197 41259
rect 14231 41256 14243 41259
rect 14734 41256 14740 41268
rect 14231 41228 14740 41256
rect 14231 41225 14243 41228
rect 14185 41219 14243 41225
rect 14734 41216 14740 41228
rect 14792 41216 14798 41268
rect 15102 41256 15108 41268
rect 15063 41228 15108 41256
rect 15102 41216 15108 41228
rect 15160 41256 15166 41268
rect 16114 41256 16120 41268
rect 15160 41228 15884 41256
rect 16075 41228 16120 41256
rect 15160 41216 15166 41228
rect 14921 41191 14979 41197
rect 14921 41188 14933 41191
rect 14108 41160 14933 41188
rect 11054 41080 11060 41132
rect 11112 41120 11118 41132
rect 14108 41129 14136 41160
rect 14921 41157 14933 41160
rect 14967 41157 14979 41191
rect 14921 41151 14979 41157
rect 15654 41148 15660 41200
rect 15712 41148 15718 41200
rect 14093 41123 14151 41129
rect 14093 41120 14105 41123
rect 11112 41092 14105 41120
rect 11112 41080 11118 41092
rect 14093 41089 14105 41092
rect 14139 41089 14151 41123
rect 14093 41083 14151 41089
rect 14277 41123 14335 41129
rect 14277 41089 14289 41123
rect 14323 41120 14335 41123
rect 14737 41123 14795 41129
rect 14737 41120 14749 41123
rect 14323 41092 14749 41120
rect 14323 41089 14335 41092
rect 14277 41083 14335 41089
rect 14737 41089 14749 41092
rect 14783 41120 14795 41123
rect 15194 41120 15200 41132
rect 14783 41092 15200 41120
rect 14783 41089 14795 41092
rect 14737 41083 14795 41089
rect 15194 41080 15200 41092
rect 15252 41080 15258 41132
rect 15672 41120 15700 41148
rect 15856 41129 15884 41228
rect 16114 41216 16120 41228
rect 16172 41216 16178 41268
rect 16942 41216 16948 41268
rect 17000 41256 17006 41268
rect 17681 41259 17739 41265
rect 17681 41256 17693 41259
rect 17000 41228 17693 41256
rect 17000 41216 17006 41228
rect 17681 41225 17693 41228
rect 17727 41225 17739 41259
rect 17681 41219 17739 41225
rect 18138 41216 18144 41268
rect 18196 41256 18202 41268
rect 19702 41256 19708 41268
rect 18196 41228 19288 41256
rect 18196 41216 18202 41228
rect 17586 41148 17592 41200
rect 17644 41188 17650 41200
rect 18693 41191 18751 41197
rect 17644 41160 18552 41188
rect 17644 41148 17650 41160
rect 15749 41123 15807 41129
rect 15749 41120 15761 41123
rect 15672 41092 15761 41120
rect 15749 41089 15761 41092
rect 15795 41089 15807 41123
rect 15749 41083 15807 41089
rect 15841 41123 15899 41129
rect 15841 41089 15853 41123
rect 15887 41089 15899 41123
rect 15841 41083 15899 41089
rect 15930 41080 15936 41132
rect 15988 41120 15994 41132
rect 16850 41120 16856 41132
rect 15988 41092 16033 41120
rect 16811 41092 16856 41120
rect 15988 41080 15994 41092
rect 16850 41080 16856 41092
rect 16908 41080 16914 41132
rect 17696 41129 17724 41160
rect 17681 41123 17739 41129
rect 17681 41089 17693 41123
rect 17727 41089 17739 41123
rect 17681 41083 17739 41089
rect 17865 41123 17923 41129
rect 17865 41089 17877 41123
rect 17911 41120 17923 41123
rect 18138 41120 18144 41132
rect 17911 41092 18144 41120
rect 17911 41089 17923 41092
rect 17865 41083 17923 41089
rect 11977 41055 12035 41061
rect 11977 41021 11989 41055
rect 12023 41052 12035 41055
rect 15654 41052 15660 41064
rect 12023 41024 15660 41052
rect 12023 41021 12035 41024
rect 11977 41015 12035 41021
rect 15654 41012 15660 41024
rect 15712 41012 15718 41064
rect 16758 41052 16764 41064
rect 16719 41024 16764 41052
rect 16758 41012 16764 41024
rect 16816 41012 16822 41064
rect 17880 41052 17908 41083
rect 18138 41080 18144 41092
rect 18196 41080 18202 41132
rect 18414 41120 18420 41132
rect 18375 41092 18420 41120
rect 18414 41080 18420 41092
rect 18472 41080 18478 41132
rect 18524 41129 18552 41160
rect 18693 41157 18705 41191
rect 18739 41188 18751 41191
rect 18874 41188 18880 41200
rect 18739 41160 18880 41188
rect 18739 41157 18751 41160
rect 18693 41151 18751 41157
rect 18874 41148 18880 41160
rect 18932 41148 18938 41200
rect 19260 41132 19288 41228
rect 19444 41228 19708 41256
rect 19444 41197 19472 41228
rect 19702 41216 19708 41228
rect 19760 41216 19766 41268
rect 19797 41259 19855 41265
rect 19797 41225 19809 41259
rect 19843 41256 19855 41259
rect 20070 41256 20076 41268
rect 19843 41228 20076 41256
rect 19843 41225 19855 41228
rect 19797 41219 19855 41225
rect 20070 41216 20076 41228
rect 20128 41216 20134 41268
rect 20346 41256 20352 41268
rect 20307 41228 20352 41256
rect 20346 41216 20352 41228
rect 20404 41216 20410 41268
rect 22002 41216 22008 41268
rect 22060 41256 22066 41268
rect 22741 41259 22799 41265
rect 22741 41256 22753 41259
rect 22060 41228 22753 41256
rect 22060 41216 22066 41228
rect 22741 41225 22753 41228
rect 22787 41256 22799 41259
rect 23014 41256 23020 41268
rect 22787 41228 23020 41256
rect 22787 41225 22799 41228
rect 22741 41219 22799 41225
rect 23014 41216 23020 41228
rect 23072 41216 23078 41268
rect 23385 41259 23443 41265
rect 23385 41225 23397 41259
rect 23431 41256 23443 41259
rect 23937 41259 23995 41265
rect 23937 41256 23949 41259
rect 23431 41228 23949 41256
rect 23431 41225 23443 41228
rect 23385 41219 23443 41225
rect 23937 41225 23949 41228
rect 23983 41256 23995 41259
rect 24302 41256 24308 41268
rect 23983 41228 24308 41256
rect 23983 41225 23995 41228
rect 23937 41219 23995 41225
rect 24302 41216 24308 41228
rect 24360 41256 24366 41268
rect 26237 41259 26295 41265
rect 26237 41256 26249 41259
rect 24360 41228 26249 41256
rect 24360 41216 24366 41228
rect 26237 41225 26249 41228
rect 26283 41256 26295 41259
rect 27430 41256 27436 41268
rect 26283 41228 27436 41256
rect 26283 41225 26295 41228
rect 26237 41219 26295 41225
rect 27430 41216 27436 41228
rect 27488 41216 27494 41268
rect 27798 41256 27804 41268
rect 27759 41228 27804 41256
rect 27798 41216 27804 41228
rect 27856 41216 27862 41268
rect 29086 41256 29092 41268
rect 29047 41228 29092 41256
rect 29086 41216 29092 41228
rect 29144 41216 29150 41268
rect 33778 41216 33784 41268
rect 33836 41256 33842 41268
rect 34333 41259 34391 41265
rect 34333 41256 34345 41259
rect 33836 41228 34345 41256
rect 33836 41216 33842 41228
rect 34333 41225 34345 41228
rect 34379 41225 34391 41259
rect 36538 41256 36544 41268
rect 36499 41228 36544 41256
rect 34333 41219 34391 41225
rect 36538 41216 36544 41228
rect 36596 41216 36602 41268
rect 38657 41259 38715 41265
rect 38657 41225 38669 41259
rect 38703 41256 38715 41259
rect 38746 41256 38752 41268
rect 38703 41228 38752 41256
rect 38703 41225 38715 41228
rect 38657 41219 38715 41225
rect 38746 41216 38752 41228
rect 38804 41216 38810 41268
rect 40218 41216 40224 41268
rect 40276 41256 40282 41268
rect 40773 41259 40831 41265
rect 40773 41256 40785 41259
rect 40276 41228 40785 41256
rect 40276 41216 40282 41228
rect 40773 41225 40785 41228
rect 40819 41225 40831 41259
rect 40773 41219 40831 41225
rect 19429 41191 19487 41197
rect 19429 41157 19441 41191
rect 19475 41157 19487 41191
rect 19978 41188 19984 41200
rect 19429 41151 19487 41157
rect 19536 41160 19984 41188
rect 18509 41123 18567 41129
rect 18509 41089 18521 41123
rect 18555 41120 18567 41123
rect 19058 41120 19064 41132
rect 18555 41092 19064 41120
rect 18555 41089 18567 41092
rect 18509 41083 18567 41089
rect 19058 41080 19064 41092
rect 19116 41080 19122 41132
rect 19153 41123 19211 41129
rect 19153 41089 19165 41123
rect 19199 41089 19211 41123
rect 19153 41083 19211 41089
rect 17144 41024 17908 41052
rect 10965 40919 11023 40925
rect 10965 40885 10977 40919
rect 11011 40916 11023 40919
rect 11054 40916 11060 40928
rect 11011 40888 11060 40916
rect 11011 40885 11023 40888
rect 10965 40879 11023 40885
rect 11054 40876 11060 40888
rect 11112 40876 11118 40928
rect 12710 40876 12716 40928
rect 12768 40916 12774 40928
rect 12989 40919 13047 40925
rect 12989 40916 13001 40919
rect 12768 40888 13001 40916
rect 12768 40876 12774 40888
rect 12989 40885 13001 40888
rect 13035 40885 13047 40919
rect 12989 40879 13047 40885
rect 13538 40876 13544 40928
rect 13596 40916 13602 40928
rect 17144 40916 17172 41024
rect 18322 41012 18328 41064
rect 18380 41052 18386 41064
rect 19168 41052 19196 41083
rect 19242 41080 19248 41132
rect 19300 41120 19306 41132
rect 19536 41129 19564 41160
rect 19978 41148 19984 41160
rect 20036 41148 20042 41200
rect 21269 41191 21327 41197
rect 21269 41188 21281 41191
rect 20180 41160 21281 41188
rect 19521 41123 19579 41129
rect 19521 41120 19533 41123
rect 19300 41092 19393 41120
rect 19444 41092 19533 41120
rect 19300 41080 19306 41092
rect 19444 41064 19472 41092
rect 19521 41089 19533 41092
rect 19567 41089 19579 41123
rect 19521 41083 19579 41089
rect 19610 41080 19616 41132
rect 19668 41129 19674 41132
rect 19668 41123 19695 41129
rect 19683 41089 19695 41123
rect 19668 41083 19695 41089
rect 19668 41080 19674 41083
rect 18380 41024 19288 41052
rect 18380 41012 18386 41024
rect 17221 40987 17279 40993
rect 17221 40953 17233 40987
rect 17267 40984 17279 40987
rect 18506 40984 18512 40996
rect 17267 40956 18512 40984
rect 17267 40953 17279 40956
rect 17221 40947 17279 40953
rect 18506 40944 18512 40956
rect 18564 40944 18570 40996
rect 19260 40984 19288 41024
rect 19426 41012 19432 41064
rect 19484 41012 19490 41064
rect 20180 41052 20208 41160
rect 21269 41157 21281 41160
rect 21315 41188 21327 41191
rect 23474 41188 23480 41200
rect 21315 41160 23480 41188
rect 21315 41157 21327 41160
rect 21269 41151 21327 41157
rect 23474 41148 23480 41160
rect 23532 41148 23538 41200
rect 25958 41148 25964 41200
rect 26016 41188 26022 41200
rect 26973 41191 27031 41197
rect 26973 41188 26985 41191
rect 26016 41160 26985 41188
rect 26016 41148 26022 41160
rect 26973 41157 26985 41160
rect 27019 41157 27031 41191
rect 26973 41151 27031 41157
rect 28994 41148 29000 41200
rect 29052 41188 29058 41200
rect 30377 41191 30435 41197
rect 30377 41188 30389 41191
rect 29052 41160 30389 41188
rect 29052 41148 29058 41160
rect 30377 41157 30389 41160
rect 30423 41157 30435 41191
rect 30377 41151 30435 41157
rect 30834 41148 30840 41200
rect 30892 41188 30898 41200
rect 32370 41191 32428 41197
rect 32370 41188 32382 41191
rect 30892 41160 32382 41188
rect 30892 41148 30898 41160
rect 32370 41157 32382 41160
rect 32416 41157 32428 41191
rect 32370 41151 32428 41157
rect 34146 41148 34152 41200
rect 34204 41188 34210 41200
rect 36262 41188 36268 41200
rect 34204 41160 36268 41188
rect 34204 41148 34210 41160
rect 36262 41148 36268 41160
rect 36320 41148 36326 41200
rect 38470 41188 38476 41200
rect 38431 41160 38476 41188
rect 38470 41148 38476 41160
rect 38528 41148 38534 41200
rect 20257 41123 20315 41129
rect 20257 41089 20269 41123
rect 20303 41089 20315 41123
rect 20438 41120 20444 41132
rect 20399 41092 20444 41120
rect 20257 41083 20315 41089
rect 19720 41024 20208 41052
rect 19720 40984 19748 41024
rect 19260 40956 19748 40984
rect 20070 40944 20076 40996
rect 20128 40984 20134 40996
rect 20272 40984 20300 41083
rect 20438 41080 20444 41092
rect 20496 41080 20502 41132
rect 21818 41120 21824 41132
rect 21779 41092 21824 41120
rect 21818 41080 21824 41092
rect 21876 41080 21882 41132
rect 22005 41123 22063 41129
rect 22005 41120 22017 41123
rect 21928 41092 22017 41120
rect 21266 41012 21272 41064
rect 21324 41052 21330 41064
rect 21726 41052 21732 41064
rect 21324 41024 21732 41052
rect 21324 41012 21330 41024
rect 21726 41012 21732 41024
rect 21784 41052 21790 41064
rect 21928 41052 21956 41092
rect 22005 41089 22017 41092
rect 22051 41089 22063 41123
rect 22005 41083 22063 41089
rect 22189 41123 22247 41129
rect 22189 41089 22201 41123
rect 22235 41120 22247 41123
rect 22649 41123 22707 41129
rect 22649 41120 22661 41123
rect 22235 41092 22661 41120
rect 22235 41089 22247 41092
rect 22189 41083 22247 41089
rect 22649 41089 22661 41092
rect 22695 41089 22707 41123
rect 22649 41083 22707 41089
rect 22738 41080 22744 41132
rect 22796 41120 22802 41132
rect 22833 41123 22891 41129
rect 22833 41120 22845 41123
rect 22796 41092 22845 41120
rect 22796 41080 22802 41092
rect 22833 41089 22845 41092
rect 22879 41089 22891 41123
rect 24394 41120 24400 41132
rect 24355 41092 24400 41120
rect 22833 41083 22891 41089
rect 24394 41080 24400 41092
rect 24452 41080 24458 41132
rect 24486 41080 24492 41132
rect 24544 41120 24550 41132
rect 24673 41123 24731 41129
rect 24544 41092 24589 41120
rect 24544 41080 24550 41092
rect 24673 41089 24685 41123
rect 24719 41120 24731 41123
rect 24946 41120 24952 41132
rect 24719 41092 24952 41120
rect 24719 41089 24731 41092
rect 24673 41083 24731 41089
rect 24946 41080 24952 41092
rect 25004 41080 25010 41132
rect 25222 41080 25228 41132
rect 25280 41120 25286 41132
rect 25409 41123 25467 41129
rect 25409 41120 25421 41123
rect 25280 41092 25421 41120
rect 25280 41080 25286 41092
rect 25409 41089 25421 41092
rect 25455 41120 25467 41123
rect 25774 41120 25780 41132
rect 25455 41092 25780 41120
rect 25455 41089 25467 41092
rect 25409 41083 25467 41089
rect 25774 41080 25780 41092
rect 25832 41080 25838 41132
rect 29086 41080 29092 41132
rect 29144 41120 29150 41132
rect 32122 41120 32128 41132
rect 29144 41092 32128 41120
rect 29144 41080 29150 41092
rect 32122 41080 32128 41092
rect 32180 41080 32186 41132
rect 32674 41080 32680 41132
rect 32732 41120 32738 41132
rect 34057 41123 34115 41129
rect 34057 41120 34069 41123
rect 32732 41092 34069 41120
rect 32732 41080 32738 41092
rect 34057 41089 34069 41092
rect 34103 41089 34115 41123
rect 34057 41083 34115 41089
rect 34698 41080 34704 41132
rect 34756 41120 34762 41132
rect 34793 41123 34851 41129
rect 34793 41120 34805 41123
rect 34756 41092 34805 41120
rect 34756 41080 34762 41092
rect 34793 41089 34805 41092
rect 34839 41089 34851 41123
rect 34793 41083 34851 41089
rect 34977 41123 35035 41129
rect 34977 41089 34989 41123
rect 35023 41089 35035 41123
rect 34977 41083 35035 41089
rect 35713 41123 35771 41129
rect 35713 41089 35725 41123
rect 35759 41089 35771 41123
rect 35713 41083 35771 41089
rect 21784 41024 21956 41052
rect 21784 41012 21790 41024
rect 23842 41012 23848 41064
rect 23900 41052 23906 41064
rect 23900 41024 25452 41052
rect 23900 41012 23906 41024
rect 25424 40996 25452 41024
rect 25498 41012 25504 41064
rect 25556 41052 25562 41064
rect 25685 41055 25743 41061
rect 25685 41052 25697 41055
rect 25556 41024 25697 41052
rect 25556 41012 25562 41024
rect 25685 41021 25697 41024
rect 25731 41021 25743 41055
rect 25685 41015 25743 41021
rect 34333 41055 34391 41061
rect 34333 41021 34345 41055
rect 34379 41052 34391 41055
rect 34514 41052 34520 41064
rect 34379 41024 34520 41052
rect 34379 41021 34391 41024
rect 34333 41015 34391 41021
rect 34514 41012 34520 41024
rect 34572 41052 34578 41064
rect 34882 41052 34888 41064
rect 34572 41024 34888 41052
rect 34572 41012 34578 41024
rect 34882 41012 34888 41024
rect 34940 41012 34946 41064
rect 24026 40984 24032 40996
rect 20128 40956 24032 40984
rect 20128 40944 20134 40956
rect 24026 40944 24032 40956
rect 24084 40944 24090 40996
rect 24670 40984 24676 40996
rect 24631 40956 24676 40984
rect 24670 40944 24676 40956
rect 24728 40944 24734 40996
rect 25406 40944 25412 40996
rect 25464 40944 25470 40996
rect 25593 40987 25651 40993
rect 25593 40953 25605 40987
rect 25639 40984 25651 40987
rect 28994 40984 29000 40996
rect 25639 40956 29000 40984
rect 25639 40953 25651 40956
rect 25593 40947 25651 40953
rect 28994 40944 29000 40956
rect 29052 40944 29058 40996
rect 34992 40984 35020 41083
rect 35728 41052 35756 41083
rect 35802 41080 35808 41132
rect 35860 41120 35866 41132
rect 36449 41123 36507 41129
rect 36449 41120 36461 41123
rect 35860 41092 36461 41120
rect 35860 41080 35866 41092
rect 36449 41089 36461 41092
rect 36495 41089 36507 41123
rect 36449 41083 36507 41089
rect 36633 41123 36691 41129
rect 36633 41089 36645 41123
rect 36679 41120 36691 41123
rect 37734 41120 37740 41132
rect 36679 41092 37740 41120
rect 36679 41089 36691 41092
rect 36633 41083 36691 41089
rect 37734 41080 37740 41092
rect 37792 41080 37798 41132
rect 37826 41080 37832 41132
rect 37884 41120 37890 41132
rect 38289 41123 38347 41129
rect 38289 41120 38301 41123
rect 37884 41092 38301 41120
rect 37884 41080 37890 41092
rect 38289 41089 38301 41092
rect 38335 41120 38347 41123
rect 38562 41120 38568 41132
rect 38335 41092 38568 41120
rect 38335 41089 38347 41092
rect 38289 41083 38347 41089
rect 38562 41080 38568 41092
rect 38620 41080 38626 41132
rect 35894 41052 35900 41064
rect 35728 41024 35900 41052
rect 35894 41012 35900 41024
rect 35952 41012 35958 41064
rect 35989 41055 36047 41061
rect 35989 41021 36001 41055
rect 36035 41052 36047 41055
rect 36078 41052 36084 41064
rect 36035 41024 36084 41052
rect 36035 41021 36047 41024
rect 35989 41015 36047 41021
rect 36078 41012 36084 41024
rect 36136 41012 36142 41064
rect 36170 41012 36176 41064
rect 36228 41052 36234 41064
rect 40221 41055 40279 41061
rect 40221 41052 40233 41055
rect 36228 41024 40233 41052
rect 36228 41012 36234 41024
rect 40221 41021 40233 41024
rect 40267 41021 40279 41055
rect 40221 41015 40279 41021
rect 35342 40984 35348 40996
rect 29196 40956 31754 40984
rect 34992 40956 35348 40984
rect 13596 40888 17172 40916
rect 18693 40919 18751 40925
rect 13596 40876 13602 40888
rect 18693 40885 18705 40919
rect 18739 40916 18751 40919
rect 19150 40916 19156 40928
rect 18739 40888 19156 40916
rect 18739 40885 18751 40888
rect 18693 40879 18751 40885
rect 19150 40876 19156 40888
rect 19208 40876 19214 40928
rect 19242 40876 19248 40928
rect 19300 40916 19306 40928
rect 24578 40916 24584 40928
rect 19300 40888 24584 40916
rect 19300 40876 19306 40888
rect 24578 40876 24584 40888
rect 24636 40876 24642 40928
rect 24762 40876 24768 40928
rect 24820 40916 24826 40928
rect 25501 40919 25559 40925
rect 25501 40916 25513 40919
rect 24820 40888 25513 40916
rect 24820 40876 24826 40888
rect 25501 40885 25513 40888
rect 25547 40885 25559 40919
rect 25501 40879 25559 40885
rect 27062 40876 27068 40928
rect 27120 40916 27126 40928
rect 29196 40916 29224 40956
rect 27120 40888 29224 40916
rect 27120 40876 27126 40888
rect 30558 40876 30564 40928
rect 30616 40916 30622 40928
rect 30837 40919 30895 40925
rect 30837 40916 30849 40919
rect 30616 40888 30849 40916
rect 30616 40876 30622 40888
rect 30837 40885 30849 40888
rect 30883 40885 30895 40919
rect 30837 40879 30895 40885
rect 31294 40876 31300 40928
rect 31352 40916 31358 40928
rect 31389 40919 31447 40925
rect 31389 40916 31401 40919
rect 31352 40888 31401 40916
rect 31352 40876 31358 40888
rect 31389 40885 31401 40888
rect 31435 40885 31447 40919
rect 31726 40916 31754 40956
rect 35342 40944 35348 40956
rect 35400 40984 35406 40996
rect 37826 40984 37832 40996
rect 35400 40956 37832 40984
rect 35400 40944 35406 40956
rect 37826 40944 37832 40956
rect 37884 40944 37890 40996
rect 39209 40987 39267 40993
rect 39209 40953 39221 40987
rect 39255 40984 39267 40987
rect 40034 40984 40040 40996
rect 39255 40956 40040 40984
rect 39255 40953 39267 40956
rect 39209 40947 39267 40953
rect 40034 40944 40040 40956
rect 40092 40944 40098 40996
rect 33226 40916 33232 40928
rect 31726 40888 33232 40916
rect 31389 40879 31447 40885
rect 33226 40876 33232 40888
rect 33284 40876 33290 40928
rect 33502 40916 33508 40928
rect 33463 40888 33508 40916
rect 33502 40876 33508 40888
rect 33560 40876 33566 40928
rect 34146 40916 34152 40928
rect 34107 40888 34152 40916
rect 34146 40876 34152 40888
rect 34204 40876 34210 40928
rect 34790 40876 34796 40928
rect 34848 40916 34854 40928
rect 34885 40919 34943 40925
rect 34885 40916 34897 40919
rect 34848 40888 34897 40916
rect 34848 40876 34854 40888
rect 34885 40885 34897 40888
rect 34931 40885 34943 40919
rect 35802 40916 35808 40928
rect 35763 40888 35808 40916
rect 34885 40879 34943 40885
rect 35802 40876 35808 40888
rect 35860 40876 35866 40928
rect 35894 40876 35900 40928
rect 35952 40916 35958 40928
rect 37274 40916 37280 40928
rect 35952 40888 35997 40916
rect 37235 40888 37280 40916
rect 35952 40876 35958 40888
rect 37274 40876 37280 40888
rect 37332 40876 37338 40928
rect 39666 40916 39672 40928
rect 39627 40888 39672 40916
rect 39666 40876 39672 40888
rect 39724 40876 39730 40928
rect 41417 40919 41475 40925
rect 41417 40885 41429 40919
rect 41463 40916 41475 40919
rect 43162 40916 43168 40928
rect 41463 40888 43168 40916
rect 41463 40885 41475 40888
rect 41417 40879 41475 40885
rect 43162 40876 43168 40888
rect 43220 40876 43226 40928
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 12437 40715 12495 40721
rect 12437 40681 12449 40715
rect 12483 40712 12495 40715
rect 12710 40712 12716 40724
rect 12483 40684 12716 40712
rect 12483 40681 12495 40684
rect 12437 40675 12495 40681
rect 12710 40672 12716 40684
rect 12768 40672 12774 40724
rect 12894 40712 12900 40724
rect 12855 40684 12900 40712
rect 12894 40672 12900 40684
rect 12952 40672 12958 40724
rect 13541 40715 13599 40721
rect 13541 40681 13553 40715
rect 13587 40712 13599 40715
rect 13814 40712 13820 40724
rect 13587 40684 13820 40712
rect 13587 40681 13599 40684
rect 13541 40675 13599 40681
rect 12066 40604 12072 40656
rect 12124 40644 12130 40656
rect 13556 40644 13584 40675
rect 13814 40672 13820 40684
rect 13872 40672 13878 40724
rect 15562 40672 15568 40724
rect 15620 40712 15626 40724
rect 15841 40715 15899 40721
rect 15841 40712 15853 40715
rect 15620 40684 15853 40712
rect 15620 40672 15626 40684
rect 15841 40681 15853 40684
rect 15887 40681 15899 40715
rect 15841 40675 15899 40681
rect 16485 40715 16543 40721
rect 16485 40681 16497 40715
rect 16531 40712 16543 40715
rect 17862 40712 17868 40724
rect 16531 40684 17868 40712
rect 16531 40681 16543 40684
rect 16485 40675 16543 40681
rect 17862 40672 17868 40684
rect 17920 40672 17926 40724
rect 18690 40712 18696 40724
rect 18651 40684 18696 40712
rect 18690 40672 18696 40684
rect 18748 40672 18754 40724
rect 18782 40672 18788 40724
rect 18840 40712 18846 40724
rect 19426 40712 19432 40724
rect 18840 40684 19432 40712
rect 18840 40672 18846 40684
rect 19426 40672 19432 40684
rect 19484 40672 19490 40724
rect 19797 40715 19855 40721
rect 19797 40681 19809 40715
rect 19843 40712 19855 40715
rect 20070 40712 20076 40724
rect 19843 40684 20076 40712
rect 19843 40681 19855 40684
rect 19797 40675 19855 40681
rect 20070 40672 20076 40684
rect 20128 40672 20134 40724
rect 20441 40715 20499 40721
rect 20441 40712 20453 40715
rect 20180 40684 20453 40712
rect 15194 40644 15200 40656
rect 12124 40616 13584 40644
rect 15107 40616 15200 40644
rect 12124 40604 12130 40616
rect 15194 40604 15200 40616
rect 15252 40644 15258 40656
rect 17586 40644 17592 40656
rect 15252 40616 17592 40644
rect 15252 40604 15258 40616
rect 17586 40604 17592 40616
rect 17644 40604 17650 40656
rect 18414 40604 18420 40656
rect 18472 40644 18478 40656
rect 19518 40644 19524 40656
rect 18472 40616 19524 40644
rect 18472 40604 18478 40616
rect 19518 40604 19524 40616
rect 19576 40644 19582 40656
rect 20180 40644 20208 40684
rect 20441 40681 20453 40684
rect 20487 40681 20499 40715
rect 20441 40675 20499 40681
rect 22281 40715 22339 40721
rect 22281 40681 22293 40715
rect 22327 40712 22339 40715
rect 24762 40712 24768 40724
rect 22327 40684 24768 40712
rect 22327 40681 22339 40684
rect 22281 40675 22339 40681
rect 24762 40672 24768 40684
rect 24820 40672 24826 40724
rect 24946 40712 24952 40724
rect 24872 40684 24952 40712
rect 19576 40616 20208 40644
rect 20257 40647 20315 40653
rect 19576 40604 19582 40616
rect 20257 40613 20269 40647
rect 20303 40613 20315 40647
rect 22833 40647 22891 40653
rect 22833 40644 22845 40647
rect 20257 40607 20315 40613
rect 22020 40616 22845 40644
rect 12710 40536 12716 40588
rect 12768 40576 12774 40588
rect 18322 40576 18328 40588
rect 12768 40548 18328 40576
rect 12768 40536 12774 40548
rect 11885 40511 11943 40517
rect 11885 40477 11897 40511
rect 11931 40508 11943 40511
rect 15010 40508 15016 40520
rect 11931 40480 15016 40508
rect 11931 40477 11943 40480
rect 11885 40471 11943 40477
rect 15010 40468 15016 40480
rect 15068 40468 15074 40520
rect 15102 40468 15108 40520
rect 15160 40508 15166 40520
rect 15749 40511 15807 40517
rect 15749 40508 15761 40511
rect 15160 40480 15761 40508
rect 15160 40468 15166 40480
rect 15749 40477 15761 40480
rect 15795 40477 15807 40511
rect 15749 40471 15807 40477
rect 16574 40468 16580 40520
rect 16632 40508 16638 40520
rect 17589 40511 17647 40517
rect 17589 40508 17601 40511
rect 16632 40480 17601 40508
rect 16632 40468 16638 40480
rect 17589 40477 17601 40480
rect 17635 40508 17647 40511
rect 17862 40508 17868 40520
rect 17635 40480 17868 40508
rect 17635 40477 17647 40480
rect 17589 40471 17647 40477
rect 17862 40468 17868 40480
rect 17920 40468 17926 40520
rect 17972 40508 18000 40548
rect 18322 40536 18328 40548
rect 18380 40536 18386 40588
rect 19058 40536 19064 40588
rect 19116 40576 19122 40588
rect 19245 40579 19303 40585
rect 19245 40576 19257 40579
rect 19116 40548 19257 40576
rect 19116 40536 19122 40548
rect 19245 40545 19257 40548
rect 19291 40545 19303 40579
rect 19794 40576 19800 40588
rect 19245 40539 19303 40545
rect 19536 40548 19800 40576
rect 18038 40511 18096 40517
rect 18038 40508 18050 40511
rect 17972 40480 18050 40508
rect 18038 40477 18050 40480
rect 18084 40477 18096 40511
rect 18038 40471 18096 40477
rect 18138 40468 18144 40520
rect 18196 40508 18202 40520
rect 18196 40480 18241 40508
rect 18196 40468 18202 40480
rect 18506 40468 18512 40520
rect 18564 40517 18570 40520
rect 18564 40508 18572 40517
rect 18564 40480 18609 40508
rect 18564 40471 18572 40480
rect 18564 40468 18570 40471
rect 18874 40468 18880 40520
rect 18932 40508 18938 40520
rect 19536 40517 19564 40548
rect 19794 40536 19800 40548
rect 19852 40536 19858 40588
rect 20070 40536 20076 40588
rect 20128 40576 20134 40588
rect 20272 40576 20300 40607
rect 22020 40585 22048 40616
rect 22833 40613 22845 40616
rect 22879 40613 22891 40647
rect 23842 40644 23848 40656
rect 23803 40616 23848 40644
rect 22833 40607 22891 40613
rect 23842 40604 23848 40616
rect 23900 40604 23906 40656
rect 20128 40548 20300 40576
rect 22005 40579 22063 40585
rect 20128 40536 20134 40548
rect 22005 40545 22017 40579
rect 22051 40545 22063 40579
rect 22738 40576 22744 40588
rect 22651 40548 22744 40576
rect 22005 40539 22063 40545
rect 22738 40536 22744 40548
rect 22796 40536 22802 40588
rect 24872 40576 24900 40684
rect 24946 40672 24952 40684
rect 25004 40672 25010 40724
rect 25133 40715 25191 40721
rect 25133 40681 25145 40715
rect 25179 40712 25191 40715
rect 25682 40712 25688 40724
rect 25179 40684 25688 40712
rect 25179 40681 25191 40684
rect 25133 40675 25191 40681
rect 25682 40672 25688 40684
rect 25740 40672 25746 40724
rect 25777 40715 25835 40721
rect 25777 40681 25789 40715
rect 25823 40681 25835 40715
rect 25777 40675 25835 40681
rect 23860 40548 24900 40576
rect 25792 40576 25820 40675
rect 25958 40672 25964 40724
rect 26016 40712 26022 40724
rect 27062 40712 27068 40724
rect 26016 40684 27068 40712
rect 26016 40672 26022 40684
rect 27062 40672 27068 40684
rect 27120 40672 27126 40724
rect 28905 40715 28963 40721
rect 28905 40681 28917 40715
rect 28951 40712 28963 40715
rect 32401 40715 32459 40721
rect 32401 40712 32413 40715
rect 28951 40684 32413 40712
rect 28951 40681 28963 40684
rect 28905 40675 28963 40681
rect 32401 40681 32413 40684
rect 32447 40712 32459 40715
rect 32490 40712 32496 40724
rect 32447 40684 32496 40712
rect 32447 40681 32459 40684
rect 32401 40675 32459 40681
rect 32490 40672 32496 40684
rect 32548 40672 32554 40724
rect 32585 40715 32643 40721
rect 32585 40681 32597 40715
rect 32631 40712 32643 40715
rect 32674 40712 32680 40724
rect 32631 40684 32680 40712
rect 32631 40681 32643 40684
rect 32585 40675 32643 40681
rect 32674 40672 32680 40684
rect 32732 40672 32738 40724
rect 34146 40712 34152 40724
rect 34107 40684 34152 40712
rect 34146 40672 34152 40684
rect 34204 40672 34210 40724
rect 35986 40672 35992 40724
rect 36044 40712 36050 40724
rect 37090 40712 37096 40724
rect 36044 40684 37096 40712
rect 36044 40672 36050 40684
rect 37090 40672 37096 40684
rect 37148 40672 37154 40724
rect 37734 40712 37740 40724
rect 37695 40684 37740 40712
rect 37734 40672 37740 40684
rect 37792 40672 37798 40724
rect 40218 40672 40224 40724
rect 40276 40712 40282 40724
rect 40405 40715 40463 40721
rect 40405 40712 40417 40715
rect 40276 40684 40417 40712
rect 40276 40672 40282 40684
rect 40405 40681 40417 40684
rect 40451 40681 40463 40715
rect 40405 40675 40463 40681
rect 25866 40604 25872 40656
rect 25924 40644 25930 40656
rect 26697 40647 26755 40653
rect 26697 40644 26709 40647
rect 25924 40616 26709 40644
rect 25924 40604 25930 40616
rect 26697 40613 26709 40616
rect 26743 40613 26755 40647
rect 26697 40607 26755 40613
rect 30929 40647 30987 40653
rect 30929 40613 30941 40647
rect 30975 40644 30987 40647
rect 32306 40644 32312 40656
rect 30975 40616 32312 40644
rect 30975 40613 30987 40616
rect 30929 40607 30987 40613
rect 32306 40604 32312 40616
rect 32364 40604 32370 40656
rect 33870 40604 33876 40656
rect 33928 40644 33934 40656
rect 34422 40644 34428 40656
rect 33928 40616 34428 40644
rect 33928 40604 33934 40616
rect 34422 40604 34428 40616
rect 34480 40604 34486 40656
rect 36170 40604 36176 40656
rect 36228 40644 36234 40656
rect 41046 40644 41052 40656
rect 36228 40616 41052 40644
rect 36228 40604 36234 40616
rect 41046 40604 41052 40616
rect 41104 40604 41110 40656
rect 26326 40576 26332 40588
rect 25792 40548 26332 40576
rect 19521 40511 19579 40517
rect 18932 40502 19196 40508
rect 19521 40502 19533 40511
rect 18932 40480 19533 40502
rect 18932 40468 18938 40480
rect 19168 40477 19533 40480
rect 19567 40477 19579 40511
rect 19168 40474 19579 40477
rect 19521 40471 19579 40474
rect 19613 40511 19671 40517
rect 19613 40477 19625 40511
rect 19659 40502 19671 40511
rect 20530 40508 20536 40520
rect 19720 40502 20536 40508
rect 19659 40480 20536 40502
rect 19659 40477 19748 40480
rect 19613 40474 19748 40477
rect 19613 40471 19671 40474
rect 20530 40468 20536 40480
rect 20588 40468 20594 40520
rect 21082 40508 21088 40520
rect 21043 40480 21088 40508
rect 21082 40468 21088 40480
rect 21140 40468 21146 40520
rect 21266 40508 21272 40520
rect 21227 40480 21272 40508
rect 21266 40468 21272 40480
rect 21324 40468 21330 40520
rect 21910 40508 21916 40520
rect 21871 40480 21916 40508
rect 21910 40468 21916 40480
rect 21968 40468 21974 40520
rect 22756 40508 22784 40536
rect 22066 40480 22784 40508
rect 22925 40511 22983 40517
rect 1578 40400 1584 40452
rect 1636 40440 1642 40452
rect 1857 40443 1915 40449
rect 1857 40440 1869 40443
rect 1636 40412 1869 40440
rect 1636 40400 1642 40412
rect 1857 40409 1869 40412
rect 1903 40409 1915 40443
rect 2038 40440 2044 40452
rect 1999 40412 2044 40440
rect 1857 40403 1915 40409
rect 2038 40400 2044 40412
rect 2096 40400 2102 40452
rect 18322 40440 18328 40452
rect 18283 40412 18328 40440
rect 18322 40400 18328 40412
rect 18380 40400 18386 40452
rect 18417 40443 18475 40449
rect 18417 40409 18429 40443
rect 18463 40440 18475 40443
rect 18782 40440 18788 40452
rect 18463 40412 18788 40440
rect 18463 40409 18475 40412
rect 18417 40403 18475 40409
rect 18782 40400 18788 40412
rect 18840 40400 18846 40452
rect 20625 40443 20683 40449
rect 20625 40440 20637 40443
rect 19352 40412 20637 40440
rect 13998 40332 14004 40384
rect 14056 40372 14062 40384
rect 14461 40375 14519 40381
rect 14461 40372 14473 40375
rect 14056 40344 14473 40372
rect 14056 40332 14062 40344
rect 14461 40341 14473 40344
rect 14507 40372 14519 40375
rect 15286 40372 15292 40384
rect 14507 40344 15292 40372
rect 14507 40341 14519 40344
rect 14461 40335 14519 40341
rect 15286 40332 15292 40344
rect 15344 40332 15350 40384
rect 17034 40372 17040 40384
rect 16995 40344 17040 40372
rect 17034 40332 17040 40344
rect 17092 40332 17098 40384
rect 19058 40332 19064 40384
rect 19116 40372 19122 40384
rect 19352 40372 19380 40412
rect 20625 40409 20637 40412
rect 20671 40409 20683 40443
rect 20625 40403 20683 40409
rect 21177 40443 21235 40449
rect 21177 40409 21189 40443
rect 21223 40440 21235 40443
rect 22066 40440 22094 40480
rect 22925 40477 22937 40511
rect 22971 40477 22983 40511
rect 22925 40471 22983 40477
rect 21223 40412 22094 40440
rect 21223 40409 21235 40412
rect 21177 40403 21235 40409
rect 22186 40400 22192 40452
rect 22244 40440 22250 40452
rect 22940 40440 22968 40471
rect 23014 40468 23020 40520
rect 23072 40508 23078 40520
rect 23569 40511 23627 40517
rect 23072 40480 23117 40508
rect 23072 40468 23078 40480
rect 23569 40477 23581 40511
rect 23615 40508 23627 40511
rect 23750 40508 23756 40520
rect 23615 40480 23756 40508
rect 23615 40477 23627 40480
rect 23569 40471 23627 40477
rect 23750 40468 23756 40480
rect 23808 40468 23814 40520
rect 23860 40517 23888 40548
rect 26326 40536 26332 40548
rect 26384 40576 26390 40588
rect 26384 40548 26740 40576
rect 26384 40536 26390 40548
rect 23845 40511 23903 40517
rect 23845 40477 23857 40511
rect 23891 40477 23903 40511
rect 23845 40471 23903 40477
rect 24210 40468 24216 40520
rect 24268 40508 24274 40520
rect 24489 40511 24547 40517
rect 24489 40508 24501 40511
rect 24268 40480 24501 40508
rect 24268 40468 24274 40480
rect 24489 40477 24501 40480
rect 24535 40477 24547 40511
rect 24489 40471 24547 40477
rect 24578 40468 24584 40520
rect 24636 40508 24642 40520
rect 25038 40517 25044 40520
rect 24993 40511 25044 40517
rect 24636 40480 24681 40508
rect 24636 40468 24642 40480
rect 24993 40477 25005 40511
rect 25039 40477 25044 40511
rect 24993 40471 25044 40477
rect 25038 40468 25044 40471
rect 25096 40468 25102 40520
rect 26712 40517 26740 40548
rect 27154 40536 27160 40588
rect 27212 40576 27218 40588
rect 27525 40579 27583 40585
rect 27525 40576 27537 40579
rect 27212 40548 27537 40576
rect 27212 40536 27218 40548
rect 27525 40545 27537 40548
rect 27571 40545 27583 40579
rect 27525 40539 27583 40545
rect 29086 40536 29092 40588
rect 29144 40576 29150 40588
rect 29549 40579 29607 40585
rect 29549 40576 29561 40579
rect 29144 40548 29561 40576
rect 29144 40536 29150 40548
rect 29549 40545 29561 40548
rect 29595 40545 29607 40579
rect 33318 40576 33324 40588
rect 29549 40539 29607 40545
rect 30576 40548 33324 40576
rect 26421 40511 26479 40517
rect 26421 40508 26433 40511
rect 25808 40480 26433 40508
rect 24762 40440 24768 40452
rect 22244 40412 22968 40440
rect 24723 40412 24768 40440
rect 22244 40400 22250 40412
rect 24762 40400 24768 40412
rect 24820 40400 24826 40452
rect 24854 40400 24860 40452
rect 24912 40440 24918 40452
rect 25590 40440 25596 40452
rect 24912 40412 24957 40440
rect 25551 40412 25596 40440
rect 24912 40400 24918 40412
rect 25590 40400 25596 40412
rect 25648 40400 25654 40452
rect 19116 40344 19380 40372
rect 19429 40375 19487 40381
rect 19116 40332 19122 40344
rect 19429 40341 19441 40375
rect 19475 40372 19487 40375
rect 19518 40372 19524 40384
rect 19475 40344 19524 40372
rect 19475 40341 19487 40344
rect 19429 40335 19487 40341
rect 19518 40332 19524 40344
rect 19576 40332 19582 40384
rect 19794 40332 19800 40384
rect 19852 40372 19858 40384
rect 20415 40375 20473 40381
rect 20415 40372 20427 40375
rect 19852 40344 20427 40372
rect 19852 40332 19858 40344
rect 20415 40341 20427 40344
rect 20461 40341 20473 40375
rect 23658 40372 23664 40384
rect 23619 40344 23664 40372
rect 20415 40335 20473 40341
rect 23658 40332 23664 40344
rect 23716 40332 23722 40384
rect 24026 40332 24032 40384
rect 24084 40372 24090 40384
rect 25808 40381 25836 40480
rect 26421 40477 26433 40480
rect 26467 40477 26479 40511
rect 26421 40471 26479 40477
rect 26697 40511 26755 40517
rect 26697 40477 26709 40511
rect 26743 40477 26755 40511
rect 26697 40471 26755 40477
rect 27792 40511 27850 40517
rect 27792 40477 27804 40511
rect 27838 40508 27850 40511
rect 30576 40508 30604 40548
rect 33318 40536 33324 40548
rect 33376 40536 33382 40588
rect 33413 40579 33471 40585
rect 33413 40545 33425 40579
rect 33459 40576 33471 40579
rect 33594 40576 33600 40588
rect 33459 40548 33600 40576
rect 33459 40545 33471 40548
rect 33413 40539 33471 40545
rect 33594 40536 33600 40548
rect 33652 40576 33658 40588
rect 34330 40576 34336 40588
rect 33652 40548 34336 40576
rect 33652 40536 33658 40548
rect 34330 40536 34336 40548
rect 34388 40536 34394 40588
rect 35802 40536 35808 40588
rect 35860 40576 35866 40588
rect 36357 40579 36415 40585
rect 36357 40576 36369 40579
rect 35860 40548 36369 40576
rect 35860 40536 35866 40548
rect 36357 40545 36369 40548
rect 36403 40545 36415 40579
rect 36357 40539 36415 40545
rect 36630 40536 36636 40588
rect 36688 40576 36694 40588
rect 38657 40579 38715 40585
rect 38657 40576 38669 40579
rect 36688 40548 38669 40576
rect 36688 40536 36694 40548
rect 38657 40545 38669 40548
rect 38703 40576 38715 40579
rect 39853 40579 39911 40585
rect 39853 40576 39865 40579
rect 38703 40548 39865 40576
rect 38703 40545 38715 40548
rect 38657 40539 38715 40545
rect 39853 40545 39865 40548
rect 39899 40576 39911 40579
rect 39899 40548 41414 40576
rect 39899 40545 39911 40548
rect 39853 40539 39911 40545
rect 27838 40480 30604 40508
rect 27838 40477 27850 40480
rect 27792 40471 27850 40477
rect 31754 40468 31760 40520
rect 31812 40508 31818 40520
rect 33226 40508 33232 40520
rect 31812 40480 31857 40508
rect 33187 40480 33232 40508
rect 31812 40468 31818 40480
rect 33226 40468 33232 40480
rect 33284 40468 33290 40520
rect 33873 40511 33931 40517
rect 33873 40477 33885 40511
rect 33919 40508 33931 40511
rect 34698 40508 34704 40520
rect 33919 40480 34704 40508
rect 33919 40477 33931 40480
rect 33873 40471 33931 40477
rect 26234 40400 26240 40452
rect 26292 40440 26298 40452
rect 26513 40443 26571 40449
rect 26513 40440 26525 40443
rect 26292 40412 26525 40440
rect 26292 40400 26298 40412
rect 26513 40409 26525 40412
rect 26559 40440 26571 40443
rect 27614 40440 27620 40452
rect 26559 40412 27620 40440
rect 26559 40409 26571 40412
rect 26513 40403 26571 40409
rect 27614 40400 27620 40412
rect 27672 40400 27678 40452
rect 29816 40443 29874 40449
rect 29816 40409 29828 40443
rect 29862 40440 29874 40443
rect 32217 40443 32275 40449
rect 29862 40412 31616 40440
rect 29862 40409 29874 40412
rect 29816 40403 29874 40409
rect 31588 40381 31616 40412
rect 32217 40409 32229 40443
rect 32263 40440 32275 40443
rect 32263 40412 32352 40440
rect 32263 40409 32275 40412
rect 32217 40403 32275 40409
rect 32324 40384 32352 40412
rect 32398 40400 32404 40452
rect 32456 40449 32462 40452
rect 32456 40443 32475 40449
rect 32463 40440 32475 40443
rect 33045 40443 33103 40449
rect 33045 40440 33057 40443
rect 32463 40412 33057 40440
rect 32463 40409 32475 40412
rect 32456 40403 32475 40409
rect 33045 40409 33057 40412
rect 33091 40440 33103 40443
rect 33888 40440 33916 40471
rect 34698 40468 34704 40480
rect 34756 40468 34762 40520
rect 34885 40511 34943 40517
rect 34885 40477 34897 40511
rect 34931 40508 34943 40511
rect 35342 40508 35348 40520
rect 34931 40480 35348 40508
rect 34931 40477 34943 40480
rect 34885 40471 34943 40477
rect 34146 40440 34152 40452
rect 33091 40412 33916 40440
rect 34107 40412 34152 40440
rect 33091 40409 33103 40412
rect 33045 40403 33103 40409
rect 32456 40400 32462 40403
rect 34146 40400 34152 40412
rect 34204 40400 34210 40452
rect 34900 40440 34928 40471
rect 35342 40468 35348 40480
rect 35400 40468 35406 40520
rect 35526 40508 35532 40520
rect 35487 40480 35532 40508
rect 35526 40468 35532 40480
rect 35584 40468 35590 40520
rect 35621 40511 35679 40517
rect 35621 40477 35633 40511
rect 35667 40508 35679 40511
rect 35894 40508 35900 40520
rect 35667 40480 35900 40508
rect 35667 40477 35679 40480
rect 35621 40471 35679 40477
rect 35894 40468 35900 40480
rect 35952 40468 35958 40520
rect 36265 40511 36323 40517
rect 36265 40477 36277 40511
rect 36311 40477 36323 40511
rect 36265 40471 36323 40477
rect 36449 40511 36507 40517
rect 36449 40477 36461 40511
rect 36495 40508 36507 40511
rect 37918 40508 37924 40520
rect 36495 40480 37924 40508
rect 36495 40477 36507 40480
rect 36449 40471 36507 40477
rect 35805 40443 35863 40449
rect 35805 40440 35817 40443
rect 34624 40412 34928 40440
rect 34992 40412 35817 40440
rect 25793 40375 25851 40381
rect 25793 40372 25805 40375
rect 24084 40344 25805 40372
rect 24084 40332 24090 40344
rect 25793 40341 25805 40344
rect 25839 40341 25851 40375
rect 25793 40335 25851 40341
rect 31573 40375 31631 40381
rect 31573 40341 31585 40375
rect 31619 40341 31631 40375
rect 31573 40335 31631 40341
rect 32306 40332 32312 40384
rect 32364 40372 32370 40384
rect 33965 40375 34023 40381
rect 33965 40372 33977 40375
rect 32364 40344 33977 40372
rect 32364 40332 32370 40344
rect 33965 40341 33977 40344
rect 34011 40372 34023 40375
rect 34624 40372 34652 40412
rect 34011 40344 34652 40372
rect 34011 40341 34023 40344
rect 33965 40335 34023 40341
rect 34698 40332 34704 40384
rect 34756 40372 34762 40384
rect 34992 40372 35020 40412
rect 35805 40409 35817 40412
rect 35851 40440 35863 40443
rect 36170 40440 36176 40452
rect 35851 40412 36176 40440
rect 35851 40409 35863 40412
rect 35805 40403 35863 40409
rect 36170 40400 36176 40412
rect 36228 40400 36234 40452
rect 34756 40344 35020 40372
rect 35069 40375 35127 40381
rect 34756 40332 34762 40344
rect 35069 40341 35081 40375
rect 35115 40372 35127 40375
rect 35342 40372 35348 40384
rect 35115 40344 35348 40372
rect 35115 40341 35127 40344
rect 35069 40335 35127 40341
rect 35342 40332 35348 40344
rect 35400 40332 35406 40384
rect 35434 40332 35440 40384
rect 35492 40372 35498 40384
rect 35706 40375 35764 40381
rect 35706 40372 35718 40375
rect 35492 40344 35718 40372
rect 35492 40332 35498 40344
rect 35706 40341 35718 40344
rect 35752 40341 35764 40375
rect 36280 40372 36308 40471
rect 37918 40468 37924 40480
rect 37976 40468 37982 40520
rect 38013 40511 38071 40517
rect 38013 40477 38025 40511
rect 38059 40477 38071 40511
rect 38013 40471 38071 40477
rect 36906 40440 36912 40452
rect 36867 40412 36912 40440
rect 36906 40400 36912 40412
rect 36964 40400 36970 40452
rect 37090 40440 37096 40452
rect 37051 40412 37096 40440
rect 37090 40400 37096 40412
rect 37148 40400 37154 40452
rect 38028 40440 38056 40471
rect 41386 40440 41414 40548
rect 47857 40511 47915 40517
rect 47857 40508 47869 40511
rect 47320 40480 47869 40508
rect 47320 40452 47348 40480
rect 47857 40477 47869 40480
rect 47903 40477 47915 40511
rect 47857 40471 47915 40477
rect 41598 40440 41604 40452
rect 37476 40412 38056 40440
rect 39684 40412 41184 40440
rect 41386 40412 41604 40440
rect 37476 40384 37504 40412
rect 39684 40384 39712 40412
rect 37277 40375 37335 40381
rect 37277 40372 37289 40375
rect 36280 40344 37289 40372
rect 35706 40335 35764 40341
rect 37277 40341 37289 40344
rect 37323 40372 37335 40375
rect 37458 40372 37464 40384
rect 37323 40344 37464 40372
rect 37323 40341 37335 40344
rect 37277 40335 37335 40341
rect 37458 40332 37464 40344
rect 37516 40332 37522 40384
rect 38654 40332 38660 40384
rect 38712 40372 38718 40384
rect 39117 40375 39175 40381
rect 39117 40372 39129 40375
rect 38712 40344 39129 40372
rect 38712 40332 38718 40344
rect 39117 40341 39129 40344
rect 39163 40372 39175 40375
rect 39666 40372 39672 40384
rect 39163 40344 39672 40372
rect 39163 40341 39175 40344
rect 39117 40335 39175 40341
rect 39666 40332 39672 40344
rect 39724 40332 39730 40384
rect 41046 40372 41052 40384
rect 41007 40344 41052 40372
rect 41046 40332 41052 40344
rect 41104 40332 41110 40384
rect 41156 40372 41184 40412
rect 41598 40400 41604 40412
rect 41656 40400 41662 40452
rect 47302 40440 47308 40452
rect 47263 40412 47308 40440
rect 47302 40400 47308 40412
rect 47360 40400 47366 40452
rect 41506 40372 41512 40384
rect 41156 40344 41512 40372
rect 41506 40332 41512 40344
rect 41564 40332 41570 40384
rect 42058 40372 42064 40384
rect 42019 40344 42064 40372
rect 42058 40332 42064 40344
rect 42116 40332 42122 40384
rect 48038 40372 48044 40384
rect 47999 40344 48044 40372
rect 48038 40332 48044 40344
rect 48096 40332 48102 40384
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 1578 40168 1584 40180
rect 1539 40140 1584 40168
rect 1578 40128 1584 40140
rect 1636 40128 1642 40180
rect 13817 40171 13875 40177
rect 13817 40137 13829 40171
rect 13863 40168 13875 40171
rect 13906 40168 13912 40180
rect 13863 40140 13912 40168
rect 13863 40137 13875 40140
rect 13817 40131 13875 40137
rect 13906 40128 13912 40140
rect 13964 40168 13970 40180
rect 14826 40168 14832 40180
rect 13964 40140 14832 40168
rect 13964 40128 13970 40140
rect 14826 40128 14832 40140
rect 14884 40168 14890 40180
rect 15470 40168 15476 40180
rect 14884 40140 15476 40168
rect 14884 40128 14890 40140
rect 15470 40128 15476 40140
rect 15528 40128 15534 40180
rect 17034 40128 17040 40180
rect 17092 40168 17098 40180
rect 20254 40168 20260 40180
rect 17092 40140 20260 40168
rect 17092 40128 17098 40140
rect 20254 40128 20260 40140
rect 20312 40128 20318 40180
rect 23109 40171 23167 40177
rect 23109 40137 23121 40171
rect 23155 40168 23167 40171
rect 23198 40168 23204 40180
rect 23155 40140 23204 40168
rect 23155 40137 23167 40140
rect 23109 40131 23167 40137
rect 23198 40128 23204 40140
rect 23256 40128 23262 40180
rect 23477 40171 23535 40177
rect 23477 40137 23489 40171
rect 23523 40168 23535 40171
rect 23658 40168 23664 40180
rect 23523 40140 23664 40168
rect 23523 40137 23535 40140
rect 23477 40131 23535 40137
rect 23658 40128 23664 40140
rect 23716 40128 23722 40180
rect 24489 40171 24547 40177
rect 24489 40137 24501 40171
rect 24535 40168 24547 40171
rect 24762 40168 24768 40180
rect 24535 40140 24768 40168
rect 24535 40137 24547 40140
rect 24489 40131 24547 40137
rect 24762 40128 24768 40140
rect 24820 40128 24826 40180
rect 25498 40168 25504 40180
rect 25459 40140 25504 40168
rect 25498 40128 25504 40140
rect 25556 40128 25562 40180
rect 26142 40168 26148 40180
rect 25608 40140 26148 40168
rect 25608 40112 25636 40140
rect 26142 40128 26148 40140
rect 26200 40128 26206 40180
rect 27150 40171 27208 40177
rect 27150 40137 27162 40171
rect 27196 40168 27208 40171
rect 27246 40168 27252 40180
rect 27196 40140 27252 40168
rect 27196 40137 27208 40140
rect 27150 40131 27208 40137
rect 27246 40128 27252 40140
rect 27304 40128 27310 40180
rect 35526 40168 35532 40180
rect 35487 40140 35532 40168
rect 35526 40128 35532 40140
rect 35584 40128 35590 40180
rect 35986 40128 35992 40180
rect 36044 40128 36050 40180
rect 36633 40171 36691 40177
rect 36633 40137 36645 40171
rect 36679 40168 36691 40171
rect 36906 40168 36912 40180
rect 36679 40140 36912 40168
rect 36679 40137 36691 40140
rect 36633 40131 36691 40137
rect 36906 40128 36912 40140
rect 36964 40128 36970 40180
rect 38742 40171 38800 40177
rect 38742 40168 38754 40171
rect 37752 40140 38754 40168
rect 11790 40060 11796 40112
rect 11848 40100 11854 40112
rect 12710 40100 12716 40112
rect 11848 40072 12716 40100
rect 11848 40060 11854 40072
rect 12710 40060 12716 40072
rect 12768 40100 12774 40112
rect 13265 40103 13323 40109
rect 13265 40100 13277 40103
rect 12768 40072 13277 40100
rect 12768 40060 12774 40072
rect 13265 40069 13277 40072
rect 13311 40100 13323 40103
rect 17218 40100 17224 40112
rect 13311 40072 17224 40100
rect 13311 40069 13323 40072
rect 13265 40063 13323 40069
rect 17218 40060 17224 40072
rect 17276 40060 17282 40112
rect 17586 40100 17592 40112
rect 17328 40072 17592 40100
rect 12066 40032 12072 40044
rect 12027 40004 12072 40032
rect 12066 39992 12072 40004
rect 12124 39992 12130 40044
rect 12434 39992 12440 40044
rect 12492 40032 12498 40044
rect 12621 40035 12679 40041
rect 12621 40032 12633 40035
rect 12492 40004 12633 40032
rect 12492 39992 12498 40004
rect 12621 40001 12633 40004
rect 12667 40001 12679 40035
rect 12621 39995 12679 40001
rect 14461 40035 14519 40041
rect 14461 40001 14473 40035
rect 14507 40032 14519 40035
rect 14642 40032 14648 40044
rect 14507 40004 14648 40032
rect 14507 40001 14519 40004
rect 14461 39995 14519 40001
rect 14642 39992 14648 40004
rect 14700 39992 14706 40044
rect 17328 40041 17356 40072
rect 17586 40060 17592 40072
rect 17644 40060 17650 40112
rect 19150 40100 19156 40112
rect 19111 40072 19156 40100
rect 19150 40060 19156 40072
rect 19208 40060 19214 40112
rect 19334 40060 19340 40112
rect 19392 40100 19398 40112
rect 20070 40100 20076 40112
rect 19392 40072 20076 40100
rect 19392 40060 19398 40072
rect 20070 40060 20076 40072
rect 20128 40060 20134 40112
rect 20530 40100 20536 40112
rect 20491 40072 20536 40100
rect 20530 40060 20536 40072
rect 20588 40060 20594 40112
rect 23934 40060 23940 40112
rect 23992 40100 23998 40112
rect 25590 40100 25596 40112
rect 23992 40072 25596 40100
rect 23992 40060 23998 40072
rect 17313 40035 17371 40041
rect 17313 40001 17325 40035
rect 17359 40001 17371 40035
rect 17313 39995 17371 40001
rect 20257 40035 20315 40041
rect 20257 40001 20269 40035
rect 20303 40001 20315 40035
rect 20257 39995 20315 40001
rect 14274 39924 14280 39976
rect 14332 39964 14338 39976
rect 14369 39967 14427 39973
rect 14369 39964 14381 39967
rect 14332 39936 14381 39964
rect 14332 39924 14338 39936
rect 14369 39933 14381 39936
rect 14415 39933 14427 39967
rect 14369 39927 14427 39933
rect 14829 39967 14887 39973
rect 14829 39933 14841 39967
rect 14875 39964 14887 39967
rect 17034 39964 17040 39976
rect 14875 39936 17040 39964
rect 14875 39933 14887 39936
rect 14829 39927 14887 39933
rect 17034 39924 17040 39936
rect 17092 39924 17098 39976
rect 17126 39924 17132 39976
rect 17184 39964 17190 39976
rect 17221 39967 17279 39973
rect 17221 39964 17233 39967
rect 17184 39936 17233 39964
rect 17184 39924 17190 39936
rect 17221 39933 17233 39936
rect 17267 39933 17279 39967
rect 17221 39927 17279 39933
rect 17402 39924 17408 39976
rect 17460 39964 17466 39976
rect 18874 39964 18880 39976
rect 17460 39936 18880 39964
rect 17460 39924 17466 39936
rect 18874 39924 18880 39936
rect 18932 39924 18938 39976
rect 18969 39967 19027 39973
rect 18969 39933 18981 39967
rect 19015 39964 19027 39967
rect 19978 39964 19984 39976
rect 19015 39936 19984 39964
rect 19015 39933 19027 39936
rect 18969 39927 19027 39933
rect 19978 39924 19984 39936
rect 20036 39924 20042 39976
rect 20272 39964 20300 39995
rect 20346 39992 20352 40044
rect 20404 40032 20410 40044
rect 20993 40035 21051 40041
rect 20404 40004 20449 40032
rect 20404 39992 20410 40004
rect 20993 40001 21005 40035
rect 21039 40001 21051 40035
rect 21174 40032 21180 40044
rect 21135 40004 21180 40032
rect 20993 39995 21051 40001
rect 20622 39964 20628 39976
rect 20272 39936 20628 39964
rect 20622 39924 20628 39936
rect 20680 39924 20686 39976
rect 14182 39856 14188 39908
rect 14240 39896 14246 39908
rect 15010 39896 15016 39908
rect 14240 39868 15016 39896
rect 14240 39856 14246 39868
rect 15010 39856 15016 39868
rect 15068 39856 15074 39908
rect 17681 39899 17739 39905
rect 17681 39865 17693 39899
rect 17727 39896 17739 39899
rect 18322 39896 18328 39908
rect 17727 39868 18328 39896
rect 17727 39865 17739 39868
rect 17681 39859 17739 39865
rect 18322 39856 18328 39868
rect 18380 39856 18386 39908
rect 20533 39899 20591 39905
rect 20533 39865 20545 39899
rect 20579 39896 20591 39899
rect 21008 39896 21036 39995
rect 21174 39992 21180 40004
rect 21232 39992 21238 40044
rect 22002 40041 22008 40044
rect 21978 40035 22008 40041
rect 21978 40001 21990 40035
rect 21978 39995 22008 40001
rect 22002 39992 22008 39995
rect 22060 39992 22066 40044
rect 23014 40032 23020 40044
rect 22975 40004 23020 40032
rect 23014 39992 23020 40004
rect 23072 39992 23078 40044
rect 23293 40035 23351 40041
rect 23293 40001 23305 40035
rect 23339 40032 23351 40035
rect 23566 40032 23572 40044
rect 23339 40004 23572 40032
rect 23339 40001 23351 40004
rect 23293 39995 23351 40001
rect 23566 39992 23572 40004
rect 23624 39992 23630 40044
rect 24136 40041 24164 40072
rect 25590 40060 25596 40072
rect 25648 40060 25654 40112
rect 25774 40060 25780 40112
rect 25832 40060 25838 40112
rect 25958 40100 25964 40112
rect 25884 40072 25964 40100
rect 24121 40035 24179 40041
rect 24121 40001 24133 40035
rect 24167 40001 24179 40035
rect 24121 39995 24179 40001
rect 25498 39992 25504 40044
rect 25556 40032 25562 40044
rect 25792 40032 25820 40060
rect 25884 40041 25912 40072
rect 25958 40060 25964 40072
rect 26016 40060 26022 40112
rect 26234 40060 26240 40112
rect 26292 40100 26298 40112
rect 26292 40072 27016 40100
rect 26292 40060 26298 40072
rect 26988 40041 27016 40072
rect 27264 40072 27844 40100
rect 25556 40004 25820 40032
rect 25869 40035 25927 40041
rect 25556 39992 25562 40004
rect 25869 40001 25881 40035
rect 25915 40001 25927 40035
rect 25869 39995 25927 40001
rect 26973 40035 27031 40041
rect 26973 40001 26985 40035
rect 27019 40001 27031 40035
rect 26973 39995 27031 40001
rect 27062 39992 27068 40044
rect 27120 40032 27126 40044
rect 27264 40041 27292 40072
rect 27249 40035 27307 40041
rect 27120 40004 27165 40032
rect 27120 39992 27126 40004
rect 27249 40001 27261 40035
rect 27295 40001 27307 40035
rect 27249 39995 27307 40001
rect 22097 39967 22155 39973
rect 22097 39933 22109 39967
rect 22143 39964 22155 39967
rect 22186 39964 22192 39976
rect 22143 39936 22192 39964
rect 22143 39933 22155 39936
rect 22097 39927 22155 39933
rect 22186 39924 22192 39936
rect 22244 39924 22250 39976
rect 24026 39964 24032 39976
rect 23987 39936 24032 39964
rect 24026 39924 24032 39936
rect 24084 39924 24090 39976
rect 25777 39967 25835 39973
rect 25777 39964 25789 39967
rect 25148 39936 25789 39964
rect 20579 39868 21036 39896
rect 22373 39899 22431 39905
rect 20579 39865 20591 39868
rect 20533 39859 20591 39865
rect 22373 39865 22385 39899
rect 22419 39896 22431 39899
rect 25038 39896 25044 39908
rect 22419 39868 25044 39896
rect 22419 39865 22431 39868
rect 22373 39859 22431 39865
rect 25038 39856 25044 39868
rect 25096 39856 25102 39908
rect 15654 39788 15660 39840
rect 15712 39828 15718 39840
rect 16117 39831 16175 39837
rect 16117 39828 16129 39831
rect 15712 39800 16129 39828
rect 15712 39788 15718 39800
rect 16117 39797 16129 39800
rect 16163 39828 16175 39831
rect 16298 39828 16304 39840
rect 16163 39800 16304 39828
rect 16163 39797 16175 39800
rect 16117 39791 16175 39797
rect 16298 39788 16304 39800
rect 16356 39788 16362 39840
rect 17218 39788 17224 39840
rect 17276 39828 17282 39840
rect 18046 39828 18052 39840
rect 17276 39800 18052 39828
rect 17276 39788 17282 39800
rect 18046 39788 18052 39800
rect 18104 39788 18110 39840
rect 18414 39828 18420 39840
rect 18375 39800 18420 39828
rect 18414 39788 18420 39800
rect 18472 39788 18478 39840
rect 19426 39788 19432 39840
rect 19484 39828 19490 39840
rect 20438 39828 20444 39840
rect 19484 39800 20444 39828
rect 19484 39788 19490 39800
rect 20438 39788 20444 39800
rect 20496 39828 20502 39840
rect 20806 39828 20812 39840
rect 20496 39800 20812 39828
rect 20496 39788 20502 39800
rect 20806 39788 20812 39800
rect 20864 39788 20870 39840
rect 21177 39831 21235 39837
rect 21177 39797 21189 39831
rect 21223 39828 21235 39831
rect 21818 39828 21824 39840
rect 21223 39800 21824 39828
rect 21223 39797 21235 39800
rect 21177 39791 21235 39797
rect 21818 39788 21824 39800
rect 21876 39788 21882 39840
rect 22278 39788 22284 39840
rect 22336 39828 22342 39840
rect 24670 39828 24676 39840
rect 22336 39800 24676 39828
rect 22336 39788 22342 39800
rect 24670 39788 24676 39800
rect 24728 39828 24734 39840
rect 24949 39831 25007 39837
rect 24949 39828 24961 39831
rect 24728 39800 24961 39828
rect 24728 39788 24734 39800
rect 24949 39797 24961 39800
rect 24995 39828 25007 39831
rect 25148 39828 25176 39936
rect 25777 39933 25789 39936
rect 25823 39964 25835 39967
rect 26694 39964 26700 39976
rect 25823 39936 26700 39964
rect 25823 39933 25835 39936
rect 25777 39927 25835 39933
rect 26694 39924 26700 39936
rect 26752 39924 26758 39976
rect 27154 39924 27160 39976
rect 27212 39964 27218 39976
rect 27264 39964 27292 39995
rect 27522 39992 27528 40044
rect 27580 40032 27586 40044
rect 27709 40035 27767 40041
rect 27709 40032 27721 40035
rect 27580 40004 27721 40032
rect 27580 39992 27586 40004
rect 27709 40001 27721 40004
rect 27755 40001 27767 40035
rect 27816 40032 27844 40072
rect 29932 40072 30420 40100
rect 27893 40035 27951 40041
rect 27893 40032 27905 40035
rect 27816 40004 27905 40032
rect 27709 39995 27767 40001
rect 27893 40001 27905 40004
rect 27939 40032 27951 40035
rect 29181 40035 29239 40041
rect 29181 40032 29193 40035
rect 27939 40004 29193 40032
rect 27939 40001 27951 40004
rect 27893 39995 27951 40001
rect 29181 40001 29193 40004
rect 29227 40001 29239 40035
rect 29181 39995 29239 40001
rect 29365 40035 29423 40041
rect 29365 40001 29377 40035
rect 29411 40032 29423 40035
rect 29932 40032 29960 40072
rect 30392 40044 30420 40072
rect 32122 40060 32128 40112
rect 32180 40100 32186 40112
rect 32585 40103 32643 40109
rect 32585 40100 32597 40103
rect 32180 40072 32597 40100
rect 32180 40060 32186 40072
rect 32585 40069 32597 40072
rect 32631 40100 32643 40103
rect 33962 40100 33968 40112
rect 32631 40072 33968 40100
rect 32631 40069 32643 40072
rect 32585 40063 32643 40069
rect 33962 40060 33968 40072
rect 34020 40060 34026 40112
rect 35434 40100 35440 40112
rect 34256 40072 34744 40100
rect 30098 40032 30104 40044
rect 29411 40004 29960 40032
rect 30059 40004 30104 40032
rect 29411 40001 29423 40004
rect 29365 39995 29423 40001
rect 30098 39992 30104 40004
rect 30156 39992 30162 40044
rect 30282 40032 30288 40044
rect 30243 40004 30288 40032
rect 30282 39992 30288 40004
rect 30340 39992 30346 40044
rect 30374 39992 30380 40044
rect 30432 39992 30438 40044
rect 30466 39992 30472 40044
rect 30524 40032 30530 40044
rect 30837 40035 30895 40041
rect 30837 40032 30849 40035
rect 30524 40004 30849 40032
rect 30524 39992 30530 40004
rect 30837 40001 30849 40004
rect 30883 40032 30895 40035
rect 32306 40032 32312 40044
rect 30883 40004 32312 40032
rect 30883 40001 30895 40004
rect 30837 39995 30895 40001
rect 32306 39992 32312 40004
rect 32364 39992 32370 40044
rect 33226 39992 33232 40044
rect 33284 40032 33290 40044
rect 33413 40035 33471 40041
rect 33413 40032 33425 40035
rect 33284 40004 33425 40032
rect 33284 39992 33290 40004
rect 33413 40001 33425 40004
rect 33459 40001 33471 40035
rect 33594 40032 33600 40044
rect 33555 40004 33600 40032
rect 33413 39995 33471 40001
rect 33594 39992 33600 40004
rect 33652 39992 33658 40044
rect 33778 39992 33784 40044
rect 33836 40032 33842 40044
rect 34256 40041 34284 40072
rect 34241 40035 34299 40041
rect 34241 40032 34253 40035
rect 33836 40004 34253 40032
rect 33836 39992 33842 40004
rect 34241 40001 34253 40004
rect 34287 40001 34299 40035
rect 34241 39995 34299 40001
rect 34330 39992 34336 40044
rect 34388 40032 34394 40044
rect 34609 40035 34667 40041
rect 34609 40032 34621 40035
rect 34388 40004 34621 40032
rect 34388 39992 34394 40004
rect 34609 40001 34621 40004
rect 34655 40001 34667 40035
rect 34609 39995 34667 40001
rect 27212 39936 27292 39964
rect 27801 39967 27859 39973
rect 27212 39924 27218 39936
rect 27801 39933 27813 39967
rect 27847 39964 27859 39967
rect 30190 39964 30196 39976
rect 27847 39936 30196 39964
rect 27847 39933 27859 39936
rect 27801 39927 27859 39933
rect 30190 39924 30196 39936
rect 30248 39924 30254 39976
rect 32030 39924 32036 39976
rect 32088 39964 32094 39976
rect 34057 39967 34115 39973
rect 34057 39964 34069 39967
rect 32088 39936 34069 39964
rect 32088 39924 32094 39936
rect 34057 39933 34069 39936
rect 34103 39933 34115 39967
rect 34057 39927 34115 39933
rect 34425 39967 34483 39973
rect 34425 39933 34437 39967
rect 34471 39933 34483 39967
rect 34425 39927 34483 39933
rect 26050 39856 26056 39908
rect 26108 39896 26114 39908
rect 29362 39896 29368 39908
rect 26108 39868 28994 39896
rect 29323 39868 29368 39896
rect 26108 39856 26114 39868
rect 25866 39828 25872 39840
rect 24995 39800 25176 39828
rect 25827 39800 25872 39828
rect 24995 39797 25007 39800
rect 24949 39791 25007 39797
rect 25866 39788 25872 39800
rect 25924 39788 25930 39840
rect 26421 39831 26479 39837
rect 26421 39797 26433 39831
rect 26467 39828 26479 39831
rect 26694 39828 26700 39840
rect 26467 39800 26700 39828
rect 26467 39797 26479 39800
rect 26421 39791 26479 39797
rect 26694 39788 26700 39800
rect 26752 39788 26758 39840
rect 28350 39828 28356 39840
rect 28311 39800 28356 39828
rect 28350 39788 28356 39800
rect 28408 39788 28414 39840
rect 28966 39828 28994 39868
rect 29362 39856 29368 39868
rect 29420 39856 29426 39908
rect 30466 39896 30472 39908
rect 29472 39868 30472 39896
rect 29472 39828 29500 39868
rect 30466 39856 30472 39868
rect 30524 39856 30530 39908
rect 33410 39896 33416 39908
rect 33371 39868 33416 39896
rect 33410 39856 33416 39868
rect 33468 39856 33474 39908
rect 34440 39896 34468 39927
rect 34514 39924 34520 39976
rect 34572 39964 34578 39976
rect 34716 39964 34744 40072
rect 34808 40072 35440 40100
rect 34808 40041 34836 40072
rect 35434 40060 35440 40072
rect 35492 40060 35498 40112
rect 36004 40100 36032 40128
rect 35728 40072 36032 40100
rect 36372 40072 36676 40100
rect 35728 40041 35756 40072
rect 36372 40044 36400 40072
rect 34793 40035 34851 40041
rect 34793 40001 34805 40035
rect 34839 40001 34851 40035
rect 34793 39995 34851 40001
rect 35713 40035 35771 40041
rect 35713 40001 35725 40035
rect 35759 40001 35771 40035
rect 35713 39995 35771 40001
rect 35894 39992 35900 40044
rect 35952 40032 35958 40044
rect 35989 40035 36047 40041
rect 35989 40032 36001 40035
rect 35952 40004 36001 40032
rect 35952 39992 35958 40004
rect 35989 40001 36001 40004
rect 36035 40001 36047 40035
rect 35989 39995 36047 40001
rect 35434 39964 35440 39976
rect 34572 39936 34617 39964
rect 34716 39936 35440 39964
rect 34572 39924 34578 39936
rect 35434 39924 35440 39936
rect 35492 39924 35498 39976
rect 35802 39964 35808 39976
rect 35763 39936 35808 39964
rect 35802 39924 35808 39936
rect 35860 39924 35866 39976
rect 36004 39964 36032 39995
rect 36354 39992 36360 40044
rect 36412 39992 36418 40044
rect 36538 40032 36544 40044
rect 36499 40004 36544 40032
rect 36538 39992 36544 40004
rect 36596 39992 36602 40044
rect 36648 40032 36676 40072
rect 36725 40035 36783 40041
rect 36725 40032 36737 40035
rect 36648 40004 36737 40032
rect 36725 40001 36737 40004
rect 36771 40001 36783 40035
rect 37458 40032 37464 40044
rect 37419 40004 37464 40032
rect 36725 39995 36783 40001
rect 37458 39992 37464 40004
rect 37516 39992 37522 40044
rect 37752 40041 37780 40140
rect 38742 40137 38754 40140
rect 38788 40137 38800 40171
rect 41598 40168 41604 40180
rect 41559 40140 41604 40168
rect 38742 40131 38800 40137
rect 41598 40128 41604 40140
rect 41656 40128 41662 40180
rect 38657 40103 38715 40109
rect 38657 40069 38669 40103
rect 38703 40100 38715 40103
rect 38703 40072 39528 40100
rect 38703 40069 38715 40072
rect 38657 40063 38715 40069
rect 39500 40044 39528 40072
rect 37737 40035 37795 40041
rect 37737 40001 37749 40035
rect 37783 40001 37795 40035
rect 37737 39995 37795 40001
rect 38565 40035 38623 40041
rect 38565 40001 38577 40035
rect 38611 40001 38623 40035
rect 38838 40032 38844 40044
rect 38799 40004 38844 40032
rect 38565 39995 38623 40001
rect 36630 39964 36636 39976
rect 36004 39936 36636 39964
rect 36630 39924 36636 39936
rect 36688 39924 36694 39976
rect 37277 39967 37335 39973
rect 37277 39933 37289 39967
rect 37323 39964 37335 39967
rect 37366 39964 37372 39976
rect 37323 39936 37372 39964
rect 37323 39933 37335 39936
rect 37277 39927 37335 39933
rect 37366 39924 37372 39936
rect 37424 39924 37430 39976
rect 37553 39967 37611 39973
rect 37553 39933 37565 39967
rect 37599 39964 37611 39967
rect 37918 39964 37924 39976
rect 37599 39936 37924 39964
rect 37599 39933 37611 39936
rect 37553 39927 37611 39933
rect 37918 39924 37924 39936
rect 37976 39924 37982 39976
rect 38010 39924 38016 39976
rect 38068 39964 38074 39976
rect 38580 39964 38608 39995
rect 38838 39992 38844 40004
rect 38896 39992 38902 40044
rect 39301 40035 39359 40041
rect 39301 40001 39313 40035
rect 39347 40001 39359 40035
rect 39482 40032 39488 40044
rect 39443 40004 39488 40032
rect 39301 39995 39359 40001
rect 39316 39964 39344 39995
rect 39482 39992 39488 40004
rect 39540 39992 39546 40044
rect 40494 40032 40500 40044
rect 40455 40004 40500 40032
rect 40494 39992 40500 40004
rect 40552 40032 40558 40044
rect 41690 40032 41696 40044
rect 40552 40004 41696 40032
rect 40552 39992 40558 40004
rect 41690 39992 41696 40004
rect 41748 39992 41754 40044
rect 40218 39964 40224 39976
rect 38068 39936 40224 39964
rect 38068 39924 38074 39936
rect 40218 39924 40224 39936
rect 40276 39924 40282 39976
rect 35897 39899 35955 39905
rect 34440 39868 35848 39896
rect 30190 39828 30196 39840
rect 28966 39800 29500 39828
rect 30151 39800 30196 39828
rect 30190 39788 30196 39800
rect 30248 39788 30254 39840
rect 31110 39788 31116 39840
rect 31168 39828 31174 39840
rect 31297 39831 31355 39837
rect 31297 39828 31309 39831
rect 31168 39800 31309 39828
rect 31168 39788 31174 39800
rect 31297 39797 31309 39800
rect 31343 39797 31355 39831
rect 32858 39828 32864 39840
rect 32819 39800 32864 39828
rect 31297 39791 31355 39797
rect 32858 39788 32864 39800
rect 32916 39788 32922 39840
rect 34514 39788 34520 39840
rect 34572 39828 34578 39840
rect 35710 39828 35716 39840
rect 34572 39800 35716 39828
rect 34572 39788 34578 39800
rect 35710 39788 35716 39800
rect 35768 39788 35774 39840
rect 35820 39828 35848 39868
rect 35897 39865 35909 39899
rect 35943 39896 35955 39899
rect 36078 39896 36084 39908
rect 35943 39868 36084 39896
rect 35943 39865 35955 39868
rect 35897 39859 35955 39865
rect 36078 39856 36084 39868
rect 36136 39896 36142 39908
rect 37645 39899 37703 39905
rect 37645 39896 37657 39899
rect 36136 39868 37657 39896
rect 36136 39856 36142 39868
rect 37645 39865 37657 39868
rect 37691 39896 37703 39899
rect 39114 39896 39120 39908
rect 37691 39868 39120 39896
rect 37691 39865 37703 39868
rect 37645 39859 37703 39865
rect 39114 39856 39120 39868
rect 39172 39856 39178 39908
rect 40034 39896 40040 39908
rect 39947 39868 40040 39896
rect 40034 39856 40040 39868
rect 40092 39896 40098 39908
rect 41322 39896 41328 39908
rect 40092 39868 41328 39896
rect 40092 39856 40098 39868
rect 41322 39856 41328 39868
rect 41380 39856 41386 39908
rect 37458 39828 37464 39840
rect 35820 39800 37464 39828
rect 37458 39788 37464 39800
rect 37516 39788 37522 39840
rect 39393 39831 39451 39837
rect 39393 39797 39405 39831
rect 39439 39828 39451 39831
rect 39850 39828 39856 39840
rect 39439 39800 39856 39828
rect 39439 39797 39451 39800
rect 39393 39791 39451 39797
rect 39850 39788 39856 39800
rect 39908 39788 39914 39840
rect 40954 39788 40960 39840
rect 41012 39828 41018 39840
rect 41049 39831 41107 39837
rect 41049 39828 41061 39831
rect 41012 39800 41061 39828
rect 41012 39788 41018 39800
rect 41049 39797 41061 39800
rect 41095 39797 41107 39831
rect 41049 39791 41107 39797
rect 42058 39788 42064 39840
rect 42116 39828 42122 39840
rect 42429 39831 42487 39837
rect 42429 39828 42441 39831
rect 42116 39800 42441 39828
rect 42116 39788 42122 39800
rect 42429 39797 42441 39800
rect 42475 39797 42487 39831
rect 42429 39791 42487 39797
rect 43073 39831 43131 39837
rect 43073 39797 43085 39831
rect 43119 39828 43131 39831
rect 43162 39828 43168 39840
rect 43119 39800 43168 39828
rect 43119 39797 43131 39800
rect 43073 39791 43131 39797
rect 43162 39788 43168 39800
rect 43220 39788 43226 39840
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 11146 39624 11152 39636
rect 11107 39596 11152 39624
rect 11146 39584 11152 39596
rect 11204 39584 11210 39636
rect 12802 39624 12808 39636
rect 12763 39596 12808 39624
rect 12802 39584 12808 39596
rect 12860 39624 12866 39636
rect 16942 39624 16948 39636
rect 12860 39596 16948 39624
rect 12860 39584 12866 39596
rect 16942 39584 16948 39596
rect 17000 39584 17006 39636
rect 17034 39584 17040 39636
rect 17092 39624 17098 39636
rect 20901 39627 20959 39633
rect 17092 39596 18460 39624
rect 17092 39584 17098 39596
rect 15565 39559 15623 39565
rect 14384 39528 15240 39556
rect 13814 39488 13820 39500
rect 13372 39460 13820 39488
rect 13372 39429 13400 39460
rect 13814 39448 13820 39460
rect 13872 39448 13878 39500
rect 13357 39423 13415 39429
rect 13357 39389 13369 39423
rect 13403 39389 13415 39423
rect 13357 39383 13415 39389
rect 13541 39423 13599 39429
rect 13541 39389 13553 39423
rect 13587 39420 13599 39423
rect 14093 39423 14151 39429
rect 14093 39420 14105 39423
rect 13587 39392 14105 39420
rect 13587 39389 13599 39392
rect 13541 39383 13599 39389
rect 14093 39389 14105 39392
rect 14139 39389 14151 39423
rect 14093 39383 14151 39389
rect 14384 39364 14412 39528
rect 14458 39448 14464 39500
rect 14516 39488 14522 39500
rect 15105 39491 15163 39497
rect 15105 39488 15117 39491
rect 14516 39460 15117 39488
rect 14516 39448 14522 39460
rect 15105 39457 15117 39460
rect 15151 39457 15163 39491
rect 15212 39488 15240 39528
rect 15565 39525 15577 39559
rect 15611 39556 15623 39559
rect 17865 39559 17923 39565
rect 17865 39556 17877 39559
rect 15611 39528 17877 39556
rect 15611 39525 15623 39528
rect 15565 39519 15623 39525
rect 17865 39525 17877 39528
rect 17911 39525 17923 39559
rect 18432 39556 18460 39596
rect 20901 39593 20913 39627
rect 20947 39624 20959 39627
rect 21174 39624 21180 39636
rect 20947 39596 21180 39624
rect 20947 39593 20959 39596
rect 20901 39587 20959 39593
rect 21174 39584 21180 39596
rect 21232 39584 21238 39636
rect 22281 39627 22339 39633
rect 22281 39593 22293 39627
rect 22327 39624 22339 39627
rect 22370 39624 22376 39636
rect 22327 39596 22376 39624
rect 22327 39593 22339 39596
rect 22281 39587 22339 39593
rect 22370 39584 22376 39596
rect 22428 39584 22434 39636
rect 23845 39627 23903 39633
rect 23845 39593 23857 39627
rect 23891 39624 23903 39627
rect 24486 39624 24492 39636
rect 23891 39596 24492 39624
rect 23891 39593 23903 39596
rect 23845 39587 23903 39593
rect 24486 39584 24492 39596
rect 24544 39584 24550 39636
rect 26697 39627 26755 39633
rect 26697 39593 26709 39627
rect 26743 39624 26755 39627
rect 27062 39624 27068 39636
rect 26743 39596 27068 39624
rect 26743 39593 26755 39596
rect 26697 39587 26755 39593
rect 27062 39584 27068 39596
rect 27120 39584 27126 39636
rect 28629 39627 28687 39633
rect 28629 39593 28641 39627
rect 28675 39624 28687 39627
rect 28810 39624 28816 39636
rect 28675 39596 28816 39624
rect 28675 39593 28687 39596
rect 28629 39587 28687 39593
rect 28810 39584 28816 39596
rect 28868 39584 28874 39636
rect 29822 39624 29828 39636
rect 28920 39596 29828 39624
rect 18432 39528 23520 39556
rect 17865 39519 17923 39525
rect 17954 39488 17960 39500
rect 15212 39460 17960 39488
rect 15105 39451 15163 39457
rect 17954 39448 17960 39460
rect 18012 39448 18018 39500
rect 18322 39488 18328 39500
rect 18064 39460 18328 39488
rect 18064 39432 18092 39460
rect 18322 39448 18328 39460
rect 18380 39448 18386 39500
rect 20346 39448 20352 39500
rect 20404 39488 20410 39500
rect 20533 39491 20591 39497
rect 20533 39488 20545 39491
rect 20404 39460 20545 39488
rect 20404 39448 20410 39460
rect 20533 39457 20545 39460
rect 20579 39457 20591 39491
rect 21818 39488 21824 39500
rect 21779 39460 21824 39488
rect 20533 39451 20591 39457
rect 21818 39448 21824 39460
rect 21876 39448 21882 39500
rect 21913 39491 21971 39497
rect 21913 39457 21925 39491
rect 21959 39488 21971 39491
rect 22646 39488 22652 39500
rect 21959 39460 22652 39488
rect 21959 39457 21971 39460
rect 21913 39451 21971 39457
rect 22646 39448 22652 39460
rect 22704 39448 22710 39500
rect 23382 39448 23388 39500
rect 23440 39448 23446 39500
rect 15197 39423 15255 39429
rect 15197 39420 15209 39423
rect 14568 39392 15209 39420
rect 10870 39312 10876 39364
rect 10928 39352 10934 39364
rect 11701 39355 11759 39361
rect 11701 39352 11713 39355
rect 10928 39324 11713 39352
rect 10928 39312 10934 39324
rect 11701 39321 11713 39324
rect 11747 39321 11759 39355
rect 11701 39315 11759 39321
rect 13630 39312 13636 39364
rect 13688 39352 13694 39364
rect 14277 39355 14335 39361
rect 14277 39352 14289 39355
rect 13688 39324 14289 39352
rect 13688 39312 13694 39324
rect 14277 39321 14289 39324
rect 14323 39321 14335 39355
rect 14277 39315 14335 39321
rect 14366 39312 14372 39364
rect 14424 39352 14430 39364
rect 14461 39355 14519 39361
rect 14461 39352 14473 39355
rect 14424 39324 14473 39352
rect 14424 39312 14430 39324
rect 14461 39321 14473 39324
rect 14507 39321 14519 39355
rect 14461 39315 14519 39321
rect 14568 39296 14596 39392
rect 15197 39389 15209 39392
rect 15243 39420 15255 39423
rect 15746 39420 15752 39432
rect 15243 39392 15752 39420
rect 15243 39389 15255 39392
rect 15197 39383 15255 39389
rect 15746 39380 15752 39392
rect 15804 39380 15810 39432
rect 16114 39380 16120 39432
rect 16172 39420 16178 39432
rect 16209 39423 16267 39429
rect 16209 39420 16221 39423
rect 16172 39392 16221 39420
rect 16172 39380 16178 39392
rect 16209 39389 16221 39392
rect 16255 39389 16267 39423
rect 16390 39420 16396 39432
rect 16351 39392 16396 39420
rect 16209 39383 16267 39389
rect 16390 39380 16396 39392
rect 16448 39380 16454 39432
rect 16942 39380 16948 39432
rect 17000 39420 17006 39432
rect 17770 39420 17776 39432
rect 17000 39392 17776 39420
rect 17000 39380 17006 39392
rect 17770 39380 17776 39392
rect 17828 39380 17834 39432
rect 18046 39420 18052 39432
rect 18007 39392 18052 39420
rect 18046 39380 18052 39392
rect 18104 39380 18110 39432
rect 18141 39423 18199 39429
rect 18141 39389 18153 39423
rect 18187 39389 18199 39423
rect 18141 39383 18199 39389
rect 17310 39312 17316 39364
rect 17368 39352 17374 39364
rect 18156 39352 18184 39383
rect 18874 39380 18880 39432
rect 18932 39420 18938 39432
rect 20441 39423 20499 39429
rect 20441 39420 20453 39423
rect 18932 39392 20453 39420
rect 18932 39380 18938 39392
rect 20441 39389 20453 39392
rect 20487 39389 20499 39423
rect 20622 39420 20628 39432
rect 20583 39392 20628 39420
rect 20441 39383 20499 39389
rect 20622 39380 20628 39392
rect 20680 39380 20686 39432
rect 20717 39423 20775 39429
rect 20717 39389 20729 39423
rect 20763 39389 20775 39423
rect 20717 39383 20775 39389
rect 17368 39324 18184 39352
rect 18325 39355 18383 39361
rect 17368 39312 17374 39324
rect 18325 39321 18337 39355
rect 18371 39352 18383 39355
rect 18371 39324 20208 39352
rect 18371 39321 18383 39324
rect 18325 39315 18383 39321
rect 12250 39284 12256 39296
rect 12211 39256 12256 39284
rect 12250 39244 12256 39256
rect 12308 39244 12314 39296
rect 13449 39287 13507 39293
rect 13449 39253 13461 39287
rect 13495 39284 13507 39287
rect 14550 39284 14556 39296
rect 13495 39256 14556 39284
rect 13495 39253 13507 39256
rect 13449 39247 13507 39253
rect 14550 39244 14556 39256
rect 14608 39244 14614 39296
rect 16206 39284 16212 39296
rect 16167 39256 16212 39284
rect 16206 39244 16212 39256
rect 16264 39244 16270 39296
rect 17221 39287 17279 39293
rect 17221 39253 17233 39287
rect 17267 39284 17279 39287
rect 19334 39284 19340 39296
rect 17267 39256 19340 39284
rect 17267 39253 17279 39256
rect 17221 39247 17279 39253
rect 19334 39244 19340 39256
rect 19392 39244 19398 39296
rect 19426 39244 19432 39296
rect 19484 39284 19490 39296
rect 19797 39287 19855 39293
rect 19797 39284 19809 39287
rect 19484 39256 19809 39284
rect 19484 39244 19490 39256
rect 19797 39253 19809 39256
rect 19843 39253 19855 39287
rect 20180 39284 20208 39324
rect 20530 39312 20536 39364
rect 20588 39352 20594 39364
rect 20732 39352 20760 39383
rect 22094 39380 22100 39432
rect 22152 39420 22158 39432
rect 22925 39423 22983 39429
rect 22925 39420 22937 39423
rect 22152 39392 22937 39420
rect 22152 39380 22158 39392
rect 22925 39389 22937 39392
rect 22971 39420 22983 39423
rect 23400 39420 23428 39448
rect 23492 39429 23520 39528
rect 23934 39516 23940 39568
rect 23992 39556 23998 39568
rect 24854 39556 24860 39568
rect 23992 39528 24860 39556
rect 23992 39516 23998 39528
rect 24854 39516 24860 39528
rect 24912 39516 24918 39568
rect 25498 39516 25504 39568
rect 25556 39556 25562 39568
rect 27249 39559 27307 39565
rect 27249 39556 27261 39559
rect 25556 39528 27261 39556
rect 25556 39516 25562 39528
rect 27249 39525 27261 39528
rect 27295 39525 27307 39559
rect 27249 39519 27307 39525
rect 27985 39559 28043 39565
rect 27985 39525 27997 39559
rect 28031 39556 28043 39559
rect 28920 39556 28948 39596
rect 29822 39584 29828 39596
rect 29880 39584 29886 39636
rect 33321 39627 33379 39633
rect 33321 39593 33333 39627
rect 33367 39624 33379 39627
rect 34330 39624 34336 39636
rect 33367 39596 34336 39624
rect 33367 39593 33379 39596
rect 33321 39587 33379 39593
rect 34330 39584 34336 39596
rect 34388 39584 34394 39636
rect 35894 39624 35900 39636
rect 34624 39596 35900 39624
rect 31386 39556 31392 39568
rect 28031 39528 28948 39556
rect 29656 39528 31392 39556
rect 28031 39525 28043 39528
rect 27985 39519 28043 39525
rect 24578 39448 24584 39500
rect 24636 39488 24642 39500
rect 25777 39491 25835 39497
rect 25777 39488 25789 39491
rect 24636 39460 25789 39488
rect 24636 39448 24642 39460
rect 25777 39457 25789 39460
rect 25823 39488 25835 39491
rect 26050 39488 26056 39500
rect 25823 39460 26056 39488
rect 25823 39457 25835 39460
rect 25777 39451 25835 39457
rect 26050 39448 26056 39460
rect 26108 39448 26114 39500
rect 26142 39448 26148 39500
rect 26200 39488 26206 39500
rect 27154 39488 27160 39500
rect 26200 39460 27160 39488
rect 26200 39448 26206 39460
rect 27154 39448 27160 39460
rect 27212 39488 27218 39500
rect 29656 39497 29684 39528
rect 31386 39516 31392 39528
rect 31444 39516 31450 39568
rect 31754 39516 31760 39568
rect 31812 39556 31818 39568
rect 33781 39559 33839 39565
rect 33781 39556 33793 39559
rect 31812 39528 33793 39556
rect 31812 39516 31818 39528
rect 33781 39525 33793 39528
rect 33827 39525 33839 39559
rect 33781 39519 33839 39525
rect 33962 39516 33968 39568
rect 34020 39556 34026 39568
rect 34624 39556 34652 39596
rect 35894 39584 35900 39596
rect 35952 39584 35958 39636
rect 35986 39584 35992 39636
rect 36044 39624 36050 39636
rect 36265 39627 36323 39633
rect 36265 39624 36277 39627
rect 36044 39596 36277 39624
rect 36044 39584 36050 39596
rect 36265 39593 36277 39596
rect 36311 39593 36323 39627
rect 36265 39587 36323 39593
rect 36354 39584 36360 39636
rect 36412 39624 36418 39636
rect 38654 39624 38660 39636
rect 36412 39596 38660 39624
rect 36412 39584 36418 39596
rect 38654 39584 38660 39596
rect 38712 39584 38718 39636
rect 38749 39627 38807 39633
rect 38749 39593 38761 39627
rect 38795 39624 38807 39627
rect 38838 39624 38844 39636
rect 38795 39596 38844 39624
rect 38795 39593 38807 39596
rect 38749 39587 38807 39593
rect 38838 39584 38844 39596
rect 38896 39584 38902 39636
rect 38933 39627 38991 39633
rect 38933 39593 38945 39627
rect 38979 39624 38991 39627
rect 39022 39624 39028 39636
rect 38979 39596 39028 39624
rect 38979 39593 38991 39596
rect 38933 39587 38991 39593
rect 39022 39584 39028 39596
rect 39080 39584 39086 39636
rect 39114 39584 39120 39636
rect 39172 39624 39178 39636
rect 39945 39627 40003 39633
rect 39945 39624 39957 39627
rect 39172 39596 39957 39624
rect 39172 39584 39178 39596
rect 39945 39593 39957 39596
rect 39991 39593 40003 39627
rect 39945 39587 40003 39593
rect 34020 39528 34652 39556
rect 34020 39516 34026 39528
rect 29641 39491 29699 39497
rect 27212 39460 28856 39488
rect 27212 39448 27218 39460
rect 22971 39392 23428 39420
rect 23477 39423 23535 39429
rect 22971 39389 22983 39392
rect 22925 39383 22983 39389
rect 23477 39389 23489 39423
rect 23523 39389 23535 39423
rect 23477 39383 23535 39389
rect 24210 39380 24216 39432
rect 24268 39420 24274 39432
rect 24765 39423 24823 39429
rect 24765 39420 24777 39423
rect 24268 39392 24777 39420
rect 24268 39380 24274 39392
rect 24765 39389 24777 39392
rect 24811 39389 24823 39423
rect 25498 39420 25504 39432
rect 25459 39392 25504 39420
rect 24765 39383 24823 39389
rect 25498 39380 25504 39392
rect 25556 39380 25562 39432
rect 25590 39380 25596 39432
rect 25648 39420 25654 39432
rect 26237 39423 26295 39429
rect 26237 39420 26249 39423
rect 25648 39392 26249 39420
rect 25648 39380 25654 39392
rect 26237 39389 26249 39392
rect 26283 39420 26295 39423
rect 26418 39420 26424 39432
rect 26283 39392 26424 39420
rect 26283 39389 26295 39392
rect 26237 39383 26295 39389
rect 26418 39380 26424 39392
rect 26476 39380 26482 39432
rect 26513 39423 26571 39429
rect 26513 39389 26525 39423
rect 26559 39389 26571 39423
rect 26513 39383 26571 39389
rect 20588 39324 20760 39352
rect 20588 39312 20594 39324
rect 20806 39312 20812 39364
rect 20864 39352 20870 39364
rect 23661 39355 23719 39361
rect 23661 39352 23673 39355
rect 20864 39324 23673 39352
rect 20864 39312 20870 39324
rect 23661 39321 23673 39324
rect 23707 39352 23719 39355
rect 25222 39352 25228 39364
rect 23707 39324 25228 39352
rect 23707 39321 23719 39324
rect 23661 39315 23719 39321
rect 25222 39312 25228 39324
rect 25280 39312 25286 39364
rect 25777 39355 25835 39361
rect 25777 39321 25789 39355
rect 25823 39352 25835 39355
rect 26528 39352 26556 39383
rect 27338 39380 27344 39432
rect 27396 39420 27402 39432
rect 27433 39423 27491 39429
rect 27433 39420 27445 39423
rect 27396 39392 27445 39420
rect 27396 39380 27402 39392
rect 27433 39389 27445 39392
rect 27479 39389 27491 39423
rect 27433 39383 27491 39389
rect 27985 39423 28043 39429
rect 27985 39389 27997 39423
rect 28031 39420 28043 39423
rect 28074 39420 28080 39432
rect 28031 39392 28080 39420
rect 28031 39389 28043 39392
rect 27985 39383 28043 39389
rect 28074 39380 28080 39392
rect 28132 39380 28138 39432
rect 28184 39429 28212 39460
rect 28169 39423 28227 39429
rect 28169 39389 28181 39423
rect 28215 39389 28227 39423
rect 28169 39383 28227 39389
rect 28350 39380 28356 39432
rect 28408 39420 28414 39432
rect 28828 39429 28856 39460
rect 29641 39457 29653 39491
rect 29687 39457 29699 39491
rect 29641 39451 29699 39457
rect 30101 39491 30159 39497
rect 30101 39457 30113 39491
rect 30147 39488 30159 39491
rect 31938 39488 31944 39500
rect 30147 39460 31944 39488
rect 30147 39457 30159 39460
rect 30101 39451 30159 39457
rect 31938 39448 31944 39460
rect 31996 39448 32002 39500
rect 32674 39448 32680 39500
rect 32732 39488 32738 39500
rect 32861 39491 32919 39497
rect 32861 39488 32873 39491
rect 32732 39460 32873 39488
rect 32732 39448 32738 39460
rect 32861 39457 32873 39460
rect 32907 39488 32919 39491
rect 33042 39488 33048 39500
rect 32907 39460 33048 39488
rect 32907 39457 32919 39460
rect 32861 39451 32919 39457
rect 33042 39448 33048 39460
rect 33100 39448 33106 39500
rect 34624 39488 34652 39528
rect 34901 39528 35296 39556
rect 34701 39491 34759 39497
rect 34701 39488 34713 39491
rect 34624 39460 34713 39488
rect 34701 39457 34713 39460
rect 34747 39457 34759 39491
rect 34701 39451 34759 39457
rect 28629 39423 28687 39429
rect 28629 39420 28641 39423
rect 28408 39392 28641 39420
rect 28408 39380 28414 39392
rect 28629 39389 28641 39392
rect 28675 39389 28687 39423
rect 28629 39383 28687 39389
rect 28813 39423 28871 39429
rect 28813 39389 28825 39423
rect 28859 39389 28871 39423
rect 28813 39383 28871 39389
rect 28994 39380 29000 39432
rect 29052 39420 29058 39432
rect 29733 39423 29791 39429
rect 29733 39420 29745 39423
rect 29052 39392 29745 39420
rect 29052 39380 29058 39392
rect 29733 39389 29745 39392
rect 29779 39389 29791 39423
rect 29733 39383 29791 39389
rect 29917 39423 29975 39429
rect 29917 39389 29929 39423
rect 29963 39420 29975 39423
rect 30558 39420 30564 39432
rect 29963 39392 30564 39420
rect 29963 39389 29975 39392
rect 29917 39383 29975 39389
rect 27356 39352 27384 39380
rect 25823 39324 26556 39352
rect 27172 39324 27384 39352
rect 25823 39321 25835 39324
rect 25777 39315 25835 39321
rect 20714 39284 20720 39296
rect 20180 39256 20720 39284
rect 19797 39247 19855 39253
rect 20714 39244 20720 39256
rect 20772 39244 20778 39296
rect 24949 39287 25007 39293
rect 24949 39253 24961 39287
rect 24995 39284 25007 39287
rect 25038 39284 25044 39296
rect 24995 39256 25044 39284
rect 24995 39253 25007 39256
rect 24949 39247 25007 39253
rect 25038 39244 25044 39256
rect 25096 39284 25102 39296
rect 26142 39284 26148 39296
rect 25096 39256 26148 39284
rect 25096 39244 25102 39256
rect 26142 39244 26148 39256
rect 26200 39244 26206 39296
rect 26329 39287 26387 39293
rect 26329 39253 26341 39287
rect 26375 39284 26387 39287
rect 27172 39284 27200 39324
rect 29086 39312 29092 39364
rect 29144 39352 29150 39364
rect 29932 39352 29960 39383
rect 30558 39380 30564 39392
rect 30616 39380 30622 39432
rect 31389 39423 31447 39429
rect 31389 39389 31401 39423
rect 31435 39420 31447 39423
rect 31570 39420 31576 39432
rect 31435 39392 31469 39420
rect 31531 39392 31576 39420
rect 31435 39389 31447 39392
rect 31389 39383 31447 39389
rect 29144 39324 29960 39352
rect 29144 39312 29150 39324
rect 31202 39312 31208 39364
rect 31260 39352 31266 39364
rect 31404 39352 31432 39383
rect 31570 39380 31576 39392
rect 31628 39380 31634 39432
rect 32953 39423 33011 39429
rect 32953 39389 32965 39423
rect 32999 39420 33011 39423
rect 33686 39420 33692 39432
rect 32999 39392 33692 39420
rect 32999 39389 33011 39392
rect 32953 39383 33011 39389
rect 33686 39380 33692 39392
rect 33744 39380 33750 39432
rect 33962 39420 33968 39432
rect 33923 39392 33968 39420
rect 33962 39380 33968 39392
rect 34020 39380 34026 39432
rect 34149 39423 34207 39429
rect 34149 39389 34161 39423
rect 34195 39420 34207 39423
rect 34330 39420 34336 39432
rect 34195 39392 34336 39420
rect 34195 39389 34207 39392
rect 34149 39383 34207 39389
rect 33134 39352 33140 39364
rect 31260 39324 33140 39352
rect 31260 39312 31266 39324
rect 33134 39312 33140 39324
rect 33192 39312 33198 39364
rect 33410 39312 33416 39364
rect 33468 39352 33474 39364
rect 33594 39352 33600 39364
rect 33468 39324 33600 39352
rect 33468 39312 33474 39324
rect 33594 39312 33600 39324
rect 33652 39352 33658 39364
rect 34164 39352 34192 39383
rect 34330 39380 34336 39392
rect 34388 39380 34394 39432
rect 34901 39429 34929 39528
rect 34974 39448 34980 39500
rect 35032 39488 35038 39500
rect 35268 39488 35296 39528
rect 35434 39516 35440 39568
rect 35492 39556 35498 39568
rect 36722 39556 36728 39568
rect 35492 39528 36728 39556
rect 35492 39516 35498 39528
rect 36722 39516 36728 39528
rect 36780 39556 36786 39568
rect 40954 39556 40960 39568
rect 36780 39528 40960 39556
rect 36780 39516 36786 39528
rect 40954 39516 40960 39528
rect 41012 39516 41018 39568
rect 35032 39460 35112 39488
rect 35268 39460 35480 39488
rect 35032 39448 35038 39460
rect 35084 39429 35112 39460
rect 34859 39423 34929 39429
rect 34859 39389 34871 39423
rect 34905 39392 34929 39423
rect 35069 39423 35127 39429
rect 34905 39389 34917 39392
rect 34859 39383 34917 39389
rect 35069 39389 35081 39423
rect 35115 39389 35127 39423
rect 35069 39383 35127 39389
rect 35161 39423 35219 39429
rect 35161 39389 35173 39423
rect 35207 39422 35219 39423
rect 35207 39420 35296 39422
rect 35342 39420 35348 39432
rect 35207 39394 35348 39420
rect 35207 39389 35219 39394
rect 35268 39392 35348 39394
rect 35161 39383 35219 39389
rect 35342 39380 35348 39392
rect 35400 39380 35406 39432
rect 33652 39324 34192 39352
rect 34977 39355 35035 39361
rect 33652 39312 33658 39324
rect 34977 39321 34989 39355
rect 35023 39321 35035 39355
rect 35452 39352 35480 39460
rect 36262 39448 36268 39500
rect 36320 39488 36326 39500
rect 37093 39491 37151 39497
rect 37093 39488 37105 39491
rect 36320 39460 37105 39488
rect 36320 39448 36326 39460
rect 37093 39457 37105 39460
rect 37139 39488 37151 39491
rect 38378 39488 38384 39500
rect 37139 39460 38384 39488
rect 37139 39457 37151 39460
rect 37093 39451 37151 39457
rect 38378 39448 38384 39460
rect 38436 39448 38442 39500
rect 42153 39491 42211 39497
rect 42153 39488 42165 39491
rect 38672 39460 42165 39488
rect 35526 39380 35532 39432
rect 35584 39420 35590 39432
rect 36354 39420 36360 39432
rect 35584 39392 36360 39420
rect 35584 39380 35590 39392
rect 36354 39380 36360 39392
rect 36412 39420 36418 39432
rect 36449 39423 36507 39429
rect 36449 39420 36461 39423
rect 36412 39392 36461 39420
rect 36412 39380 36418 39392
rect 36449 39389 36461 39392
rect 36495 39389 36507 39423
rect 36449 39383 36507 39389
rect 36538 39380 36544 39432
rect 36596 39420 36602 39432
rect 38102 39420 38108 39432
rect 36596 39392 36641 39420
rect 38063 39392 38108 39420
rect 36596 39380 36602 39392
rect 38102 39380 38108 39392
rect 38160 39380 38166 39432
rect 38289 39423 38347 39429
rect 38289 39389 38301 39423
rect 38335 39389 38347 39423
rect 38289 39383 38347 39389
rect 36998 39352 37004 39364
rect 35452 39324 37004 39352
rect 34977 39315 35035 39321
rect 26375 39256 27200 39284
rect 26375 39253 26387 39256
rect 26329 39247 26387 39253
rect 30466 39244 30472 39296
rect 30524 39284 30530 39296
rect 30837 39287 30895 39293
rect 30837 39284 30849 39287
rect 30524 39256 30849 39284
rect 30524 39244 30530 39256
rect 30837 39253 30849 39256
rect 30883 39253 30895 39287
rect 30837 39247 30895 39253
rect 33502 39244 33508 39296
rect 33560 39284 33566 39296
rect 34992 39284 35020 39315
rect 36998 39312 37004 39324
rect 37056 39312 37062 39364
rect 37642 39312 37648 39364
rect 37700 39352 37706 39364
rect 38304 39352 38332 39383
rect 38672 39364 38700 39460
rect 42153 39457 42165 39460
rect 42199 39488 42211 39491
rect 43530 39488 43536 39500
rect 42199 39460 43536 39488
rect 42199 39457 42211 39460
rect 42153 39451 42211 39457
rect 43530 39448 43536 39460
rect 43588 39488 43594 39500
rect 43809 39491 43867 39497
rect 43809 39488 43821 39491
rect 43588 39460 43821 39488
rect 43588 39448 43594 39460
rect 43809 39457 43821 39460
rect 43855 39488 43867 39491
rect 47118 39488 47124 39500
rect 43855 39460 47124 39488
rect 43855 39457 43867 39460
rect 43809 39451 43867 39457
rect 47118 39448 47124 39460
rect 47176 39448 47182 39500
rect 39850 39420 39856 39432
rect 39811 39392 39856 39420
rect 39850 39380 39856 39392
rect 39908 39380 39914 39432
rect 40037 39423 40095 39429
rect 40037 39389 40049 39423
rect 40083 39389 40095 39423
rect 40037 39383 40095 39389
rect 41141 39423 41199 39429
rect 41141 39389 41153 39423
rect 41187 39420 41199 39423
rect 41506 39420 41512 39432
rect 41187 39392 41512 39420
rect 41187 39389 41199 39392
rect 41141 39383 41199 39389
rect 38654 39352 38660 39364
rect 37700 39324 38660 39352
rect 37700 39312 37706 39324
rect 38654 39312 38660 39324
rect 38712 39312 38718 39364
rect 39114 39352 39120 39364
rect 39075 39324 39120 39352
rect 39114 39312 39120 39324
rect 39172 39312 39178 39364
rect 40052 39352 40080 39383
rect 41506 39380 41512 39392
rect 41564 39420 41570 39432
rect 43257 39423 43315 39429
rect 43257 39420 43269 39423
rect 41564 39392 43269 39420
rect 41564 39380 41570 39392
rect 43257 39389 43269 39392
rect 43303 39389 43315 39423
rect 43257 39383 43315 39389
rect 41598 39352 41604 39364
rect 39868 39324 40080 39352
rect 41559 39324 41604 39352
rect 39868 39296 39896 39324
rect 41598 39312 41604 39324
rect 41656 39352 41662 39364
rect 42058 39352 42064 39364
rect 41656 39324 42064 39352
rect 41656 39312 41662 39324
rect 42058 39312 42064 39324
rect 42116 39312 42122 39364
rect 35342 39284 35348 39296
rect 33560 39256 35020 39284
rect 35303 39256 35348 39284
rect 33560 39244 33566 39256
rect 35342 39244 35348 39256
rect 35400 39244 35406 39296
rect 38289 39287 38347 39293
rect 38289 39253 38301 39287
rect 38335 39284 38347 39287
rect 38746 39284 38752 39296
rect 38335 39256 38752 39284
rect 38335 39253 38347 39256
rect 38289 39247 38347 39253
rect 38746 39244 38752 39256
rect 38804 39244 38810 39296
rect 38917 39287 38975 39293
rect 38917 39253 38929 39287
rect 38963 39284 38975 39287
rect 39850 39284 39856 39296
rect 38963 39256 39856 39284
rect 38963 39253 38975 39256
rect 38917 39247 38975 39253
rect 39850 39244 39856 39256
rect 39908 39244 39914 39296
rect 40586 39284 40592 39296
rect 40547 39256 40592 39284
rect 40586 39244 40592 39256
rect 40644 39244 40650 39296
rect 42702 39284 42708 39296
rect 42663 39256 42708 39284
rect 42702 39244 42708 39256
rect 42760 39244 42766 39296
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 11793 39083 11851 39089
rect 11793 39049 11805 39083
rect 11839 39080 11851 39083
rect 12894 39080 12900 39092
rect 11839 39052 12900 39080
rect 11839 39049 11851 39052
rect 11793 39043 11851 39049
rect 12894 39040 12900 39052
rect 12952 39040 12958 39092
rect 13449 39083 13507 39089
rect 13449 39049 13461 39083
rect 13495 39080 13507 39083
rect 13814 39080 13820 39092
rect 13495 39052 13820 39080
rect 13495 39049 13507 39052
rect 13449 39043 13507 39049
rect 13814 39040 13820 39052
rect 13872 39040 13878 39092
rect 14274 39080 14280 39092
rect 14235 39052 14280 39080
rect 14274 39040 14280 39052
rect 14332 39040 14338 39092
rect 15289 39083 15347 39089
rect 15289 39049 15301 39083
rect 15335 39080 15347 39083
rect 15838 39080 15844 39092
rect 15335 39052 15844 39080
rect 15335 39049 15347 39052
rect 15289 39043 15347 39049
rect 15838 39040 15844 39052
rect 15896 39040 15902 39092
rect 16114 39080 16120 39092
rect 16075 39052 16120 39080
rect 16114 39040 16120 39052
rect 16172 39040 16178 39092
rect 17770 39040 17776 39092
rect 17828 39080 17834 39092
rect 18509 39083 18567 39089
rect 18509 39080 18521 39083
rect 17828 39052 18521 39080
rect 17828 39040 17834 39052
rect 18509 39049 18521 39052
rect 18555 39080 18567 39083
rect 19426 39080 19432 39092
rect 18555 39052 19432 39080
rect 18555 39049 18567 39052
rect 18509 39043 18567 39049
rect 19426 39040 19432 39052
rect 19484 39040 19490 39092
rect 20990 39080 20996 39092
rect 19536 39052 20996 39080
rect 13630 39012 13636 39024
rect 13372 38984 13636 39012
rect 11146 38904 11152 38956
rect 11204 38944 11210 38956
rect 13372 38953 13400 38984
rect 13630 38972 13636 38984
rect 13688 38972 13694 39024
rect 13832 39012 13860 39040
rect 14182 39012 14188 39024
rect 13832 38984 14188 39012
rect 14182 38972 14188 38984
rect 14240 38972 14246 39024
rect 14366 39012 14372 39024
rect 14292 38984 14372 39012
rect 13357 38947 13415 38953
rect 13357 38944 13369 38947
rect 11204 38916 13369 38944
rect 11204 38904 11210 38916
rect 13357 38913 13369 38916
rect 13403 38913 13415 38947
rect 13357 38907 13415 38913
rect 13541 38947 13599 38953
rect 13541 38913 13553 38947
rect 13587 38944 13599 38947
rect 14292 38944 14320 38984
rect 14366 38972 14372 38984
rect 14424 38972 14430 39024
rect 15933 39015 15991 39021
rect 15933 39012 15945 39015
rect 15304 38984 15945 39012
rect 14458 38944 14464 38956
rect 13587 38916 14320 38944
rect 14419 38916 14464 38944
rect 13587 38913 13599 38916
rect 13541 38907 13599 38913
rect 12894 38876 12900 38888
rect 12855 38848 12900 38876
rect 12894 38836 12900 38848
rect 12952 38836 12958 38888
rect 13556 38808 13584 38907
rect 14458 38904 14464 38916
rect 14516 38904 14522 38956
rect 14550 38904 14556 38956
rect 14608 38944 14614 38956
rect 14608 38916 14653 38944
rect 14608 38904 14614 38916
rect 15010 38904 15016 38956
rect 15068 38944 15074 38956
rect 15304 38953 15332 38984
rect 15933 38981 15945 38984
rect 15979 38981 15991 39015
rect 15933 38975 15991 38981
rect 18417 39015 18475 39021
rect 18417 38981 18429 39015
rect 18463 39012 18475 39015
rect 18874 39012 18880 39024
rect 18463 38984 18880 39012
rect 18463 38981 18475 38984
rect 18417 38975 18475 38981
rect 18874 38972 18880 38984
rect 18932 38972 18938 39024
rect 19334 38972 19340 39024
rect 19392 39012 19398 39024
rect 19536 39012 19564 39052
rect 20990 39040 20996 39052
rect 21048 39040 21054 39092
rect 21085 39083 21143 39089
rect 21085 39049 21097 39083
rect 21131 39080 21143 39083
rect 21913 39083 21971 39089
rect 21913 39080 21925 39083
rect 21131 39052 21925 39080
rect 21131 39049 21143 39052
rect 21085 39043 21143 39049
rect 21913 39049 21925 39052
rect 21959 39049 21971 39083
rect 23106 39080 23112 39092
rect 21913 39043 21971 39049
rect 22756 39052 23112 39080
rect 19392 38984 19564 39012
rect 20441 39015 20499 39021
rect 19392 38972 19398 38984
rect 20441 38981 20453 39015
rect 20487 39012 20499 39015
rect 20622 39012 20628 39024
rect 20487 38984 20628 39012
rect 20487 38981 20499 38984
rect 20441 38975 20499 38981
rect 20622 38972 20628 38984
rect 20680 39012 20686 39024
rect 22756 39021 22784 39052
rect 23106 39040 23112 39052
rect 23164 39040 23170 39092
rect 23566 39080 23572 39092
rect 23527 39052 23572 39080
rect 23566 39040 23572 39052
rect 23624 39040 23630 39092
rect 25590 39080 25596 39092
rect 24780 39052 25596 39080
rect 22741 39015 22799 39021
rect 20680 38984 21864 39012
rect 20680 38972 20686 38984
rect 15105 38947 15163 38953
rect 15105 38944 15117 38947
rect 15068 38916 15117 38944
rect 15068 38904 15074 38916
rect 15105 38913 15117 38916
rect 15151 38913 15163 38947
rect 15289 38947 15347 38953
rect 15289 38944 15301 38947
rect 15105 38907 15163 38913
rect 15212 38916 15301 38944
rect 14274 38876 14280 38888
rect 14235 38848 14280 38876
rect 14274 38836 14280 38848
rect 14332 38836 14338 38888
rect 10888 38780 13584 38808
rect 10888 38752 10916 38780
rect 10226 38700 10232 38752
rect 10284 38740 10290 38752
rect 10870 38740 10876 38752
rect 10284 38712 10876 38740
rect 10284 38700 10290 38712
rect 10870 38700 10876 38712
rect 10928 38700 10934 38752
rect 12250 38740 12256 38752
rect 12211 38712 12256 38740
rect 12250 38700 12256 38712
rect 12308 38740 12314 38752
rect 15212 38740 15240 38916
rect 15289 38913 15301 38916
rect 15335 38913 15347 38947
rect 15289 38907 15347 38913
rect 15378 38904 15384 38956
rect 15436 38944 15442 38956
rect 15749 38947 15807 38953
rect 15749 38944 15761 38947
rect 15436 38916 15761 38944
rect 15436 38904 15442 38916
rect 15749 38913 15761 38916
rect 15795 38913 15807 38947
rect 15749 38907 15807 38913
rect 16022 38904 16028 38956
rect 16080 38944 16086 38956
rect 16853 38947 16911 38953
rect 16853 38944 16865 38947
rect 16080 38916 16865 38944
rect 16080 38904 16086 38916
rect 16853 38913 16865 38916
rect 16899 38913 16911 38947
rect 16853 38907 16911 38913
rect 18598 38904 18604 38956
rect 18656 38944 18662 38956
rect 19429 38947 19487 38953
rect 19429 38944 19441 38947
rect 18656 38916 19441 38944
rect 18656 38904 18662 38916
rect 19429 38913 19441 38916
rect 19475 38913 19487 38947
rect 20070 38944 20076 38956
rect 20031 38916 20076 38944
rect 19429 38907 19487 38913
rect 20070 38904 20076 38916
rect 20128 38904 20134 38956
rect 20257 38947 20315 38953
rect 20257 38913 20269 38947
rect 20303 38944 20315 38947
rect 20806 38944 20812 38956
rect 20303 38916 20812 38944
rect 20303 38913 20315 38916
rect 20257 38907 20315 38913
rect 20806 38904 20812 38916
rect 20864 38904 20870 38956
rect 21836 38953 21864 38984
rect 22741 38981 22753 39015
rect 22787 38981 22799 39015
rect 22741 38975 22799 38981
rect 22925 39015 22983 39021
rect 22925 38981 22937 39015
rect 22971 39012 22983 39015
rect 23290 39012 23296 39024
rect 22971 38984 23296 39012
rect 22971 38981 22983 38984
rect 22925 38975 22983 38981
rect 20901 38947 20959 38953
rect 20901 38913 20913 38947
rect 20947 38944 20959 38947
rect 21085 38947 21143 38953
rect 20947 38916 21036 38944
rect 20947 38913 20959 38916
rect 20901 38907 20959 38913
rect 15930 38836 15936 38888
rect 15988 38876 15994 38888
rect 16390 38876 16396 38888
rect 15988 38848 16396 38876
rect 15988 38836 15994 38848
rect 16390 38836 16396 38848
rect 16448 38876 16454 38888
rect 16669 38879 16727 38885
rect 16669 38876 16681 38879
rect 16448 38848 16681 38876
rect 16448 38836 16454 38848
rect 16669 38845 16681 38848
rect 16715 38845 16727 38879
rect 19242 38876 19248 38888
rect 19203 38848 19248 38876
rect 16669 38839 16727 38845
rect 19242 38836 19248 38848
rect 19300 38836 19306 38888
rect 20088 38876 20116 38904
rect 21008 38876 21036 38916
rect 21085 38913 21097 38947
rect 21131 38913 21143 38947
rect 21085 38907 21143 38913
rect 21821 38947 21879 38953
rect 21821 38913 21833 38947
rect 21867 38913 21879 38947
rect 21821 38907 21879 38913
rect 20088 38848 21036 38876
rect 17865 38811 17923 38817
rect 17865 38777 17877 38811
rect 17911 38808 17923 38811
rect 19334 38808 19340 38820
rect 17911 38780 19340 38808
rect 17911 38777 17923 38780
rect 17865 38771 17923 38777
rect 19334 38768 19340 38780
rect 19392 38768 19398 38820
rect 20806 38768 20812 38820
rect 20864 38808 20870 38820
rect 21100 38808 21128 38907
rect 21910 38904 21916 38956
rect 21968 38944 21974 38956
rect 22189 38947 22247 38953
rect 22189 38944 22201 38947
rect 21968 38916 22201 38944
rect 21968 38904 21974 38916
rect 22189 38913 22201 38916
rect 22235 38913 22247 38947
rect 22189 38907 22247 38913
rect 22002 38876 22008 38888
rect 21963 38848 22008 38876
rect 22002 38836 22008 38848
rect 22060 38836 22066 38888
rect 22940 38876 22968 38975
rect 23290 38972 23296 38984
rect 23348 39012 23354 39024
rect 23348 38984 23888 39012
rect 23348 38972 23354 38984
rect 23014 38904 23020 38956
rect 23072 38944 23078 38956
rect 23860 38953 23888 38984
rect 24026 38972 24032 39024
rect 24084 39012 24090 39024
rect 24641 39015 24699 39021
rect 24641 39012 24653 39015
rect 24084 38984 24653 39012
rect 24084 38972 24090 38984
rect 24641 38981 24653 38984
rect 24687 39012 24699 39015
rect 24780 39012 24808 39052
rect 25590 39040 25596 39052
rect 25648 39040 25654 39092
rect 28350 39080 28356 39092
rect 28311 39052 28356 39080
rect 28350 39040 28356 39052
rect 28408 39040 28414 39092
rect 28442 39040 28448 39092
rect 28500 39080 28506 39092
rect 30377 39083 30435 39089
rect 30377 39080 30389 39083
rect 28500 39052 30389 39080
rect 28500 39040 28506 39052
rect 30377 39049 30389 39052
rect 30423 39049 30435 39083
rect 30377 39043 30435 39049
rect 24687 38984 24808 39012
rect 24687 38981 24699 38984
rect 24641 38975 24699 38981
rect 24854 38972 24860 39024
rect 24912 39012 24918 39024
rect 25498 39012 25504 39024
rect 24912 38984 25504 39012
rect 24912 38972 24918 38984
rect 25498 38972 25504 38984
rect 25556 38972 25562 39024
rect 23753 38947 23811 38953
rect 23753 38944 23765 38947
rect 23072 38916 23765 38944
rect 23072 38904 23078 38916
rect 23753 38913 23765 38916
rect 23799 38913 23811 38947
rect 23753 38907 23811 38913
rect 23845 38947 23903 38953
rect 23845 38913 23857 38947
rect 23891 38913 23903 38947
rect 23845 38907 23903 38913
rect 24302 38904 24308 38956
rect 24360 38944 24366 38956
rect 24762 38944 24768 38956
rect 24360 38916 24768 38944
rect 24360 38904 24366 38916
rect 24762 38904 24768 38916
rect 24820 38944 24826 38956
rect 25608 38953 25636 39040
rect 25317 38947 25375 38953
rect 25317 38944 25329 38947
rect 24820 38916 25329 38944
rect 24820 38904 24826 38916
rect 25317 38913 25329 38916
rect 25363 38913 25375 38947
rect 25317 38907 25375 38913
rect 25593 38947 25651 38953
rect 25593 38913 25605 38947
rect 25639 38913 25651 38947
rect 25593 38907 25651 38913
rect 28258 38904 28264 38956
rect 28316 38944 28322 38956
rect 28537 38947 28595 38953
rect 28537 38944 28549 38947
rect 28316 38916 28549 38944
rect 28316 38904 28322 38916
rect 28537 38913 28549 38916
rect 28583 38913 28595 38947
rect 28537 38907 28595 38913
rect 28626 38904 28632 38956
rect 28684 38944 28690 38956
rect 28810 38944 28816 38956
rect 28684 38916 28816 38944
rect 28684 38904 28690 38916
rect 28810 38904 28816 38916
rect 28868 38904 28874 38956
rect 28905 38947 28963 38953
rect 28905 38913 28917 38947
rect 28951 38913 28963 38947
rect 29730 38944 29736 38956
rect 29691 38916 29736 38944
rect 28905 38907 28963 38913
rect 22112 38848 22968 38876
rect 23569 38879 23627 38885
rect 20864 38780 21128 38808
rect 20864 38768 20870 38780
rect 17034 38740 17040 38752
rect 12308 38712 15240 38740
rect 16995 38712 17040 38740
rect 12308 38700 12314 38712
rect 17034 38700 17040 38712
rect 17092 38700 17098 38752
rect 18322 38700 18328 38752
rect 18380 38740 18386 38752
rect 19150 38740 19156 38752
rect 18380 38712 19156 38740
rect 18380 38700 18386 38712
rect 19150 38700 19156 38712
rect 19208 38700 19214 38752
rect 19610 38740 19616 38752
rect 19571 38712 19616 38740
rect 19610 38700 19616 38712
rect 19668 38700 19674 38752
rect 21082 38700 21088 38752
rect 21140 38740 21146 38752
rect 22112 38740 22140 38848
rect 23569 38845 23581 38879
rect 23615 38876 23627 38879
rect 23658 38876 23664 38888
rect 23615 38848 23664 38876
rect 23615 38845 23627 38848
rect 23569 38839 23627 38845
rect 23658 38836 23664 38848
rect 23716 38836 23722 38888
rect 24486 38836 24492 38888
rect 24544 38876 24550 38888
rect 27522 38876 27528 38888
rect 24544 38848 25360 38876
rect 24544 38836 24550 38848
rect 25332 38817 25360 38848
rect 25424 38848 27528 38876
rect 22189 38811 22247 38817
rect 22189 38777 22201 38811
rect 22235 38808 22247 38811
rect 25317 38811 25375 38817
rect 22235 38780 24992 38808
rect 22235 38777 22247 38780
rect 22189 38771 22247 38777
rect 22738 38740 22744 38752
rect 21140 38712 22140 38740
rect 22699 38712 22744 38740
rect 21140 38700 21146 38712
rect 22738 38700 22744 38712
rect 22796 38700 22802 38752
rect 24489 38743 24547 38749
rect 24489 38709 24501 38743
rect 24535 38740 24547 38743
rect 24578 38740 24584 38752
rect 24535 38712 24584 38740
rect 24535 38709 24547 38712
rect 24489 38703 24547 38709
rect 24578 38700 24584 38712
rect 24636 38700 24642 38752
rect 24673 38743 24731 38749
rect 24673 38709 24685 38743
rect 24719 38740 24731 38743
rect 24762 38740 24768 38752
rect 24719 38712 24768 38740
rect 24719 38709 24731 38712
rect 24673 38703 24731 38709
rect 24762 38700 24768 38712
rect 24820 38700 24826 38752
rect 24964 38740 24992 38780
rect 25317 38777 25329 38811
rect 25363 38777 25375 38811
rect 25317 38771 25375 38777
rect 25424 38740 25452 38848
rect 27522 38836 27528 38848
rect 27580 38836 27586 38888
rect 28442 38836 28448 38888
rect 28500 38876 28506 38888
rect 28920 38876 28948 38907
rect 29730 38904 29736 38916
rect 29788 38904 29794 38956
rect 29638 38876 29644 38888
rect 28500 38848 28948 38876
rect 29599 38848 29644 38876
rect 28500 38836 28506 38848
rect 29638 38836 29644 38848
rect 29696 38836 29702 38888
rect 30392 38876 30420 39043
rect 30558 39040 30564 39092
rect 30616 39080 30622 39092
rect 31113 39083 31171 39089
rect 31113 39080 31125 39083
rect 30616 39052 31125 39080
rect 30616 39040 30622 39052
rect 30558 38904 30564 38956
rect 30616 38944 30622 38956
rect 30742 38944 30748 38956
rect 30616 38916 30748 38944
rect 30616 38904 30622 38916
rect 30742 38904 30748 38916
rect 30800 38904 30806 38956
rect 30944 38944 30972 39052
rect 31113 39049 31125 39052
rect 31159 39049 31171 39083
rect 31113 39043 31171 39049
rect 31938 39040 31944 39092
rect 31996 39080 32002 39092
rect 32398 39080 32404 39092
rect 31996 39052 32404 39080
rect 31996 39040 32002 39052
rect 32398 39040 32404 39052
rect 32456 39040 32462 39092
rect 33410 39080 33416 39092
rect 32508 39052 33416 39080
rect 31021 39015 31079 39021
rect 31021 38981 31033 39015
rect 31067 39012 31079 39015
rect 32508 39012 32536 39052
rect 33410 39040 33416 39052
rect 33468 39040 33474 39092
rect 37553 39083 37611 39089
rect 37553 39049 37565 39083
rect 37599 39080 37611 39083
rect 37642 39080 37648 39092
rect 37599 39052 37648 39080
rect 37599 39049 37611 39052
rect 37553 39043 37611 39049
rect 37642 39040 37648 39052
rect 37700 39040 37706 39092
rect 38197 39083 38255 39089
rect 38197 39080 38209 39083
rect 37752 39052 38209 39080
rect 31067 38984 32536 39012
rect 32585 39015 32643 39021
rect 31067 38981 31079 38984
rect 31021 38975 31079 38981
rect 32585 38981 32597 39015
rect 32631 39012 32643 39015
rect 32766 39012 32772 39024
rect 32631 38984 32772 39012
rect 32631 38981 32643 38984
rect 32585 38975 32643 38981
rect 32766 38972 32772 38984
rect 32824 38972 32830 39024
rect 33502 39012 33508 39024
rect 33463 38984 33508 39012
rect 33502 38972 33508 38984
rect 33560 38972 33566 39024
rect 33594 38972 33600 39024
rect 33652 39012 33658 39024
rect 33873 39015 33931 39021
rect 33873 39012 33885 39015
rect 33652 38984 33885 39012
rect 33652 38972 33658 38984
rect 33873 38981 33885 38984
rect 33919 39012 33931 39015
rect 34422 39012 34428 39024
rect 33919 38984 34428 39012
rect 33919 38981 33931 38984
rect 33873 38975 33931 38981
rect 34422 38972 34428 38984
rect 34480 38972 34486 39024
rect 37752 39021 37780 39052
rect 38197 39049 38209 39052
rect 38243 39049 38255 39083
rect 38197 39043 38255 39049
rect 38365 39083 38423 39089
rect 38365 39049 38377 39083
rect 38411 39080 38423 39083
rect 38930 39080 38936 39092
rect 38411 39052 38936 39080
rect 38411 39049 38423 39052
rect 38365 39043 38423 39049
rect 38930 39040 38936 39052
rect 38988 39080 38994 39092
rect 39025 39083 39083 39089
rect 39025 39080 39037 39083
rect 38988 39052 39037 39080
rect 38988 39040 38994 39052
rect 39025 39049 39037 39052
rect 39071 39049 39083 39083
rect 39850 39080 39856 39092
rect 39811 39052 39856 39080
rect 39025 39043 39083 39049
rect 39850 39040 39856 39052
rect 39908 39040 39914 39092
rect 43530 39080 43536 39092
rect 43491 39052 43536 39080
rect 43530 39040 43536 39052
rect 43588 39040 43594 39092
rect 37737 39015 37795 39021
rect 34624 38984 37688 39012
rect 31754 38944 31760 38956
rect 30944 38916 31760 38944
rect 31754 38904 31760 38916
rect 31812 38904 31818 38956
rect 32490 38904 32496 38956
rect 32548 38944 32554 38956
rect 32953 38947 33011 38953
rect 32953 38944 32965 38947
rect 32548 38916 32965 38944
rect 32548 38904 32554 38916
rect 32953 38913 32965 38916
rect 32999 38944 33011 38947
rect 33686 38944 33692 38956
rect 32999 38916 33692 38944
rect 32999 38913 33011 38916
rect 32953 38907 33011 38913
rect 33686 38904 33692 38916
rect 33744 38904 33750 38956
rect 34146 38904 34152 38956
rect 34204 38944 34210 38956
rect 34624 38953 34652 38984
rect 34333 38947 34391 38953
rect 34333 38944 34345 38947
rect 34204 38916 34345 38944
rect 34204 38904 34210 38916
rect 34333 38913 34345 38916
rect 34379 38913 34391 38947
rect 34333 38907 34391 38913
rect 34517 38947 34575 38953
rect 34517 38913 34529 38947
rect 34563 38913 34575 38947
rect 34517 38907 34575 38913
rect 34609 38947 34667 38953
rect 34609 38913 34621 38947
rect 34655 38913 34667 38947
rect 36170 38944 36176 38956
rect 36131 38916 36176 38944
rect 34609 38907 34667 38913
rect 31386 38876 31392 38888
rect 30392 38848 31392 38876
rect 31386 38836 31392 38848
rect 31444 38836 31450 38888
rect 31570 38836 31576 38888
rect 31628 38876 31634 38888
rect 34238 38876 34244 38888
rect 31628 38848 34244 38876
rect 31628 38836 31634 38848
rect 34238 38836 34244 38848
rect 34296 38836 34302 38888
rect 34532 38876 34560 38907
rect 36170 38904 36176 38916
rect 36228 38904 36234 38956
rect 36357 38947 36415 38953
rect 36357 38913 36369 38947
rect 36403 38944 36415 38947
rect 36446 38944 36452 38956
rect 36403 38916 36452 38944
rect 36403 38913 36415 38916
rect 36357 38907 36415 38913
rect 36446 38904 36452 38916
rect 36504 38904 36510 38956
rect 37461 38947 37519 38953
rect 37461 38913 37473 38947
rect 37507 38913 37519 38947
rect 37660 38944 37688 38984
rect 37737 38981 37749 39015
rect 37783 38981 37795 39015
rect 38562 39012 38568 39024
rect 38523 38984 38568 39012
rect 37737 38975 37795 38981
rect 38562 38972 38568 38984
rect 38620 38972 38626 39024
rect 38654 38972 38660 39024
rect 38712 39012 38718 39024
rect 39209 39015 39267 39021
rect 39209 39012 39221 39015
rect 38712 38984 39221 39012
rect 38712 38972 38718 38984
rect 39209 38981 39221 38984
rect 39255 38981 39267 39015
rect 39209 38975 39267 38981
rect 39482 38972 39488 39024
rect 39540 39012 39546 39024
rect 40037 39015 40095 39021
rect 40037 39012 40049 39015
rect 39540 38984 40049 39012
rect 39540 38972 39546 38984
rect 40037 38981 40049 38984
rect 40083 39012 40095 39015
rect 43162 39012 43168 39024
rect 40083 38984 43168 39012
rect 40083 38981 40095 38984
rect 40037 38975 40095 38981
rect 43162 38972 43168 38984
rect 43220 38972 43226 39024
rect 39022 38944 39028 38956
rect 37660 38916 39028 38944
rect 37461 38907 37519 38913
rect 35710 38876 35716 38888
rect 34532 38848 35716 38876
rect 35710 38836 35716 38848
rect 35768 38836 35774 38888
rect 37476 38876 37504 38907
rect 39022 38904 39028 38916
rect 39080 38904 39086 38956
rect 39393 38947 39451 38953
rect 39393 38913 39405 38947
rect 39439 38913 39451 38947
rect 40218 38944 40224 38956
rect 40131 38916 40224 38944
rect 39393 38907 39451 38913
rect 38102 38876 38108 38888
rect 37476 38848 38108 38876
rect 38102 38836 38108 38848
rect 38160 38876 38166 38888
rect 39408 38876 39436 38907
rect 40218 38904 40224 38916
rect 40276 38944 40282 38956
rect 40862 38944 40868 38956
rect 40276 38916 40868 38944
rect 40276 38904 40282 38916
rect 40862 38904 40868 38916
rect 40920 38904 40926 38956
rect 41785 38879 41843 38885
rect 41785 38876 41797 38879
rect 38160 38848 41797 38876
rect 38160 38836 38166 38848
rect 41785 38845 41797 38848
rect 41831 38876 41843 38879
rect 42702 38876 42708 38888
rect 41831 38848 42708 38876
rect 41831 38845 41843 38848
rect 41785 38839 41843 38845
rect 42702 38836 42708 38848
rect 42760 38836 42766 38888
rect 27433 38811 27491 38817
rect 27433 38777 27445 38811
rect 27479 38808 27491 38811
rect 28166 38808 28172 38820
rect 27479 38780 28172 38808
rect 27479 38777 27491 38780
rect 27433 38771 27491 38777
rect 28166 38768 28172 38780
rect 28224 38768 28230 38820
rect 29086 38808 29092 38820
rect 28736 38780 29092 38808
rect 24964 38712 25452 38740
rect 26234 38700 26240 38752
rect 26292 38740 26298 38752
rect 26329 38743 26387 38749
rect 26329 38740 26341 38743
rect 26292 38712 26341 38740
rect 26292 38700 26298 38712
rect 26329 38709 26341 38712
rect 26375 38740 26387 38743
rect 27246 38740 27252 38752
rect 26375 38712 27252 38740
rect 26375 38709 26387 38712
rect 26329 38703 26387 38709
rect 27246 38700 27252 38712
rect 27304 38740 27310 38752
rect 28736 38740 28764 38780
rect 29086 38768 29092 38780
rect 29144 38768 29150 38820
rect 29454 38768 29460 38820
rect 29512 38808 29518 38820
rect 32398 38808 32404 38820
rect 29512 38780 32404 38808
rect 29512 38768 29518 38780
rect 32398 38768 32404 38780
rect 32456 38808 32462 38820
rect 32858 38808 32864 38820
rect 32456 38780 32864 38808
rect 32456 38768 32462 38780
rect 32858 38768 32864 38780
rect 32916 38768 32922 38820
rect 33686 38768 33692 38820
rect 33744 38808 33750 38820
rect 38010 38808 38016 38820
rect 33744 38780 38016 38808
rect 33744 38768 33750 38780
rect 38010 38768 38016 38780
rect 38068 38768 38074 38820
rect 41233 38811 41291 38817
rect 41233 38808 41245 38811
rect 38396 38780 41245 38808
rect 27304 38712 28764 38740
rect 28813 38743 28871 38749
rect 27304 38700 27310 38712
rect 28813 38709 28825 38743
rect 28859 38740 28871 38743
rect 29365 38743 29423 38749
rect 29365 38740 29377 38743
rect 28859 38712 29377 38740
rect 28859 38709 28871 38712
rect 28813 38703 28871 38709
rect 29365 38709 29377 38712
rect 29411 38709 29423 38743
rect 29365 38703 29423 38709
rect 30558 38700 30564 38752
rect 30616 38740 30622 38752
rect 31294 38740 31300 38752
rect 30616 38712 31300 38740
rect 30616 38700 30622 38712
rect 31294 38700 31300 38712
rect 31352 38700 31358 38752
rect 32306 38700 32312 38752
rect 32364 38740 32370 38752
rect 33594 38740 33600 38752
rect 32364 38712 33600 38740
rect 32364 38700 32370 38712
rect 33594 38700 33600 38712
rect 33652 38700 33658 38752
rect 34330 38740 34336 38752
rect 34291 38712 34336 38740
rect 34330 38700 34336 38712
rect 34388 38700 34394 38752
rect 35161 38743 35219 38749
rect 35161 38709 35173 38743
rect 35207 38740 35219 38743
rect 35434 38740 35440 38752
rect 35207 38712 35440 38740
rect 35207 38709 35219 38712
rect 35161 38703 35219 38709
rect 35434 38700 35440 38712
rect 35492 38700 35498 38752
rect 35710 38740 35716 38752
rect 35671 38712 35716 38740
rect 35710 38700 35716 38712
rect 35768 38700 35774 38752
rect 36262 38740 36268 38752
rect 36223 38712 36268 38740
rect 36262 38700 36268 38712
rect 36320 38700 36326 38752
rect 37737 38743 37795 38749
rect 37737 38709 37749 38743
rect 37783 38740 37795 38743
rect 38194 38740 38200 38752
rect 37783 38712 38200 38740
rect 37783 38709 37795 38712
rect 37737 38703 37795 38709
rect 38194 38700 38200 38712
rect 38252 38700 38258 38752
rect 38396 38749 38424 38780
rect 41233 38777 41245 38780
rect 41279 38808 41291 38811
rect 41279 38780 41414 38808
rect 41279 38777 41291 38780
rect 41233 38771 41291 38777
rect 38381 38743 38439 38749
rect 38381 38709 38393 38743
rect 38427 38709 38439 38743
rect 38381 38703 38439 38709
rect 39666 38700 39672 38752
rect 39724 38740 39730 38752
rect 40681 38743 40739 38749
rect 40681 38740 40693 38743
rect 39724 38712 40693 38740
rect 39724 38700 39730 38712
rect 40681 38709 40693 38712
rect 40727 38709 40739 38743
rect 41386 38740 41414 38780
rect 42521 38743 42579 38749
rect 42521 38740 42533 38743
rect 41386 38712 42533 38740
rect 40681 38703 40739 38709
rect 42521 38709 42533 38712
rect 42567 38740 42579 38743
rect 42702 38740 42708 38752
rect 42567 38712 42708 38740
rect 42567 38709 42579 38712
rect 42521 38703 42579 38709
rect 42702 38700 42708 38712
rect 42760 38700 42766 38752
rect 42978 38740 42984 38752
rect 42939 38712 42984 38740
rect 42978 38700 42984 38712
rect 43036 38700 43042 38752
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 11146 38496 11152 38548
rect 11204 38536 11210 38548
rect 11241 38539 11299 38545
rect 11241 38536 11253 38539
rect 11204 38508 11253 38536
rect 11204 38496 11210 38508
rect 11241 38505 11253 38508
rect 11287 38505 11299 38539
rect 11241 38499 11299 38505
rect 14090 38496 14096 38548
rect 14148 38536 14154 38548
rect 14185 38539 14243 38545
rect 14185 38536 14197 38539
rect 14148 38508 14197 38536
rect 14148 38496 14154 38508
rect 14185 38505 14197 38508
rect 14231 38505 14243 38539
rect 14185 38499 14243 38505
rect 14458 38496 14464 38548
rect 14516 38536 14522 38548
rect 14737 38539 14795 38545
rect 14737 38536 14749 38539
rect 14516 38508 14749 38536
rect 14516 38496 14522 38508
rect 14737 38505 14749 38508
rect 14783 38505 14795 38539
rect 14737 38499 14795 38505
rect 15933 38539 15991 38545
rect 15933 38505 15945 38539
rect 15979 38505 15991 38539
rect 16666 38536 16672 38548
rect 16579 38508 16672 38536
rect 15933 38499 15991 38505
rect 13446 38428 13452 38480
rect 13504 38468 13510 38480
rect 13541 38471 13599 38477
rect 13541 38468 13553 38471
rect 13504 38440 13553 38468
rect 13504 38428 13510 38440
rect 13541 38437 13553 38440
rect 13587 38468 13599 38471
rect 15654 38468 15660 38480
rect 13587 38440 15660 38468
rect 13587 38437 13599 38440
rect 13541 38431 13599 38437
rect 15654 38428 15660 38440
rect 15712 38428 15718 38480
rect 15746 38400 15752 38412
rect 15707 38372 15752 38400
rect 15746 38360 15752 38372
rect 15804 38360 15810 38412
rect 15948 38400 15976 38499
rect 16666 38496 16672 38508
rect 16724 38536 16730 38548
rect 17034 38536 17040 38548
rect 16724 38508 17040 38536
rect 16724 38496 16730 38508
rect 17034 38496 17040 38508
rect 17092 38496 17098 38548
rect 17681 38539 17739 38545
rect 17681 38505 17693 38539
rect 17727 38536 17739 38539
rect 19242 38536 19248 38548
rect 17727 38508 19248 38536
rect 17727 38505 17739 38508
rect 17681 38499 17739 38505
rect 19242 38496 19248 38508
rect 19300 38496 19306 38548
rect 19889 38539 19947 38545
rect 19889 38505 19901 38539
rect 19935 38536 19947 38539
rect 20346 38536 20352 38548
rect 19935 38508 20352 38536
rect 19935 38505 19947 38508
rect 19889 38499 19947 38505
rect 20346 38496 20352 38508
rect 20404 38496 20410 38548
rect 20530 38536 20536 38548
rect 20491 38508 20536 38536
rect 20530 38496 20536 38508
rect 20588 38496 20594 38548
rect 21910 38496 21916 38548
rect 21968 38536 21974 38548
rect 22005 38539 22063 38545
rect 22005 38536 22017 38539
rect 21968 38508 22017 38536
rect 21968 38496 21974 38508
rect 22005 38505 22017 38508
rect 22051 38505 22063 38539
rect 22005 38499 22063 38505
rect 22235 38539 22293 38545
rect 22235 38505 22247 38539
rect 22281 38536 22293 38539
rect 22738 38536 22744 38548
rect 22281 38508 22744 38536
rect 22281 38505 22293 38508
rect 22235 38499 22293 38505
rect 22738 38496 22744 38508
rect 22796 38496 22802 38548
rect 22830 38496 22836 38548
rect 22888 38536 22894 38548
rect 23109 38539 23167 38545
rect 23109 38536 23121 38539
rect 22888 38508 23121 38536
rect 22888 38496 22894 38508
rect 23109 38505 23121 38508
rect 23155 38536 23167 38539
rect 23198 38536 23204 38548
rect 23155 38508 23204 38536
rect 23155 38505 23167 38508
rect 23109 38499 23167 38505
rect 23198 38496 23204 38508
rect 23256 38496 23262 38548
rect 23842 38536 23848 38548
rect 23803 38508 23848 38536
rect 23842 38496 23848 38508
rect 23900 38496 23906 38548
rect 25133 38539 25191 38545
rect 25133 38505 25145 38539
rect 25179 38536 25191 38539
rect 25314 38536 25320 38548
rect 25179 38508 25320 38536
rect 25179 38505 25191 38508
rect 25133 38499 25191 38505
rect 25314 38496 25320 38508
rect 25372 38496 25378 38548
rect 25406 38496 25412 38548
rect 25464 38536 25470 38548
rect 27798 38536 27804 38548
rect 25464 38508 27804 38536
rect 25464 38496 25470 38508
rect 27798 38496 27804 38508
rect 27856 38496 27862 38548
rect 27982 38536 27988 38548
rect 27943 38508 27988 38536
rect 27982 38496 27988 38508
rect 28040 38496 28046 38548
rect 28905 38539 28963 38545
rect 28905 38505 28917 38539
rect 28951 38536 28963 38539
rect 29638 38536 29644 38548
rect 28951 38508 29644 38536
rect 28951 38505 28963 38508
rect 28905 38499 28963 38505
rect 29638 38496 29644 38508
rect 29696 38496 29702 38548
rect 30374 38496 30380 38548
rect 30432 38536 30438 38548
rect 32493 38539 32551 38545
rect 32493 38536 32505 38539
rect 30432 38508 32505 38536
rect 30432 38496 30438 38508
rect 32493 38505 32505 38508
rect 32539 38505 32551 38539
rect 32493 38499 32551 38505
rect 32858 38496 32864 38548
rect 32916 38536 32922 38548
rect 32916 38508 33916 38536
rect 32916 38496 32922 38508
rect 16022 38428 16028 38480
rect 16080 38468 16086 38480
rect 18598 38468 18604 38480
rect 16080 38440 18604 38468
rect 16080 38428 16086 38440
rect 18598 38428 18604 38440
rect 18656 38428 18662 38480
rect 19150 38428 19156 38480
rect 19208 38468 19214 38480
rect 21361 38471 21419 38477
rect 21361 38468 21373 38471
rect 19208 38440 21373 38468
rect 19208 38428 19214 38440
rect 21361 38437 21373 38440
rect 21407 38468 21419 38471
rect 21818 38468 21824 38480
rect 21407 38440 21824 38468
rect 21407 38437 21419 38440
rect 21361 38431 21419 38437
rect 21818 38428 21824 38440
rect 21876 38428 21882 38480
rect 22097 38471 22155 38477
rect 22097 38437 22109 38471
rect 22143 38468 22155 38471
rect 23014 38468 23020 38480
rect 22143 38440 23020 38468
rect 22143 38437 22155 38440
rect 22097 38431 22155 38437
rect 23014 38428 23020 38440
rect 23072 38468 23078 38480
rect 23293 38471 23351 38477
rect 23293 38468 23305 38471
rect 23072 38440 23305 38468
rect 23072 38428 23078 38440
rect 23293 38437 23305 38440
rect 23339 38437 23351 38471
rect 27706 38468 27712 38480
rect 23293 38431 23351 38437
rect 24688 38440 27712 38468
rect 16482 38400 16488 38412
rect 15948 38372 16488 38400
rect 16482 38360 16488 38372
rect 16540 38400 16546 38412
rect 16577 38403 16635 38409
rect 16577 38400 16589 38403
rect 16540 38372 16589 38400
rect 16540 38360 16546 38372
rect 16577 38369 16589 38372
rect 16623 38369 16635 38403
rect 18138 38400 18144 38412
rect 16577 38363 16635 38369
rect 17788 38372 18144 38400
rect 2041 38335 2099 38341
rect 2041 38301 2053 38335
rect 2087 38332 2099 38335
rect 12250 38332 12256 38344
rect 2087 38304 12256 38332
rect 2087 38301 2099 38304
rect 2041 38295 2099 38301
rect 12250 38292 12256 38304
rect 12308 38332 12314 38344
rect 12526 38332 12532 38344
rect 12308 38304 12532 38332
rect 12308 38292 12314 38304
rect 12526 38292 12532 38304
rect 12584 38292 12590 38344
rect 14921 38335 14979 38341
rect 14921 38301 14933 38335
rect 14967 38332 14979 38335
rect 15102 38332 15108 38344
rect 14967 38304 15108 38332
rect 14967 38301 14979 38304
rect 14921 38295 14979 38301
rect 15102 38292 15108 38304
rect 15160 38292 15166 38344
rect 15197 38335 15255 38341
rect 15197 38301 15209 38335
rect 15243 38332 15255 38335
rect 15286 38332 15292 38344
rect 15243 38304 15292 38332
rect 15243 38301 15255 38304
rect 15197 38295 15255 38301
rect 15286 38292 15292 38304
rect 15344 38292 15350 38344
rect 15933 38335 15991 38341
rect 15933 38301 15945 38335
rect 15979 38301 15991 38335
rect 16850 38332 16856 38344
rect 16811 38304 16856 38332
rect 15933 38295 15991 38301
rect 1578 38224 1584 38276
rect 1636 38264 1642 38276
rect 1857 38267 1915 38273
rect 1857 38264 1869 38267
rect 1636 38236 1869 38264
rect 1636 38224 1642 38236
rect 1857 38233 1869 38236
rect 1903 38233 1915 38267
rect 1857 38227 1915 38233
rect 11885 38267 11943 38273
rect 11885 38233 11897 38267
rect 11931 38264 11943 38267
rect 12989 38267 13047 38273
rect 11931 38236 12940 38264
rect 11931 38233 11943 38236
rect 11885 38227 11943 38233
rect 12434 38156 12440 38208
rect 12492 38196 12498 38208
rect 12912 38196 12940 38236
rect 12989 38233 13001 38267
rect 13035 38264 13047 38267
rect 13814 38264 13820 38276
rect 13035 38236 13820 38264
rect 13035 38233 13047 38236
rect 12989 38227 13047 38233
rect 13814 38224 13820 38236
rect 13872 38224 13878 38276
rect 14642 38224 14648 38276
rect 14700 38264 14706 38276
rect 15470 38264 15476 38276
rect 14700 38236 15476 38264
rect 14700 38224 14706 38236
rect 15470 38224 15476 38236
rect 15528 38264 15534 38276
rect 15657 38267 15715 38273
rect 15657 38264 15669 38267
rect 15528 38236 15669 38264
rect 15528 38224 15534 38236
rect 15657 38233 15669 38236
rect 15703 38233 15715 38267
rect 15948 38264 15976 38295
rect 16850 38292 16856 38304
rect 16908 38292 16914 38344
rect 17586 38332 17592 38344
rect 17547 38304 17592 38332
rect 17586 38292 17592 38304
rect 17644 38292 17650 38344
rect 17788 38341 17816 38372
rect 18138 38360 18144 38372
rect 18196 38360 18202 38412
rect 18230 38360 18236 38412
rect 18288 38400 18294 38412
rect 24688 38409 24716 38440
rect 24673 38403 24731 38409
rect 18288 38372 24624 38400
rect 18288 38360 18294 38372
rect 17773 38335 17831 38341
rect 17773 38301 17785 38335
rect 17819 38301 17831 38335
rect 17773 38295 17831 38301
rect 18417 38335 18475 38341
rect 18417 38301 18429 38335
rect 18463 38332 18475 38335
rect 18506 38332 18512 38344
rect 18463 38304 18512 38332
rect 18463 38301 18475 38304
rect 18417 38295 18475 38301
rect 18506 38292 18512 38304
rect 18564 38292 18570 38344
rect 19797 38335 19855 38341
rect 19797 38301 19809 38335
rect 19843 38332 19855 38335
rect 19886 38332 19892 38344
rect 19843 38304 19892 38332
rect 19843 38301 19855 38304
rect 19797 38295 19855 38301
rect 19886 38292 19892 38304
rect 19944 38292 19950 38344
rect 19981 38335 20039 38341
rect 19981 38301 19993 38335
rect 20027 38332 20039 38335
rect 20162 38332 20168 38344
rect 20027 38304 20168 38332
rect 20027 38301 20039 38304
rect 19981 38295 20039 38301
rect 20162 38292 20168 38304
rect 20220 38292 20226 38344
rect 20438 38332 20444 38344
rect 20399 38304 20444 38332
rect 20438 38292 20444 38304
rect 20496 38292 20502 38344
rect 20625 38335 20683 38341
rect 20625 38301 20637 38335
rect 20671 38332 20683 38335
rect 20714 38332 20720 38344
rect 20671 38304 20720 38332
rect 20671 38301 20683 38304
rect 20625 38295 20683 38301
rect 20714 38292 20720 38304
rect 20772 38292 20778 38344
rect 21910 38332 21916 38344
rect 21871 38304 21916 38332
rect 21910 38292 21916 38304
rect 21968 38292 21974 38344
rect 22278 38292 22284 38344
rect 22336 38332 22342 38344
rect 22373 38335 22431 38341
rect 22373 38332 22385 38335
rect 22336 38304 22385 38332
rect 22336 38292 22342 38304
rect 22373 38301 22385 38304
rect 22419 38301 22431 38335
rect 23290 38332 23296 38344
rect 22373 38295 22431 38301
rect 22940 38304 23296 38332
rect 16206 38264 16212 38276
rect 15948 38236 16212 38264
rect 15657 38227 15715 38233
rect 16206 38224 16212 38236
rect 16264 38264 16270 38276
rect 17604 38264 17632 38292
rect 16264 38236 17632 38264
rect 16264 38224 16270 38236
rect 18138 38224 18144 38276
rect 18196 38264 18202 38276
rect 18233 38267 18291 38273
rect 18233 38264 18245 38267
rect 18196 38236 18245 38264
rect 18196 38224 18202 38236
rect 18233 38233 18245 38236
rect 18279 38264 18291 38267
rect 18966 38264 18972 38276
rect 18279 38236 18972 38264
rect 18279 38233 18291 38236
rect 18233 38227 18291 38233
rect 18966 38224 18972 38236
rect 19024 38224 19030 38276
rect 19904 38264 19932 38292
rect 22830 38264 22836 38276
rect 19904 38236 22836 38264
rect 22830 38224 22836 38236
rect 22888 38224 22894 38276
rect 22940 38273 22968 38304
rect 23290 38292 23296 38304
rect 23348 38292 23354 38344
rect 23474 38292 23480 38344
rect 23532 38332 23538 38344
rect 24596 38341 24624 38372
rect 24673 38369 24685 38403
rect 24719 38369 24731 38403
rect 24673 38363 24731 38369
rect 25685 38403 25743 38409
rect 25685 38369 25697 38403
rect 25731 38400 25743 38403
rect 26326 38400 26332 38412
rect 25731 38372 26332 38400
rect 25731 38369 25743 38372
rect 25685 38363 25743 38369
rect 26326 38360 26332 38372
rect 26384 38360 26390 38412
rect 26513 38403 26571 38409
rect 26513 38369 26525 38403
rect 26559 38400 26571 38403
rect 27062 38400 27068 38412
rect 26559 38372 27068 38400
rect 26559 38369 26571 38372
rect 26513 38363 26571 38369
rect 27062 38360 27068 38372
rect 27120 38360 27126 38412
rect 27540 38409 27568 38440
rect 27706 38428 27712 38440
rect 27764 38468 27770 38480
rect 28442 38468 28448 38480
rect 27764 38440 28448 38468
rect 27764 38428 27770 38440
rect 28442 38428 28448 38440
rect 28500 38428 28506 38480
rect 28813 38471 28871 38477
rect 28813 38437 28825 38471
rect 28859 38468 28871 38471
rect 29825 38471 29883 38477
rect 29825 38468 29837 38471
rect 28859 38440 29837 38468
rect 28859 38437 28871 38440
rect 28813 38431 28871 38437
rect 29825 38437 29837 38440
rect 29871 38468 29883 38471
rect 29871 38440 31340 38468
rect 29871 38437 29883 38440
rect 29825 38431 29883 38437
rect 27525 38403 27583 38409
rect 27525 38369 27537 38403
rect 27571 38369 27583 38403
rect 28994 38400 29000 38412
rect 28955 38372 29000 38400
rect 27525 38363 27583 38369
rect 28994 38360 29000 38372
rect 29052 38360 29058 38412
rect 31312 38409 31340 38440
rect 33594 38428 33600 38480
rect 33652 38468 33658 38480
rect 33781 38471 33839 38477
rect 33781 38468 33793 38471
rect 33652 38440 33793 38468
rect 33652 38428 33658 38440
rect 33781 38437 33793 38440
rect 33827 38437 33839 38471
rect 33888 38468 33916 38508
rect 33962 38496 33968 38548
rect 34020 38536 34026 38548
rect 34701 38539 34759 38545
rect 34701 38536 34713 38539
rect 34020 38508 34713 38536
rect 34020 38496 34026 38508
rect 34701 38505 34713 38508
rect 34747 38505 34759 38539
rect 40405 38539 40463 38545
rect 40405 38536 40417 38539
rect 34701 38499 34759 38505
rect 34808 38508 40417 38536
rect 34808 38468 34836 38508
rect 40405 38505 40417 38508
rect 40451 38505 40463 38539
rect 42610 38536 42616 38548
rect 42571 38508 42616 38536
rect 40405 38499 40463 38505
rect 42610 38496 42616 38508
rect 42668 38496 42674 38548
rect 33888 38440 34836 38468
rect 33781 38431 33839 38437
rect 36354 38428 36360 38480
rect 36412 38468 36418 38480
rect 37737 38471 37795 38477
rect 37737 38468 37749 38471
rect 36412 38440 37749 38468
rect 36412 38428 36418 38440
rect 37737 38437 37749 38440
rect 37783 38437 37795 38471
rect 38841 38471 38899 38477
rect 38841 38468 38853 38471
rect 37737 38431 37795 38437
rect 38120 38440 38853 38468
rect 31297 38403 31355 38409
rect 29472 38372 29960 38400
rect 24397 38335 24455 38341
rect 24397 38332 24409 38335
rect 23532 38304 24409 38332
rect 23532 38292 23538 38304
rect 24397 38301 24409 38304
rect 24443 38301 24455 38335
rect 24397 38295 24455 38301
rect 24581 38335 24639 38341
rect 24581 38301 24593 38335
rect 24627 38301 24639 38335
rect 24581 38295 24639 38301
rect 22925 38267 22983 38273
rect 22925 38233 22937 38267
rect 22971 38233 22983 38267
rect 22925 38227 22983 38233
rect 13170 38196 13176 38208
rect 12492 38168 12537 38196
rect 12912 38168 13176 38196
rect 12492 38156 12498 38168
rect 13170 38156 13176 38168
rect 13228 38156 13234 38208
rect 15105 38199 15163 38205
rect 15105 38165 15117 38199
rect 15151 38196 15163 38199
rect 16022 38196 16028 38208
rect 15151 38168 16028 38196
rect 15151 38165 15163 38168
rect 15105 38159 15163 38165
rect 16022 38156 16028 38168
rect 16080 38156 16086 38208
rect 16114 38156 16120 38208
rect 16172 38196 16178 38208
rect 17034 38196 17040 38208
rect 16172 38168 16217 38196
rect 16995 38168 17040 38196
rect 16172 38156 16178 38168
rect 17034 38156 17040 38168
rect 17092 38156 17098 38208
rect 17954 38156 17960 38208
rect 18012 38196 18018 38208
rect 19337 38199 19395 38205
rect 19337 38196 19349 38199
rect 18012 38168 19349 38196
rect 18012 38156 18018 38168
rect 19337 38165 19349 38168
rect 19383 38196 19395 38199
rect 21818 38196 21824 38208
rect 19383 38168 21824 38196
rect 19383 38165 19395 38168
rect 19337 38159 19395 38165
rect 21818 38156 21824 38168
rect 21876 38156 21882 38208
rect 23106 38156 23112 38208
rect 23164 38205 23170 38208
rect 23164 38199 23183 38205
rect 23171 38165 23183 38199
rect 23164 38159 23183 38165
rect 23164 38156 23170 38159
rect 23290 38156 23296 38208
rect 23348 38196 23354 38208
rect 24302 38196 24308 38208
rect 23348 38168 24308 38196
rect 23348 38156 23354 38168
rect 24302 38156 24308 38168
rect 24360 38156 24366 38208
rect 24412 38196 24440 38295
rect 24762 38292 24768 38344
rect 24820 38332 24826 38344
rect 24820 38304 24865 38332
rect 24820 38292 24826 38304
rect 24946 38292 24952 38344
rect 25004 38332 25010 38344
rect 25406 38332 25412 38344
rect 25004 38304 25412 38332
rect 25004 38292 25010 38304
rect 25406 38292 25412 38304
rect 25464 38292 25470 38344
rect 26421 38335 26479 38341
rect 26421 38301 26433 38335
rect 26467 38332 26479 38335
rect 26694 38332 26700 38344
rect 26467 38304 26700 38332
rect 26467 38301 26479 38304
rect 26421 38295 26479 38301
rect 26694 38292 26700 38304
rect 26752 38292 26758 38344
rect 27246 38332 27252 38344
rect 27207 38304 27252 38332
rect 27246 38292 27252 38304
rect 27304 38292 27310 38344
rect 27430 38332 27436 38344
rect 27391 38304 27436 38332
rect 27430 38292 27436 38304
rect 27488 38292 27494 38344
rect 27614 38292 27620 38344
rect 27672 38332 27678 38344
rect 27672 38304 27717 38332
rect 27672 38292 27678 38304
rect 27798 38292 27804 38344
rect 27856 38332 27862 38344
rect 28626 38332 28632 38344
rect 27856 38304 28632 38332
rect 27856 38292 27862 38304
rect 28626 38292 28632 38304
rect 28684 38292 28690 38344
rect 28721 38335 28779 38341
rect 28721 38301 28733 38335
rect 28767 38332 28779 38335
rect 29472 38332 29500 38372
rect 29638 38332 29644 38344
rect 28767 38304 29500 38332
rect 29599 38304 29644 38332
rect 28767 38301 28779 38304
rect 28721 38295 28779 38301
rect 29638 38292 29644 38304
rect 29696 38292 29702 38344
rect 29730 38292 29736 38344
rect 29788 38332 29794 38344
rect 29932 38341 29960 38372
rect 31297 38369 31309 38403
rect 31343 38400 31355 38403
rect 31386 38400 31392 38412
rect 31343 38372 31392 38400
rect 31343 38369 31355 38372
rect 31297 38363 31355 38369
rect 31386 38360 31392 38372
rect 31444 38360 31450 38412
rect 32953 38403 33011 38409
rect 31726 38372 32812 38400
rect 29917 38335 29975 38341
rect 29788 38304 29833 38332
rect 29788 38292 29794 38304
rect 29917 38301 29929 38335
rect 29963 38332 29975 38335
rect 30190 38332 30196 38344
rect 29963 38304 30196 38332
rect 29963 38301 29975 38304
rect 29917 38295 29975 38301
rect 30190 38292 30196 38304
rect 30248 38332 30254 38344
rect 31205 38335 31263 38341
rect 31205 38332 31217 38335
rect 30248 38304 31217 38332
rect 30248 38292 30254 38304
rect 31205 38301 31217 38304
rect 31251 38301 31263 38335
rect 31205 38295 31263 38301
rect 28442 38224 28448 38276
rect 28500 38264 28506 38276
rect 31726 38264 31754 38372
rect 32784 38344 32812 38372
rect 32953 38369 32965 38403
rect 32999 38400 33011 38403
rect 33226 38400 33232 38412
rect 32999 38372 33232 38400
rect 32999 38369 33011 38372
rect 32953 38363 33011 38369
rect 33226 38360 33232 38372
rect 33284 38360 33290 38412
rect 34885 38403 34943 38409
rect 34885 38369 34897 38403
rect 34931 38369 34943 38403
rect 35066 38400 35072 38412
rect 35027 38372 35072 38400
rect 34885 38363 34943 38369
rect 32677 38335 32735 38341
rect 32677 38301 32689 38335
rect 32723 38301 32735 38335
rect 32677 38295 32735 38301
rect 28500 38236 31754 38264
rect 32692 38264 32720 38295
rect 32766 38292 32772 38344
rect 32824 38332 32830 38344
rect 33042 38332 33048 38344
rect 32824 38304 32869 38332
rect 33003 38304 33048 38332
rect 32824 38292 32830 38304
rect 33042 38292 33048 38304
rect 33100 38292 33106 38344
rect 33134 38292 33140 38344
rect 33192 38332 33198 38344
rect 33505 38335 33563 38341
rect 33505 38332 33517 38335
rect 33192 38304 33517 38332
rect 33192 38292 33198 38304
rect 33505 38301 33517 38304
rect 33551 38301 33563 38335
rect 33505 38295 33563 38301
rect 33597 38335 33655 38341
rect 33597 38301 33609 38335
rect 33643 38332 33655 38335
rect 33686 38332 33692 38344
rect 33643 38304 33692 38332
rect 33643 38301 33655 38304
rect 33597 38295 33655 38301
rect 33686 38292 33692 38304
rect 33744 38292 33750 38344
rect 34900 38334 34928 38363
rect 35066 38360 35072 38372
rect 35124 38360 35130 38412
rect 35161 38403 35219 38409
rect 35161 38369 35173 38403
rect 35207 38400 35219 38403
rect 35342 38400 35348 38412
rect 35207 38372 35348 38400
rect 35207 38369 35219 38372
rect 35161 38363 35219 38369
rect 35342 38360 35348 38372
rect 35400 38360 35406 38412
rect 35710 38360 35716 38412
rect 35768 38400 35774 38412
rect 35989 38403 36047 38409
rect 35989 38400 36001 38403
rect 35768 38372 36001 38400
rect 35768 38360 35774 38372
rect 35989 38369 36001 38372
rect 36035 38369 36047 38403
rect 35989 38363 36047 38369
rect 37185 38403 37243 38409
rect 37185 38369 37197 38403
rect 37231 38400 37243 38403
rect 37366 38400 37372 38412
rect 37231 38372 37372 38400
rect 37231 38369 37243 38372
rect 37185 38363 37243 38369
rect 37366 38360 37372 38372
rect 37424 38400 37430 38412
rect 38013 38403 38071 38409
rect 38013 38400 38025 38403
rect 37424 38372 38025 38400
rect 37424 38360 37430 38372
rect 38013 38369 38025 38372
rect 38059 38369 38071 38403
rect 38013 38363 38071 38369
rect 34977 38335 35035 38341
rect 34900 38306 34929 38334
rect 34901 38276 34929 38306
rect 34977 38301 34989 38335
rect 35023 38301 35035 38335
rect 35084 38332 35112 38360
rect 38120 38344 38148 38440
rect 38841 38437 38853 38440
rect 38887 38437 38899 38471
rect 38841 38431 38899 38437
rect 42153 38471 42211 38477
rect 42153 38437 42165 38471
rect 42199 38468 42211 38471
rect 42978 38468 42984 38480
rect 42199 38440 42984 38468
rect 42199 38437 42211 38440
rect 42153 38431 42211 38437
rect 38562 38360 38568 38412
rect 38620 38400 38626 38412
rect 42168 38400 42196 38431
rect 42978 38428 42984 38440
rect 43036 38428 43042 38480
rect 38620 38372 42196 38400
rect 38620 38360 38626 38372
rect 35084 38304 36032 38332
rect 34977 38295 35035 38301
rect 32692 38236 33088 38264
rect 28500 38224 28506 38236
rect 25958 38196 25964 38208
rect 24412 38168 25964 38196
rect 25958 38156 25964 38168
rect 26016 38196 26022 38208
rect 26234 38196 26240 38208
rect 26016 38168 26240 38196
rect 26016 38156 26022 38168
rect 26234 38156 26240 38168
rect 26292 38156 26298 38208
rect 26789 38199 26847 38205
rect 26789 38165 26801 38199
rect 26835 38196 26847 38199
rect 29546 38196 29552 38208
rect 26835 38168 29552 38196
rect 26835 38165 26847 38168
rect 26789 38159 26847 38165
rect 29546 38156 29552 38168
rect 29604 38156 29610 38208
rect 29730 38156 29736 38208
rect 29788 38196 29794 38208
rect 30101 38199 30159 38205
rect 30101 38196 30113 38199
rect 29788 38168 30113 38196
rect 29788 38156 29794 38168
rect 30101 38165 30113 38168
rect 30147 38165 30159 38199
rect 30101 38159 30159 38165
rect 31573 38199 31631 38205
rect 31573 38165 31585 38199
rect 31619 38196 31631 38199
rect 32950 38196 32956 38208
rect 31619 38168 32956 38196
rect 31619 38165 31631 38168
rect 31573 38159 31631 38165
rect 32950 38156 32956 38168
rect 33008 38156 33014 38208
rect 33060 38196 33088 38236
rect 33410 38224 33416 38276
rect 33468 38264 33474 38276
rect 33781 38267 33839 38273
rect 33781 38264 33793 38267
rect 33468 38236 33793 38264
rect 33468 38224 33474 38236
rect 33781 38233 33793 38236
rect 33827 38233 33839 38267
rect 33781 38227 33839 38233
rect 34882 38224 34888 38276
rect 34940 38224 34946 38276
rect 34992 38264 35020 38295
rect 35342 38264 35348 38276
rect 34992 38236 35348 38264
rect 35342 38224 35348 38236
rect 35400 38224 35406 38276
rect 36004 38264 36032 38304
rect 36078 38292 36084 38344
rect 36136 38332 36142 38344
rect 36136 38304 36181 38332
rect 36136 38292 36142 38304
rect 36262 38292 36268 38344
rect 36320 38332 36326 38344
rect 37093 38335 37151 38341
rect 37093 38332 37105 38335
rect 36320 38304 37105 38332
rect 36320 38292 36326 38304
rect 37093 38301 37105 38304
rect 37139 38332 37151 38335
rect 37921 38335 37979 38341
rect 37921 38332 37933 38335
rect 37139 38304 37933 38332
rect 37139 38301 37151 38304
rect 37093 38295 37151 38301
rect 37921 38301 37933 38304
rect 37967 38301 37979 38335
rect 38102 38332 38108 38344
rect 38063 38304 38108 38332
rect 37921 38295 37979 38301
rect 38102 38292 38108 38304
rect 38160 38292 38166 38344
rect 38194 38292 38200 38344
rect 38252 38332 38258 38344
rect 38746 38332 38752 38344
rect 38252 38304 38297 38332
rect 38707 38304 38752 38332
rect 38252 38292 38258 38304
rect 38746 38292 38752 38304
rect 38804 38292 38810 38344
rect 38930 38332 38936 38344
rect 38891 38304 38936 38332
rect 38930 38292 38936 38304
rect 38988 38292 38994 38344
rect 40586 38292 40592 38344
rect 40644 38332 40650 38344
rect 41601 38335 41659 38341
rect 40644 38304 41552 38332
rect 40644 38292 40650 38304
rect 36004 38236 36860 38264
rect 34790 38196 34796 38208
rect 33060 38168 34796 38196
rect 34790 38156 34796 38168
rect 34848 38156 34854 38208
rect 34974 38156 34980 38208
rect 35032 38196 35038 38208
rect 35713 38199 35771 38205
rect 35713 38196 35725 38199
rect 35032 38168 35725 38196
rect 35032 38156 35038 38168
rect 35713 38165 35725 38168
rect 35759 38165 35771 38199
rect 35713 38159 35771 38165
rect 35802 38156 35808 38208
rect 35860 38196 35866 38208
rect 36725 38199 36783 38205
rect 36725 38196 36737 38199
rect 35860 38168 36737 38196
rect 35860 38156 35866 38168
rect 36725 38165 36737 38168
rect 36771 38165 36783 38199
rect 36832 38196 36860 38236
rect 37826 38224 37832 38276
rect 37884 38264 37890 38276
rect 40957 38267 41015 38273
rect 40957 38264 40969 38267
rect 37884 38236 40969 38264
rect 37884 38224 37890 38236
rect 40957 38233 40969 38236
rect 41003 38233 41015 38267
rect 41524 38264 41552 38304
rect 41601 38301 41613 38335
rect 41647 38332 41659 38335
rect 42702 38332 42708 38344
rect 41647 38304 42708 38332
rect 41647 38301 41659 38304
rect 41601 38295 41659 38301
rect 42702 38292 42708 38304
rect 42760 38332 42766 38344
rect 43346 38332 43352 38344
rect 42760 38304 43352 38332
rect 42760 38292 42766 38304
rect 43346 38292 43352 38304
rect 43404 38332 43410 38344
rect 47397 38335 47455 38341
rect 47397 38332 47409 38335
rect 43404 38304 47409 38332
rect 43404 38292 43410 38304
rect 47397 38301 47409 38304
rect 47443 38332 47455 38335
rect 47857 38335 47915 38341
rect 47857 38332 47869 38335
rect 47443 38304 47869 38332
rect 47443 38301 47455 38304
rect 47397 38295 47455 38301
rect 47857 38301 47869 38304
rect 47903 38301 47915 38335
rect 47857 38295 47915 38301
rect 42150 38264 42156 38276
rect 41524 38236 42156 38264
rect 40957 38227 41015 38233
rect 42150 38224 42156 38236
rect 42208 38224 42214 38276
rect 39666 38196 39672 38208
rect 36832 38168 39672 38196
rect 36725 38159 36783 38165
rect 39666 38156 39672 38168
rect 39724 38156 39730 38208
rect 39850 38196 39856 38208
rect 39811 38168 39856 38196
rect 39850 38156 39856 38168
rect 39908 38156 39914 38208
rect 43162 38196 43168 38208
rect 43123 38168 43168 38196
rect 43162 38156 43168 38168
rect 43220 38156 43226 38208
rect 48038 38196 48044 38208
rect 47999 38168 48044 38196
rect 48038 38156 48044 38168
rect 48096 38156 48102 38208
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 1578 37992 1584 38004
rect 1539 37964 1584 37992
rect 1578 37952 1584 37964
rect 1636 37952 1642 38004
rect 12345 37995 12403 38001
rect 12345 37961 12357 37995
rect 12391 37992 12403 37995
rect 12434 37992 12440 38004
rect 12391 37964 12440 37992
rect 12391 37961 12403 37964
rect 12345 37955 12403 37961
rect 12434 37952 12440 37964
rect 12492 37992 12498 38004
rect 14182 37992 14188 38004
rect 12492 37964 14188 37992
rect 12492 37952 12498 37964
rect 14182 37952 14188 37964
rect 14240 37952 14246 38004
rect 16850 38001 16856 38004
rect 16846 37992 16856 38001
rect 16811 37964 16856 37992
rect 16846 37955 16856 37964
rect 16850 37952 16856 37955
rect 16908 37952 16914 38004
rect 17218 37952 17224 38004
rect 17276 37992 17282 38004
rect 17276 37964 18092 37992
rect 17276 37952 17282 37964
rect 13262 37884 13268 37936
rect 13320 37924 13326 37936
rect 13446 37924 13452 37936
rect 13320 37896 13452 37924
rect 13320 37884 13326 37896
rect 13446 37884 13452 37896
rect 13504 37884 13510 37936
rect 13538 37884 13544 37936
rect 13596 37924 13602 37936
rect 14550 37924 14556 37936
rect 13596 37896 14228 37924
rect 14511 37896 14556 37924
rect 13596 37884 13602 37896
rect 13906 37856 13912 37868
rect 13867 37828 13912 37856
rect 13906 37816 13912 37828
rect 13964 37816 13970 37868
rect 14200 37865 14228 37896
rect 14550 37884 14556 37896
rect 14608 37884 14614 37936
rect 16482 37884 16488 37936
rect 16540 37924 16546 37936
rect 16761 37927 16819 37933
rect 16761 37924 16773 37927
rect 16540 37896 16773 37924
rect 16540 37884 16546 37896
rect 16761 37893 16773 37896
rect 16807 37893 16819 37927
rect 18064 37924 18092 37964
rect 18138 37952 18144 38004
rect 18196 37992 18202 38004
rect 18693 37995 18751 38001
rect 18693 37992 18705 37995
rect 18196 37964 18705 37992
rect 18196 37952 18202 37964
rect 18693 37961 18705 37964
rect 18739 37961 18751 37995
rect 18693 37955 18751 37961
rect 21450 37952 21456 38004
rect 21508 37992 21514 38004
rect 22005 37995 22063 38001
rect 22005 37992 22017 37995
rect 21508 37964 22017 37992
rect 21508 37952 21514 37964
rect 22005 37961 22017 37964
rect 22051 37961 22063 37995
rect 22005 37955 22063 37961
rect 23198 37952 23204 38004
rect 23256 37992 23262 38004
rect 23385 37995 23443 38001
rect 23385 37992 23397 37995
rect 23256 37964 23397 37992
rect 23256 37952 23262 37964
rect 23385 37961 23397 37964
rect 23431 37961 23443 37995
rect 23385 37955 23443 37961
rect 23477 37995 23535 38001
rect 23477 37961 23489 37995
rect 23523 37992 23535 37995
rect 23842 37992 23848 38004
rect 23523 37964 23848 37992
rect 23523 37961 23535 37964
rect 23477 37955 23535 37961
rect 23842 37952 23848 37964
rect 23900 37952 23906 38004
rect 24394 37952 24400 38004
rect 24452 37992 24458 38004
rect 24857 37995 24915 38001
rect 24857 37992 24869 37995
rect 24452 37964 24869 37992
rect 24452 37952 24458 37964
rect 24857 37961 24869 37964
rect 24903 37961 24915 37995
rect 24857 37955 24915 37961
rect 25409 37995 25467 38001
rect 25409 37961 25421 37995
rect 25455 37992 25467 37995
rect 25682 37992 25688 38004
rect 25455 37964 25688 37992
rect 25455 37961 25467 37964
rect 25409 37955 25467 37961
rect 25682 37952 25688 37964
rect 25740 37952 25746 38004
rect 26421 37995 26479 38001
rect 26421 37961 26433 37995
rect 26467 37992 26479 37995
rect 29914 37992 29920 38004
rect 26467 37964 29920 37992
rect 26467 37961 26479 37964
rect 26421 37955 26479 37961
rect 29914 37952 29920 37964
rect 29972 37952 29978 38004
rect 30098 37992 30104 38004
rect 30059 37964 30104 37992
rect 30098 37952 30104 37964
rect 30156 37952 30162 38004
rect 30282 37952 30288 38004
rect 30340 37952 30346 38004
rect 33042 37992 33048 38004
rect 32416 37964 33048 37992
rect 23216 37924 23244 37952
rect 18064 37896 23244 37924
rect 16761 37887 16819 37893
rect 23290 37884 23296 37936
rect 23348 37924 23354 37936
rect 27154 37924 27160 37936
rect 23348 37896 26280 37924
rect 27115 37896 27160 37924
rect 23348 37884 23354 37896
rect 14093 37859 14151 37865
rect 14093 37825 14105 37859
rect 14139 37825 14151 37859
rect 14093 37819 14151 37825
rect 14185 37859 14243 37865
rect 14185 37825 14197 37859
rect 14231 37825 14243 37859
rect 14185 37819 14243 37825
rect 14108 37788 14136 37819
rect 14274 37816 14280 37868
rect 14332 37856 14338 37868
rect 15194 37856 15200 37868
rect 14332 37828 14377 37856
rect 15155 37828 15200 37856
rect 14332 37816 14338 37828
rect 15194 37816 15200 37828
rect 15252 37816 15258 37868
rect 15470 37856 15476 37868
rect 15431 37828 15476 37856
rect 15470 37816 15476 37828
rect 15528 37816 15534 37868
rect 16666 37856 16672 37868
rect 16627 37828 16672 37856
rect 16666 37816 16672 37828
rect 16724 37816 16730 37868
rect 16942 37856 16948 37868
rect 16903 37828 16948 37856
rect 16942 37816 16948 37828
rect 17000 37816 17006 37868
rect 17862 37856 17868 37868
rect 17823 37828 17868 37856
rect 17862 37816 17868 37828
rect 17920 37816 17926 37868
rect 18966 37856 18972 37868
rect 18879 37828 18972 37856
rect 18966 37816 18972 37828
rect 19024 37816 19030 37868
rect 20346 37856 20352 37868
rect 20307 37828 20352 37856
rect 20346 37816 20352 37828
rect 20404 37816 20410 37868
rect 22097 37859 22155 37865
rect 22097 37825 22109 37859
rect 22143 37856 22155 37859
rect 22281 37859 22339 37865
rect 22143 37828 22232 37856
rect 22143 37825 22155 37828
rect 22097 37819 22155 37825
rect 15286 37788 15292 37800
rect 14108 37760 15056 37788
rect 15247 37760 15292 37788
rect 12805 37723 12863 37729
rect 12805 37689 12817 37723
rect 12851 37720 12863 37723
rect 12894 37720 12900 37732
rect 12851 37692 12900 37720
rect 12851 37689 12863 37692
rect 12805 37683 12863 37689
rect 12894 37680 12900 37692
rect 12952 37720 12958 37732
rect 14918 37720 14924 37732
rect 12952 37692 14924 37720
rect 12952 37680 12958 37692
rect 14918 37680 14924 37692
rect 14976 37680 14982 37732
rect 15028 37729 15056 37760
rect 15286 37748 15292 37760
rect 15344 37748 15350 37800
rect 17678 37748 17684 37800
rect 17736 37788 17742 37800
rect 17773 37791 17831 37797
rect 17773 37788 17785 37791
rect 17736 37760 17785 37788
rect 17736 37748 17742 37760
rect 17773 37757 17785 37760
rect 17819 37757 17831 37791
rect 18690 37788 18696 37800
rect 18651 37760 18696 37788
rect 17773 37751 17831 37757
rect 15013 37723 15071 37729
rect 15013 37689 15025 37723
rect 15059 37689 15071 37723
rect 17218 37720 17224 37732
rect 15013 37683 15071 37689
rect 15120 37692 17224 37720
rect 10318 37612 10324 37664
rect 10376 37652 10382 37664
rect 10873 37655 10931 37661
rect 10873 37652 10885 37655
rect 10376 37624 10885 37652
rect 10376 37612 10382 37624
rect 10873 37621 10885 37624
rect 10919 37652 10931 37655
rect 11701 37655 11759 37661
rect 11701 37652 11713 37655
rect 10919 37624 11713 37652
rect 10919 37621 10931 37624
rect 10873 37615 10931 37621
rect 11701 37621 11713 37624
rect 11747 37621 11759 37655
rect 11701 37615 11759 37621
rect 13170 37612 13176 37664
rect 13228 37652 13234 37664
rect 15120 37652 15148 37692
rect 17218 37680 17224 37692
rect 17276 37680 17282 37732
rect 17788 37720 17816 37751
rect 18690 37748 18696 37760
rect 18748 37748 18754 37800
rect 18984 37788 19012 37816
rect 22204 37800 22232 37828
rect 22281 37825 22293 37859
rect 22327 37856 22339 37859
rect 22462 37856 22468 37868
rect 22327 37828 22468 37856
rect 22327 37825 22339 37828
rect 22281 37819 22339 37825
rect 22462 37816 22468 37828
rect 22520 37816 22526 37868
rect 23569 37859 23627 37865
rect 23569 37825 23581 37859
rect 23615 37856 23627 37859
rect 24026 37856 24032 37868
rect 23615 37828 24032 37856
rect 23615 37825 23627 37828
rect 23569 37819 23627 37825
rect 24026 37816 24032 37828
rect 24084 37816 24090 37868
rect 24210 37856 24216 37868
rect 24171 37828 24216 37856
rect 24210 37816 24216 37828
rect 24268 37816 24274 37868
rect 24486 37856 24492 37868
rect 24447 37828 24492 37856
rect 24486 37816 24492 37828
rect 24544 37816 24550 37868
rect 24670 37856 24676 37868
rect 24631 37828 24676 37856
rect 24670 37816 24676 37828
rect 24728 37816 24734 37868
rect 24854 37856 24860 37868
rect 24780 37828 24860 37856
rect 21726 37788 21732 37800
rect 18984 37760 21732 37788
rect 21726 37748 21732 37760
rect 21784 37748 21790 37800
rect 21818 37748 21824 37800
rect 21876 37788 21882 37800
rect 21876 37760 22094 37788
rect 21876 37748 21882 37760
rect 18138 37720 18144 37732
rect 17788 37692 18144 37720
rect 18138 37680 18144 37692
rect 18196 37680 18202 37732
rect 18230 37680 18236 37732
rect 18288 37720 18294 37732
rect 21634 37720 21640 37732
rect 18288 37692 18333 37720
rect 18892 37692 21640 37720
rect 18288 37680 18294 37692
rect 13228 37624 15148 37652
rect 15473 37655 15531 37661
rect 13228 37612 13234 37624
rect 15473 37621 15485 37655
rect 15519 37652 15531 37655
rect 15746 37652 15752 37664
rect 15519 37624 15752 37652
rect 15519 37621 15531 37624
rect 15473 37615 15531 37621
rect 15746 37612 15752 37624
rect 15804 37612 15810 37664
rect 16022 37652 16028 37664
rect 15983 37624 16028 37652
rect 16022 37612 16028 37624
rect 16080 37612 16086 37664
rect 16114 37612 16120 37664
rect 16172 37652 16178 37664
rect 18892 37661 18920 37692
rect 21634 37680 21640 37692
rect 21692 37680 21698 37732
rect 22066 37720 22094 37760
rect 22186 37748 22192 37800
rect 22244 37748 22250 37800
rect 23106 37748 23112 37800
rect 23164 37788 23170 37800
rect 23753 37791 23811 37797
rect 23753 37788 23765 37791
rect 23164 37760 23765 37788
rect 23164 37748 23170 37760
rect 23753 37757 23765 37760
rect 23799 37757 23811 37791
rect 23753 37751 23811 37757
rect 24394 37748 24400 37800
rect 24452 37788 24458 37800
rect 24578 37788 24584 37800
rect 24452 37760 24497 37788
rect 24539 37760 24584 37788
rect 24452 37748 24458 37760
rect 24578 37748 24584 37760
rect 24636 37748 24642 37800
rect 23201 37723 23259 37729
rect 23201 37720 23213 37723
rect 22066 37692 23213 37720
rect 23201 37689 23213 37692
rect 23247 37720 23259 37723
rect 24780 37720 24808 37828
rect 24854 37816 24860 37828
rect 24912 37816 24918 37868
rect 25958 37856 25964 37868
rect 25919 37828 25964 37856
rect 25958 37816 25964 37828
rect 26016 37816 26022 37868
rect 26252 37865 26280 37896
rect 27154 37884 27160 37896
rect 27212 37884 27218 37936
rect 28169 37927 28227 37933
rect 28169 37893 28181 37927
rect 28215 37893 28227 37927
rect 28169 37887 28227 37893
rect 28261 37927 28319 37933
rect 28261 37893 28273 37927
rect 28307 37893 28319 37927
rect 28261 37887 28319 37893
rect 26237 37859 26295 37865
rect 26237 37825 26249 37859
rect 26283 37825 26295 37859
rect 26237 37819 26295 37825
rect 26418 37816 26424 37868
rect 26476 37856 26482 37868
rect 27525 37859 27583 37865
rect 27525 37856 27537 37859
rect 26476 37828 27537 37856
rect 26476 37816 26482 37828
rect 27525 37825 27537 37828
rect 27571 37856 27583 37859
rect 27985 37859 28043 37865
rect 27985 37856 27997 37859
rect 27571 37828 27997 37856
rect 27571 37825 27583 37828
rect 27525 37819 27583 37825
rect 27985 37825 27997 37828
rect 28031 37825 28043 37859
rect 27985 37819 28043 37825
rect 26053 37791 26111 37797
rect 26053 37757 26065 37791
rect 26099 37788 26111 37791
rect 26099 37760 27016 37788
rect 26099 37757 26111 37760
rect 26053 37751 26111 37757
rect 23247 37692 24808 37720
rect 23247 37689 23259 37692
rect 23201 37683 23259 37689
rect 24854 37680 24860 37732
rect 24912 37720 24918 37732
rect 26988 37729 27016 37760
rect 26145 37723 26203 37729
rect 26145 37720 26157 37723
rect 24912 37692 26157 37720
rect 24912 37680 24918 37692
rect 26145 37689 26157 37692
rect 26191 37689 26203 37723
rect 26145 37683 26203 37689
rect 26973 37723 27031 37729
rect 26973 37689 26985 37723
rect 27019 37689 27031 37723
rect 28184 37720 28212 37887
rect 28276 37788 28304 37887
rect 28994 37884 29000 37936
rect 29052 37924 29058 37936
rect 30300 37924 30328 37952
rect 31021 37927 31079 37933
rect 31021 37924 31033 37927
rect 29052 37896 31033 37924
rect 29052 37884 29058 37896
rect 31021 37893 31033 37896
rect 31067 37893 31079 37927
rect 31021 37887 31079 37893
rect 28350 37816 28356 37868
rect 28408 37856 28414 37868
rect 28626 37856 28632 37868
rect 28408 37828 28632 37856
rect 28408 37816 28414 37828
rect 28626 37816 28632 37828
rect 28684 37816 28690 37868
rect 29365 37859 29423 37865
rect 29365 37825 29377 37859
rect 29411 37856 29423 37859
rect 29546 37856 29552 37868
rect 29411 37828 29552 37856
rect 29411 37825 29423 37828
rect 29365 37819 29423 37825
rect 29546 37816 29552 37828
rect 29604 37816 29610 37868
rect 30282 37856 30288 37868
rect 30243 37828 30288 37856
rect 30282 37816 30288 37828
rect 30340 37816 30346 37868
rect 30469 37859 30527 37865
rect 30469 37825 30481 37859
rect 30515 37856 30527 37859
rect 30558 37856 30564 37868
rect 30515 37828 30564 37856
rect 30515 37825 30527 37828
rect 30469 37819 30527 37825
rect 30558 37816 30564 37828
rect 30616 37856 30622 37868
rect 30742 37856 30748 37868
rect 30616 37828 30748 37856
rect 30616 37816 30622 37828
rect 30742 37816 30748 37828
rect 30800 37816 30806 37868
rect 30926 37856 30932 37868
rect 30887 37828 30932 37856
rect 30926 37816 30932 37828
rect 30984 37816 30990 37868
rect 31113 37859 31171 37865
rect 31113 37825 31125 37859
rect 31159 37856 31171 37859
rect 31294 37856 31300 37868
rect 31159 37828 31300 37856
rect 31159 37825 31171 37828
rect 31113 37819 31171 37825
rect 31294 37816 31300 37828
rect 31352 37816 31358 37868
rect 32030 37816 32036 37868
rect 32088 37856 32094 37868
rect 32416 37865 32444 37964
rect 33042 37952 33048 37964
rect 33100 37952 33106 38004
rect 33134 37952 33140 38004
rect 33192 37992 33198 38004
rect 33502 37992 33508 38004
rect 33192 37964 33508 37992
rect 33192 37952 33198 37964
rect 33502 37952 33508 37964
rect 33560 37952 33566 38004
rect 34882 37992 34888 38004
rect 34843 37964 34888 37992
rect 34882 37952 34888 37964
rect 34940 37952 34946 38004
rect 35710 37952 35716 38004
rect 35768 37992 35774 38004
rect 35989 37995 36047 38001
rect 35989 37992 36001 37995
rect 35768 37964 36001 37992
rect 35768 37952 35774 37964
rect 35989 37961 36001 37964
rect 36035 37961 36047 37995
rect 35989 37955 36047 37961
rect 37458 37952 37464 38004
rect 37516 37992 37522 38004
rect 38197 37995 38255 38001
rect 38197 37992 38209 37995
rect 37516 37964 38209 37992
rect 37516 37952 37522 37964
rect 38197 37961 38209 37964
rect 38243 37961 38255 37995
rect 38197 37955 38255 37961
rect 38378 37952 38384 38004
rect 38436 37952 38442 38004
rect 41046 37952 41052 38004
rect 41104 37992 41110 38004
rect 41141 37995 41199 38001
rect 41141 37992 41153 37995
rect 41104 37964 41153 37992
rect 41104 37952 41110 37964
rect 41141 37961 41153 37964
rect 41187 37961 41199 37995
rect 41690 37992 41696 38004
rect 41651 37964 41696 37992
rect 41141 37955 41199 37961
rect 41690 37952 41696 37964
rect 41748 37952 41754 38004
rect 42521 37995 42579 38001
rect 42521 37961 42533 37995
rect 42567 37992 42579 37995
rect 42978 37992 42984 38004
rect 42567 37964 42984 37992
rect 42567 37961 42579 37964
rect 42521 37955 42579 37961
rect 42978 37952 42984 37964
rect 43036 37952 43042 38004
rect 34330 37924 34336 37936
rect 32508 37896 34336 37924
rect 32508 37865 32536 37896
rect 34330 37884 34336 37896
rect 34388 37884 34394 37936
rect 35069 37927 35127 37933
rect 35069 37893 35081 37927
rect 35115 37924 35127 37927
rect 35526 37924 35532 37936
rect 35115 37896 35532 37924
rect 35115 37893 35127 37896
rect 35069 37887 35127 37893
rect 35526 37884 35532 37896
rect 35584 37884 35590 37936
rect 37369 37927 37427 37933
rect 37369 37924 37381 37927
rect 36188 37896 37381 37924
rect 36188 37868 36216 37896
rect 37369 37893 37381 37896
rect 37415 37893 37427 37927
rect 37369 37887 37427 37893
rect 38102 37884 38108 37936
rect 38160 37924 38166 37936
rect 38396 37924 38424 37952
rect 38160 37896 38424 37924
rect 38160 37884 38166 37896
rect 32401 37859 32459 37865
rect 32401 37856 32413 37859
rect 32088 37828 32413 37856
rect 32088 37816 32094 37828
rect 32401 37825 32413 37828
rect 32447 37825 32459 37859
rect 32401 37819 32459 37825
rect 32493 37859 32551 37865
rect 32493 37825 32505 37859
rect 32539 37825 32551 37859
rect 32493 37819 32551 37825
rect 32582 37816 32588 37868
rect 32640 37856 32646 37868
rect 32640 37828 32685 37856
rect 32640 37816 32646 37828
rect 32766 37816 32772 37868
rect 32824 37856 32830 37868
rect 32824 37828 32869 37856
rect 32824 37816 32830 37828
rect 33502 37816 33508 37868
rect 33560 37856 33566 37868
rect 33597 37859 33655 37865
rect 33597 37856 33609 37859
rect 33560 37828 33609 37856
rect 33560 37816 33566 37828
rect 33597 37825 33609 37828
rect 33643 37825 33655 37859
rect 33597 37819 33655 37825
rect 33781 37859 33839 37865
rect 33781 37825 33793 37859
rect 33827 37856 33839 37859
rect 34514 37856 34520 37868
rect 33827 37828 34520 37856
rect 33827 37825 33839 37828
rect 33781 37819 33839 37825
rect 34514 37816 34520 37828
rect 34572 37816 34578 37868
rect 35253 37859 35311 37865
rect 35253 37825 35265 37859
rect 35299 37825 35311 37859
rect 36170 37856 36176 37868
rect 36131 37828 36176 37856
rect 35253 37819 35311 37825
rect 28442 37788 28448 37800
rect 28276 37760 28448 37788
rect 28442 37748 28448 37760
rect 28500 37748 28506 37800
rect 30006 37748 30012 37800
rect 30064 37788 30070 37800
rect 32125 37791 32183 37797
rect 32125 37788 32137 37791
rect 30064 37760 32137 37788
rect 30064 37748 30070 37760
rect 32125 37757 32137 37760
rect 32171 37757 32183 37791
rect 35268 37788 35296 37819
rect 36170 37816 36176 37828
rect 36228 37816 36234 37868
rect 36262 37816 36268 37868
rect 36320 37856 36326 37868
rect 36449 37859 36507 37865
rect 36449 37856 36461 37859
rect 36320 37828 36461 37856
rect 36320 37816 36326 37828
rect 36449 37825 36461 37828
rect 36495 37825 36507 37859
rect 36449 37819 36507 37825
rect 37277 37859 37335 37865
rect 37277 37825 37289 37859
rect 37323 37825 37335 37859
rect 37458 37856 37464 37868
rect 37419 37828 37464 37856
rect 37277 37819 37335 37825
rect 35986 37788 35992 37800
rect 35268 37760 35992 37788
rect 32125 37751 32183 37757
rect 35986 37748 35992 37760
rect 36044 37788 36050 37800
rect 36538 37788 36544 37800
rect 36044 37760 36544 37788
rect 36044 37748 36050 37760
rect 36538 37748 36544 37760
rect 36596 37748 36602 37800
rect 37292 37788 37320 37819
rect 37458 37816 37464 37828
rect 37516 37816 37522 37868
rect 38565 37859 38623 37865
rect 38565 37825 38577 37859
rect 38611 37856 38623 37859
rect 39114 37856 39120 37868
rect 38611 37828 39120 37856
rect 38611 37825 38623 37828
rect 38565 37819 38623 37825
rect 39114 37816 39120 37828
rect 39172 37816 39178 37868
rect 40126 37816 40132 37868
rect 40184 37856 40190 37868
rect 40497 37859 40555 37865
rect 40497 37856 40509 37859
rect 40184 37828 40509 37856
rect 40184 37816 40190 37828
rect 40497 37825 40509 37828
rect 40543 37825 40555 37859
rect 40497 37819 40555 37825
rect 37550 37788 37556 37800
rect 37292 37760 37556 37788
rect 37550 37748 37556 37760
rect 37608 37748 37614 37800
rect 38470 37788 38476 37800
rect 38431 37760 38476 37788
rect 38470 37748 38476 37760
rect 38528 37748 38534 37800
rect 40589 37791 40647 37797
rect 40589 37757 40601 37791
rect 40635 37788 40647 37791
rect 41138 37788 41144 37800
rect 40635 37760 41144 37788
rect 40635 37757 40647 37760
rect 40589 37751 40647 37757
rect 41138 37748 41144 37760
rect 41196 37748 41202 37800
rect 28350 37720 28356 37732
rect 28184 37692 28356 37720
rect 26973 37683 27031 37689
rect 28350 37680 28356 37692
rect 28408 37680 28414 37732
rect 28537 37723 28595 37729
rect 28537 37689 28549 37723
rect 28583 37720 28595 37723
rect 29549 37723 29607 37729
rect 29549 37720 29561 37723
rect 28583 37692 29561 37720
rect 28583 37689 28595 37692
rect 28537 37683 28595 37689
rect 29549 37689 29561 37692
rect 29595 37720 29607 37723
rect 30190 37720 30196 37732
rect 29595 37692 30196 37720
rect 29595 37689 29607 37692
rect 29549 37683 29607 37689
rect 18877 37655 18935 37661
rect 18877 37652 18889 37655
rect 16172 37624 18889 37652
rect 16172 37612 16178 37624
rect 18877 37621 18889 37624
rect 18923 37621 18935 37655
rect 19886 37652 19892 37664
rect 19847 37624 19892 37652
rect 18877 37615 18935 37621
rect 19886 37612 19892 37624
rect 19944 37612 19950 37664
rect 20622 37652 20628 37664
rect 20583 37624 20628 37652
rect 20622 37612 20628 37624
rect 20680 37612 20686 37664
rect 20806 37652 20812 37664
rect 20767 37624 20812 37652
rect 20806 37612 20812 37624
rect 20864 37612 20870 37664
rect 21818 37652 21824 37664
rect 21779 37624 21824 37652
rect 21818 37612 21824 37624
rect 21876 37612 21882 37664
rect 22002 37612 22008 37664
rect 22060 37652 22066 37664
rect 24118 37652 24124 37664
rect 22060 37624 24124 37652
rect 22060 37612 22066 37624
rect 24118 37612 24124 37624
rect 24176 37652 24182 37664
rect 24394 37652 24400 37664
rect 24176 37624 24400 37652
rect 24176 37612 24182 37624
rect 24394 37612 24400 37624
rect 24452 37652 24458 37664
rect 25774 37652 25780 37664
rect 24452 37624 25780 37652
rect 24452 37612 24458 37624
rect 25774 37612 25780 37624
rect 25832 37612 25838 37664
rect 26050 37612 26056 37664
rect 26108 37652 26114 37664
rect 27157 37655 27215 37661
rect 27157 37652 27169 37655
rect 26108 37624 27169 37652
rect 26108 37612 26114 37624
rect 27157 37621 27169 37624
rect 27203 37621 27215 37655
rect 27157 37615 27215 37621
rect 28442 37612 28448 37664
rect 28500 37652 28506 37664
rect 28552 37652 28580 37683
rect 30190 37680 30196 37692
rect 30248 37680 30254 37732
rect 32674 37680 32680 37732
rect 32732 37720 32738 37732
rect 34054 37720 34060 37732
rect 32732 37692 34060 37720
rect 32732 37680 32738 37692
rect 34054 37680 34060 37692
rect 34112 37680 34118 37732
rect 36357 37723 36415 37729
rect 36357 37689 36369 37723
rect 36403 37720 36415 37723
rect 37366 37720 37372 37732
rect 36403 37692 37372 37720
rect 36403 37689 36415 37692
rect 36357 37683 36415 37689
rect 37366 37680 37372 37692
rect 37424 37680 37430 37732
rect 39206 37720 39212 37732
rect 39167 37692 39212 37720
rect 39206 37680 39212 37692
rect 39264 37680 39270 37732
rect 33594 37652 33600 37664
rect 28500 37624 28580 37652
rect 33555 37624 33600 37652
rect 28500 37612 28506 37624
rect 33594 37612 33600 37624
rect 33652 37612 33658 37664
rect 33686 37612 33692 37664
rect 33744 37652 33750 37664
rect 33965 37655 34023 37661
rect 33965 37652 33977 37655
rect 33744 37624 33977 37652
rect 33744 37612 33750 37624
rect 33965 37621 33977 37624
rect 34011 37621 34023 37655
rect 34072 37652 34100 37680
rect 37826 37652 37832 37664
rect 34072 37624 37832 37652
rect 33965 37615 34023 37621
rect 37826 37612 37832 37624
rect 37884 37612 37890 37664
rect 39022 37612 39028 37664
rect 39080 37652 39086 37664
rect 40129 37655 40187 37661
rect 40129 37652 40141 37655
rect 39080 37624 40141 37652
rect 39080 37612 39086 37624
rect 40129 37621 40141 37624
rect 40175 37621 40187 37655
rect 40129 37615 40187 37621
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 11517 37451 11575 37457
rect 11517 37417 11529 37451
rect 11563 37448 11575 37451
rect 11790 37448 11796 37460
rect 11563 37420 11796 37448
rect 11563 37417 11575 37420
rect 11517 37411 11575 37417
rect 11790 37408 11796 37420
rect 11848 37448 11854 37460
rect 13814 37448 13820 37460
rect 11848 37420 13820 37448
rect 11848 37408 11854 37420
rect 13814 37408 13820 37420
rect 13872 37448 13878 37460
rect 14369 37451 14427 37457
rect 13872 37420 14320 37448
rect 13872 37408 13878 37420
rect 10962 37380 10968 37392
rect 10875 37352 10968 37380
rect 10962 37340 10968 37352
rect 11020 37380 11026 37392
rect 12434 37380 12440 37392
rect 11020 37352 12440 37380
rect 11020 37340 11026 37352
rect 12434 37340 12440 37352
rect 12492 37340 12498 37392
rect 14292 37380 14320 37420
rect 14369 37417 14381 37451
rect 14415 37448 14427 37451
rect 15194 37448 15200 37460
rect 14415 37420 15200 37448
rect 14415 37417 14427 37420
rect 14369 37411 14427 37417
rect 15194 37408 15200 37420
rect 15252 37408 15258 37460
rect 16025 37451 16083 37457
rect 16025 37417 16037 37451
rect 16071 37448 16083 37451
rect 16482 37448 16488 37460
rect 16071 37420 16488 37448
rect 16071 37417 16083 37420
rect 16025 37411 16083 37417
rect 16482 37408 16488 37420
rect 16540 37408 16546 37460
rect 16942 37408 16948 37460
rect 17000 37408 17006 37460
rect 18046 37408 18052 37460
rect 18104 37448 18110 37460
rect 18601 37451 18659 37457
rect 18601 37448 18613 37451
rect 18104 37420 18613 37448
rect 18104 37408 18110 37420
rect 18601 37417 18613 37420
rect 18647 37448 18659 37451
rect 19150 37448 19156 37460
rect 18647 37420 19156 37448
rect 18647 37417 18659 37420
rect 18601 37411 18659 37417
rect 19150 37408 19156 37420
rect 19208 37408 19214 37460
rect 19613 37451 19671 37457
rect 19613 37417 19625 37451
rect 19659 37448 19671 37451
rect 20530 37448 20536 37460
rect 19659 37420 20536 37448
rect 19659 37417 19671 37420
rect 19613 37411 19671 37417
rect 20530 37408 20536 37420
rect 20588 37408 20594 37460
rect 20901 37451 20959 37457
rect 20901 37417 20913 37451
rect 20947 37448 20959 37451
rect 21818 37448 21824 37460
rect 20947 37420 21824 37448
rect 20947 37417 20959 37420
rect 20901 37411 20959 37417
rect 21818 37408 21824 37420
rect 21876 37408 21882 37460
rect 22094 37408 22100 37460
rect 22152 37448 22158 37460
rect 23934 37448 23940 37460
rect 22152 37420 23940 37448
rect 22152 37408 22158 37420
rect 23934 37408 23940 37420
rect 23992 37408 23998 37460
rect 24762 37408 24768 37460
rect 24820 37448 24826 37460
rect 24949 37451 25007 37457
rect 24949 37448 24961 37451
rect 24820 37420 24961 37448
rect 24820 37408 24826 37420
rect 24949 37417 24961 37420
rect 24995 37417 25007 37451
rect 25682 37448 25688 37460
rect 25643 37420 25688 37448
rect 24949 37411 25007 37417
rect 25682 37408 25688 37420
rect 25740 37408 25746 37460
rect 26237 37451 26295 37457
rect 26237 37417 26249 37451
rect 26283 37448 26295 37451
rect 26326 37448 26332 37460
rect 26283 37420 26332 37448
rect 26283 37417 26295 37420
rect 26237 37411 26295 37417
rect 14292 37352 14412 37380
rect 10318 37312 10324 37324
rect 10279 37284 10324 37312
rect 10318 37272 10324 37284
rect 10376 37312 10382 37324
rect 14384 37312 14412 37352
rect 16298 37340 16304 37392
rect 16356 37380 16362 37392
rect 16960 37380 16988 37408
rect 19058 37380 19064 37392
rect 16356 37352 19064 37380
rect 16356 37340 16362 37352
rect 19058 37340 19064 37352
rect 19116 37340 19122 37392
rect 20806 37380 20812 37392
rect 19536 37352 20812 37380
rect 10376 37284 12664 37312
rect 10376 37272 10382 37284
rect 12434 37204 12440 37256
rect 12492 37244 12498 37256
rect 12529 37247 12587 37253
rect 12529 37244 12541 37247
rect 12492 37216 12541 37244
rect 12492 37204 12498 37216
rect 12529 37213 12541 37216
rect 12575 37213 12587 37247
rect 12636 37244 12664 37284
rect 14384 37284 15056 37312
rect 12713 37247 12771 37253
rect 12713 37244 12725 37247
rect 12636 37216 12725 37244
rect 12529 37207 12587 37213
rect 12713 37213 12725 37216
rect 12759 37244 12771 37247
rect 13357 37247 13415 37253
rect 13357 37244 13369 37247
rect 12759 37216 13369 37244
rect 12759 37213 12771 37216
rect 12713 37207 12771 37213
rect 13357 37213 13369 37216
rect 13403 37244 13415 37247
rect 13446 37244 13452 37256
rect 13403 37216 13452 37244
rect 13403 37213 13415 37216
rect 13357 37207 13415 37213
rect 12544 37176 12572 37207
rect 13446 37204 13452 37216
rect 13504 37204 13510 37256
rect 14182 37244 14188 37256
rect 14143 37216 14188 37244
rect 14182 37204 14188 37216
rect 14240 37204 14246 37256
rect 14384 37253 14412 37284
rect 15028 37256 15056 37284
rect 16942 37272 16948 37324
rect 17000 37312 17006 37324
rect 18049 37315 18107 37321
rect 18049 37312 18061 37315
rect 17000 37284 18061 37312
rect 17000 37272 17006 37284
rect 18049 37281 18061 37284
rect 18095 37312 18107 37315
rect 18414 37312 18420 37324
rect 18095 37284 18420 37312
rect 18095 37281 18107 37284
rect 18049 37275 18107 37281
rect 18414 37272 18420 37284
rect 18472 37312 18478 37324
rect 19242 37312 19248 37324
rect 18472 37284 19248 37312
rect 18472 37272 18478 37284
rect 19242 37272 19248 37284
rect 19300 37272 19306 37324
rect 19536 37321 19564 37352
rect 20806 37340 20812 37352
rect 20864 37340 20870 37392
rect 21634 37380 21640 37392
rect 21595 37352 21640 37380
rect 21634 37340 21640 37352
rect 21692 37340 21698 37392
rect 23106 37340 23112 37392
rect 23164 37380 23170 37392
rect 23164 37352 23704 37380
rect 23164 37340 23170 37352
rect 19521 37315 19579 37321
rect 19521 37281 19533 37315
rect 19567 37281 19579 37315
rect 20346 37312 20352 37324
rect 19521 37275 19579 37281
rect 20272 37284 20352 37312
rect 14369 37247 14427 37253
rect 14369 37213 14381 37247
rect 14415 37213 14427 37247
rect 14369 37207 14427 37213
rect 14829 37247 14887 37253
rect 14829 37213 14841 37247
rect 14875 37213 14887 37247
rect 15010 37244 15016 37256
rect 14971 37216 15016 37244
rect 14829 37207 14887 37213
rect 13170 37176 13176 37188
rect 12544 37148 13176 37176
rect 13170 37136 13176 37148
rect 13228 37136 13234 37188
rect 13906 37176 13912 37188
rect 13464 37148 13912 37176
rect 12069 37111 12127 37117
rect 12069 37077 12081 37111
rect 12115 37108 12127 37111
rect 12526 37108 12532 37120
rect 12115 37080 12532 37108
rect 12115 37077 12127 37080
rect 12069 37071 12127 37077
rect 12526 37068 12532 37080
rect 12584 37068 12590 37120
rect 12713 37111 12771 37117
rect 12713 37077 12725 37111
rect 12759 37108 12771 37111
rect 13464 37108 13492 37148
rect 13906 37136 13912 37148
rect 13964 37136 13970 37188
rect 14200 37176 14228 37204
rect 14844 37176 14872 37207
rect 15010 37204 15016 37216
rect 15068 37204 15074 37256
rect 15197 37247 15255 37253
rect 15197 37213 15209 37247
rect 15243 37244 15255 37247
rect 15378 37244 15384 37256
rect 15243 37216 15384 37244
rect 15243 37213 15255 37216
rect 15197 37207 15255 37213
rect 15378 37204 15384 37216
rect 15436 37244 15442 37256
rect 15841 37247 15899 37253
rect 15841 37244 15853 37247
rect 15436 37216 15853 37244
rect 15436 37204 15442 37216
rect 15841 37213 15853 37216
rect 15887 37213 15899 37247
rect 15841 37207 15899 37213
rect 17313 37247 17371 37253
rect 17313 37213 17325 37247
rect 17359 37213 17371 37247
rect 17494 37244 17500 37256
rect 17455 37216 17500 37244
rect 17313 37207 17371 37213
rect 14200 37148 14872 37176
rect 15657 37179 15715 37185
rect 15657 37145 15669 37179
rect 15703 37145 15715 37179
rect 15657 37139 15715 37145
rect 12759 37080 13492 37108
rect 13541 37111 13599 37117
rect 12759 37077 12771 37080
rect 12713 37071 12771 37077
rect 13541 37077 13553 37111
rect 13587 37108 13599 37111
rect 14090 37108 14096 37120
rect 13587 37080 14096 37108
rect 13587 37077 13599 37080
rect 13541 37071 13599 37077
rect 14090 37068 14096 37080
rect 14148 37068 14154 37120
rect 15194 37068 15200 37120
rect 15252 37108 15258 37120
rect 15672 37108 15700 37139
rect 17218 37136 17224 37188
rect 17276 37176 17282 37188
rect 17328 37176 17356 37207
rect 17494 37204 17500 37216
rect 17552 37204 17558 37256
rect 18506 37204 18512 37256
rect 18564 37244 18570 37256
rect 20272 37253 20300 37284
rect 20346 37272 20352 37284
rect 20404 37272 20410 37324
rect 21542 37312 21548 37324
rect 21503 37284 21548 37312
rect 21542 37272 21548 37284
rect 21600 37272 21606 37324
rect 22094 37272 22100 37324
rect 22152 37312 22158 37324
rect 23201 37315 23259 37321
rect 23201 37312 23213 37315
rect 22152 37284 23213 37312
rect 22152 37272 22158 37284
rect 23201 37281 23213 37284
rect 23247 37312 23259 37315
rect 23382 37312 23388 37324
rect 23247 37284 23388 37312
rect 23247 37281 23259 37284
rect 23201 37275 23259 37281
rect 23382 37272 23388 37284
rect 23440 37272 23446 37324
rect 19429 37247 19487 37253
rect 19429 37244 19441 37247
rect 18564 37216 19441 37244
rect 18564 37204 18570 37216
rect 19429 37213 19441 37216
rect 19475 37213 19487 37247
rect 19429 37207 19487 37213
rect 20257 37247 20315 37253
rect 20257 37213 20269 37247
rect 20303 37213 20315 37247
rect 20441 37247 20499 37253
rect 20671 37247 20729 37253
rect 20441 37234 20453 37247
rect 20487 37234 20499 37247
rect 20552 37241 20610 37247
rect 20671 37244 20683 37247
rect 20552 37238 20564 37241
rect 20548 37234 20564 37238
rect 20257 37207 20315 37213
rect 18874 37176 18880 37188
rect 17276 37148 18880 37176
rect 17276 37136 17282 37148
rect 18874 37136 18880 37148
rect 18932 37136 18938 37188
rect 20438 37182 20444 37234
rect 20496 37182 20502 37234
rect 20530 37182 20536 37234
rect 20598 37207 20610 37241
rect 20588 37201 20610 37207
rect 20656 37213 20683 37244
rect 20717 37213 20729 37247
rect 21450 37244 21456 37256
rect 21411 37216 21456 37244
rect 20656 37207 20729 37213
rect 20588 37182 20594 37201
rect 20656 37176 20684 37207
rect 21450 37204 21456 37216
rect 21508 37204 21514 37256
rect 21726 37244 21732 37256
rect 21639 37216 21732 37244
rect 21726 37204 21732 37216
rect 21784 37204 21790 37256
rect 23014 37244 23020 37256
rect 22975 37216 23020 37244
rect 23014 37204 23020 37216
rect 23072 37204 23078 37256
rect 23676 37253 23704 37352
rect 23842 37340 23848 37392
rect 23900 37380 23906 37392
rect 24118 37380 24124 37392
rect 23900 37352 24124 37380
rect 23900 37340 23906 37352
rect 24118 37340 24124 37352
rect 24176 37340 24182 37392
rect 24302 37340 24308 37392
rect 24360 37380 24366 37392
rect 24360 37352 25084 37380
rect 24360 37340 24366 37352
rect 24486 37312 24492 37324
rect 24447 37284 24492 37312
rect 24486 37272 24492 37284
rect 24544 37272 24550 37324
rect 25056 37312 25084 37352
rect 25130 37340 25136 37392
rect 25188 37380 25194 37392
rect 25406 37380 25412 37392
rect 25188 37352 25412 37380
rect 25188 37340 25194 37352
rect 25406 37340 25412 37352
rect 25464 37380 25470 37392
rect 26252 37380 26280 37411
rect 26326 37408 26332 37420
rect 26384 37408 26390 37460
rect 27154 37408 27160 37460
rect 27212 37448 27218 37460
rect 27433 37451 27491 37457
rect 27433 37448 27445 37451
rect 27212 37420 27445 37448
rect 27212 37408 27218 37420
rect 27433 37417 27445 37420
rect 27479 37417 27491 37451
rect 27433 37411 27491 37417
rect 27985 37451 28043 37457
rect 27985 37417 27997 37451
rect 28031 37448 28043 37451
rect 28166 37448 28172 37460
rect 28031 37420 28172 37448
rect 28031 37417 28043 37420
rect 27985 37411 28043 37417
rect 28166 37408 28172 37420
rect 28224 37408 28230 37460
rect 28534 37408 28540 37460
rect 28592 37448 28598 37460
rect 32125 37451 32183 37457
rect 28592 37420 31754 37448
rect 28592 37408 28598 37420
rect 27798 37380 27804 37392
rect 25464 37352 26280 37380
rect 27172 37352 27804 37380
rect 25464 37340 25470 37352
rect 26050 37312 26056 37324
rect 24688 37284 24992 37312
rect 25056 37284 26056 37312
rect 23661 37247 23719 37253
rect 23661 37213 23673 37247
rect 23707 37213 23719 37247
rect 23842 37244 23848 37256
rect 23803 37216 23848 37244
rect 23661 37207 23719 37213
rect 23842 37204 23848 37216
rect 23900 37204 23906 37256
rect 24394 37244 24400 37256
rect 24355 37216 24400 37244
rect 24394 37204 24400 37216
rect 24452 37204 24458 37256
rect 24688 37253 24716 37284
rect 24673 37247 24731 37253
rect 24673 37213 24685 37247
rect 24719 37213 24731 37247
rect 24673 37207 24731 37213
rect 24765 37247 24823 37253
rect 24765 37213 24777 37247
rect 24811 37213 24823 37247
rect 24964 37244 24992 37284
rect 26050 37272 26056 37284
rect 26108 37272 26114 37324
rect 27062 37312 27068 37324
rect 27023 37284 27068 37312
rect 27062 37272 27068 37284
rect 27120 37272 27126 37324
rect 27172 37321 27200 37352
rect 27798 37340 27804 37352
rect 27856 37340 27862 37392
rect 28350 37340 28356 37392
rect 28408 37380 28414 37392
rect 28408 37352 28672 37380
rect 28408 37340 28414 37352
rect 27157 37315 27215 37321
rect 27157 37281 27169 37315
rect 27203 37281 27215 37315
rect 27157 37275 27215 37281
rect 27249 37315 27307 37321
rect 27249 37281 27261 37315
rect 27295 37312 27307 37315
rect 27706 37312 27712 37324
rect 27295 37284 27712 37312
rect 27295 37281 27307 37284
rect 27249 37275 27307 37281
rect 27706 37272 27712 37284
rect 27764 37312 27770 37324
rect 28368 37312 28396 37340
rect 27764 37284 28396 37312
rect 27764 37272 27770 37284
rect 25958 37244 25964 37256
rect 24964 37216 25964 37244
rect 24765 37207 24823 37213
rect 20640 37148 20684 37176
rect 21744 37176 21772 37204
rect 23753 37179 23811 37185
rect 21744 37148 23704 37176
rect 20640 37120 20668 37148
rect 15252 37080 15700 37108
rect 16853 37111 16911 37117
rect 15252 37068 15258 37080
rect 16853 37077 16865 37111
rect 16899 37108 16911 37111
rect 16942 37108 16948 37120
rect 16899 37080 16948 37108
rect 16899 37077 16911 37080
rect 16853 37071 16911 37077
rect 16942 37068 16948 37080
rect 17000 37068 17006 37120
rect 17497 37111 17555 37117
rect 17497 37077 17509 37111
rect 17543 37108 17555 37111
rect 17770 37108 17776 37120
rect 17543 37080 17776 37108
rect 17543 37077 17555 37080
rect 17497 37071 17555 37077
rect 17770 37068 17776 37080
rect 17828 37068 17834 37120
rect 19797 37111 19855 37117
rect 19797 37077 19809 37111
rect 19843 37108 19855 37111
rect 20162 37108 20168 37120
rect 19843 37080 20168 37108
rect 19843 37077 19855 37080
rect 19797 37071 19855 37077
rect 20162 37068 20168 37080
rect 20220 37068 20226 37120
rect 20622 37068 20628 37120
rect 20680 37068 20686 37120
rect 21913 37111 21971 37117
rect 21913 37077 21925 37111
rect 21959 37108 21971 37111
rect 22186 37108 22192 37120
rect 21959 37080 22192 37108
rect 21959 37077 21971 37080
rect 21913 37071 21971 37077
rect 22186 37068 22192 37080
rect 22244 37068 22250 37120
rect 22830 37108 22836 37120
rect 22791 37080 22836 37108
rect 22830 37068 22836 37080
rect 22888 37068 22894 37120
rect 23676 37108 23704 37148
rect 23753 37145 23765 37179
rect 23799 37176 23811 37179
rect 24780 37176 24808 37207
rect 25958 37204 25964 37216
rect 26016 37204 26022 37256
rect 26970 37244 26976 37256
rect 26931 37216 26976 37244
rect 26970 37204 26976 37216
rect 27028 37204 27034 37256
rect 27080 37244 27108 37272
rect 28644 37256 28672 37352
rect 30190 37340 30196 37392
rect 30248 37380 30254 37392
rect 31297 37383 31355 37389
rect 30248 37352 30325 37380
rect 30248 37340 30254 37352
rect 30098 37272 30104 37324
rect 30156 37312 30162 37324
rect 30156 37284 30236 37312
rect 30156 37272 30162 37284
rect 27982 37244 27988 37256
rect 27080 37216 27988 37244
rect 27982 37204 27988 37216
rect 28040 37244 28046 37256
rect 28442 37244 28448 37256
rect 28040 37216 28448 37244
rect 28040 37204 28046 37216
rect 28442 37204 28448 37216
rect 28500 37204 28506 37256
rect 28626 37244 28632 37256
rect 28587 37216 28632 37244
rect 28626 37204 28632 37216
rect 28684 37204 28690 37256
rect 28718 37204 28724 37256
rect 28776 37244 28782 37256
rect 30208 37253 30236 37284
rect 30297 37253 30325 37352
rect 31297 37349 31309 37383
rect 31343 37349 31355 37383
rect 31726 37380 31754 37420
rect 32125 37417 32137 37451
rect 32171 37448 32183 37451
rect 32582 37448 32588 37460
rect 32171 37420 32588 37448
rect 32171 37417 32183 37420
rect 32125 37411 32183 37417
rect 32582 37408 32588 37420
rect 32640 37408 32646 37460
rect 32861 37451 32919 37457
rect 32861 37417 32873 37451
rect 32907 37448 32919 37451
rect 33410 37448 33416 37460
rect 32907 37420 33416 37448
rect 32907 37417 32919 37420
rect 32861 37411 32919 37417
rect 32876 37380 32904 37411
rect 33410 37408 33416 37420
rect 33468 37408 33474 37460
rect 35342 37408 35348 37460
rect 35400 37448 35406 37460
rect 35805 37451 35863 37457
rect 35805 37448 35817 37451
rect 35400 37420 35817 37448
rect 35400 37408 35406 37420
rect 35805 37417 35817 37420
rect 35851 37448 35863 37451
rect 36630 37448 36636 37460
rect 35851 37420 36636 37448
rect 35851 37417 35863 37420
rect 35805 37411 35863 37417
rect 36630 37408 36636 37420
rect 36688 37408 36694 37460
rect 37918 37408 37924 37460
rect 37976 37448 37982 37460
rect 38473 37451 38531 37457
rect 38473 37448 38485 37451
rect 37976 37420 38485 37448
rect 37976 37408 37982 37420
rect 38473 37417 38485 37420
rect 38519 37448 38531 37451
rect 40586 37448 40592 37460
rect 38519 37420 40592 37448
rect 38519 37417 38531 37420
rect 38473 37411 38531 37417
rect 40586 37408 40592 37420
rect 40644 37408 40650 37460
rect 41138 37448 41144 37460
rect 41099 37420 41144 37448
rect 41138 37408 41144 37420
rect 41196 37408 41202 37460
rect 41693 37451 41751 37457
rect 41693 37417 41705 37451
rect 41739 37448 41751 37451
rect 42797 37451 42855 37457
rect 42797 37448 42809 37451
rect 41739 37420 42809 37448
rect 41739 37417 41751 37420
rect 41693 37411 41751 37417
rect 42797 37417 42809 37420
rect 42843 37448 42855 37451
rect 43346 37448 43352 37460
rect 42843 37420 43352 37448
rect 42843 37417 42855 37420
rect 42797 37411 42855 37417
rect 31726 37352 32904 37380
rect 33428 37380 33456 37408
rect 37366 37380 37372 37392
rect 33428 37352 36860 37380
rect 37327 37352 37372 37380
rect 31297 37343 31355 37349
rect 31018 37312 31024 37324
rect 30392 37284 31024 37312
rect 30392 37256 30420 37284
rect 31018 37272 31024 37284
rect 31076 37272 31082 37324
rect 31312 37312 31340 37343
rect 31754 37312 31760 37324
rect 31312 37284 31760 37312
rect 31754 37272 31760 37284
rect 31812 37272 31818 37324
rect 34054 37312 34060 37324
rect 31864 37284 34060 37312
rect 30193 37247 30251 37253
rect 28776 37216 30144 37244
rect 28776 37204 28782 37216
rect 29730 37176 29736 37188
rect 23799 37148 24808 37176
rect 24872 37148 29736 37176
rect 23799 37145 23811 37148
rect 23753 37139 23811 37145
rect 24872 37108 24900 37148
rect 29730 37136 29736 37148
rect 29788 37136 29794 37188
rect 30116 37176 30144 37216
rect 30193 37213 30205 37247
rect 30239 37213 30251 37247
rect 30193 37207 30251 37213
rect 30282 37247 30340 37253
rect 30282 37213 30294 37247
rect 30328 37213 30340 37247
rect 30282 37207 30340 37213
rect 30374 37204 30380 37256
rect 30432 37244 30438 37256
rect 30561 37247 30619 37253
rect 30432 37216 30477 37244
rect 30432 37204 30438 37216
rect 30561 37213 30573 37247
rect 30607 37244 30619 37247
rect 30742 37244 30748 37256
rect 30607 37216 30748 37244
rect 30607 37213 30619 37216
rect 30561 37207 30619 37213
rect 30742 37204 30748 37216
rect 30800 37204 30806 37256
rect 31205 37247 31263 37253
rect 31205 37213 31217 37247
rect 31251 37213 31263 37247
rect 31386 37244 31392 37256
rect 31347 37216 31392 37244
rect 31205 37207 31263 37213
rect 31220 37176 31248 37207
rect 31386 37204 31392 37216
rect 31444 37204 31450 37256
rect 31864 37176 31892 37284
rect 32030 37244 32036 37256
rect 31991 37216 32036 37244
rect 32030 37204 32036 37216
rect 32088 37204 32094 37256
rect 33520 37253 33548 37284
rect 34054 37272 34060 37284
rect 34112 37272 34118 37324
rect 34330 37272 34336 37324
rect 34388 37312 34394 37324
rect 36722 37312 36728 37324
rect 34388 37284 36728 37312
rect 34388 37272 34394 37284
rect 36722 37272 36728 37284
rect 36780 37272 36786 37324
rect 32217 37247 32275 37253
rect 32217 37213 32229 37247
rect 32263 37244 32275 37247
rect 33505 37247 33563 37253
rect 32263 37216 33180 37244
rect 32263 37213 32275 37216
rect 32217 37207 32275 37213
rect 30116 37148 31892 37176
rect 32490 37136 32496 37188
rect 32548 37176 32554 37188
rect 32677 37179 32735 37185
rect 32677 37176 32689 37179
rect 32548 37148 32689 37176
rect 32548 37136 32554 37148
rect 32677 37145 32689 37148
rect 32723 37145 32735 37179
rect 32677 37139 32735 37145
rect 32858 37136 32864 37188
rect 32916 37185 32922 37188
rect 32916 37179 32935 37185
rect 32923 37145 32935 37179
rect 33152 37176 33180 37216
rect 33505 37213 33517 37247
rect 33551 37213 33563 37247
rect 33686 37244 33692 37256
rect 33647 37216 33692 37244
rect 33505 37207 33563 37213
rect 33686 37204 33692 37216
rect 33744 37204 33750 37256
rect 33781 37247 33839 37253
rect 33781 37213 33793 37247
rect 33827 37213 33839 37247
rect 33781 37207 33839 37213
rect 33796 37176 33824 37207
rect 33870 37204 33876 37256
rect 33928 37244 33934 37256
rect 33928 37216 33973 37244
rect 33928 37204 33934 37216
rect 34238 37204 34244 37256
rect 34296 37244 34302 37256
rect 34701 37247 34759 37253
rect 34701 37244 34713 37247
rect 34296 37216 34713 37244
rect 34296 37204 34302 37216
rect 34701 37213 34713 37216
rect 34747 37213 34759 37247
rect 34701 37207 34759 37213
rect 35802 37204 35808 37256
rect 35860 37204 35866 37256
rect 36446 37244 36452 37256
rect 36407 37216 36452 37244
rect 36446 37204 36452 37216
rect 36504 37204 36510 37256
rect 36832 37253 36860 37352
rect 37366 37340 37372 37352
rect 37424 37340 37430 37392
rect 37829 37383 37887 37389
rect 37829 37349 37841 37383
rect 37875 37380 37887 37383
rect 38102 37380 38108 37392
rect 37875 37352 38108 37380
rect 37875 37349 37887 37352
rect 37829 37343 37887 37349
rect 38102 37340 38108 37352
rect 38160 37340 38166 37392
rect 41230 37380 41236 37392
rect 40972 37352 41236 37380
rect 37274 37272 37280 37324
rect 37332 37312 37338 37324
rect 40972 37321 41000 37352
rect 41230 37340 41236 37352
rect 41288 37340 41294 37392
rect 39209 37315 39267 37321
rect 39209 37312 39221 37315
rect 37332 37284 39221 37312
rect 37332 37272 37338 37284
rect 39209 37281 39221 37284
rect 39255 37281 39267 37315
rect 39209 37275 39267 37281
rect 40957 37315 41015 37321
rect 40957 37281 40969 37315
rect 41003 37281 41015 37315
rect 40957 37275 41015 37281
rect 36817 37247 36875 37253
rect 36817 37213 36829 37247
rect 36863 37244 36875 37247
rect 37458 37244 37464 37256
rect 36863 37216 37464 37244
rect 36863 37213 36875 37216
rect 36817 37207 36875 37213
rect 37458 37204 37464 37216
rect 37516 37244 37522 37256
rect 38562 37244 38568 37256
rect 37516 37216 38568 37244
rect 37516 37204 37522 37216
rect 38562 37204 38568 37216
rect 38620 37204 38626 37256
rect 39114 37244 39120 37256
rect 39075 37216 39120 37244
rect 39114 37204 39120 37216
rect 39172 37204 39178 37256
rect 39301 37247 39359 37253
rect 39301 37213 39313 37247
rect 39347 37213 39359 37247
rect 39301 37207 39359 37213
rect 34146 37176 34152 37188
rect 33152 37148 33824 37176
rect 34107 37148 34152 37176
rect 32916 37139 32935 37145
rect 32916 37136 32922 37139
rect 28534 37108 28540 37120
rect 23676 37080 24900 37108
rect 28495 37080 28540 37108
rect 28534 37068 28540 37080
rect 28592 37068 28598 37120
rect 29822 37068 29828 37120
rect 29880 37108 29886 37120
rect 29917 37111 29975 37117
rect 29917 37108 29929 37111
rect 29880 37080 29929 37108
rect 29880 37068 29886 37080
rect 29917 37077 29929 37080
rect 29963 37077 29975 37111
rect 29917 37071 29975 37077
rect 33045 37111 33103 37117
rect 33045 37077 33057 37111
rect 33091 37108 33103 37111
rect 33502 37108 33508 37120
rect 33091 37080 33508 37108
rect 33091 37077 33103 37080
rect 33045 37071 33103 37077
rect 33502 37068 33508 37080
rect 33560 37068 33566 37120
rect 33796 37108 33824 37148
rect 34146 37136 34152 37148
rect 34204 37136 34210 37188
rect 35820 37176 35848 37204
rect 34256 37148 35848 37176
rect 35989 37179 36047 37185
rect 34256 37108 34284 37148
rect 35989 37145 36001 37179
rect 36035 37176 36047 37179
rect 36262 37176 36268 37188
rect 36035 37148 36268 37176
rect 36035 37145 36047 37148
rect 35989 37139 36047 37145
rect 36262 37136 36268 37148
rect 36320 37136 36326 37188
rect 36633 37179 36691 37185
rect 36633 37145 36645 37179
rect 36679 37176 36691 37179
rect 37090 37176 37096 37188
rect 36679 37148 37096 37176
rect 36679 37145 36691 37148
rect 36633 37139 36691 37145
rect 37090 37136 37096 37148
rect 37148 37176 37154 37188
rect 37550 37176 37556 37188
rect 37148 37148 37556 37176
rect 37148 37136 37154 37148
rect 37550 37136 37556 37148
rect 37608 37136 37614 37188
rect 39316 37176 39344 37207
rect 39482 37204 39488 37256
rect 39540 37244 39546 37256
rect 39853 37247 39911 37253
rect 39853 37244 39865 37247
rect 39540 37216 39865 37244
rect 39540 37204 39546 37216
rect 39853 37213 39865 37216
rect 39899 37213 39911 37247
rect 39853 37207 39911 37213
rect 39942 37204 39948 37256
rect 40000 37244 40006 37256
rect 40037 37247 40095 37253
rect 40037 37244 40049 37247
rect 40000 37216 40049 37244
rect 40000 37204 40006 37216
rect 40037 37213 40049 37216
rect 40083 37244 40095 37247
rect 40083 37216 40724 37244
rect 40083 37213 40095 37216
rect 40037 37207 40095 37213
rect 40126 37176 40132 37188
rect 39316 37148 40132 37176
rect 40126 37136 40132 37148
rect 40184 37136 40190 37188
rect 40696 37176 40724 37216
rect 40770 37204 40776 37256
rect 40828 37246 40834 37256
rect 40865 37247 40923 37253
rect 40865 37246 40877 37247
rect 40828 37218 40877 37246
rect 40828 37204 40834 37218
rect 40865 37213 40877 37218
rect 40911 37213 40923 37247
rect 40865 37207 40923 37213
rect 41708 37176 41736 37411
rect 43346 37408 43352 37420
rect 43404 37408 43410 37460
rect 42150 37380 42156 37392
rect 42111 37352 42156 37380
rect 42150 37340 42156 37352
rect 42208 37340 42214 37392
rect 40696 37148 41736 37176
rect 33796 37080 34284 37108
rect 34698 37068 34704 37120
rect 34756 37108 34762 37120
rect 34793 37111 34851 37117
rect 34793 37108 34805 37111
rect 34756 37080 34805 37108
rect 34756 37068 34762 37080
rect 34793 37077 34805 37080
rect 34839 37077 34851 37111
rect 35618 37108 35624 37120
rect 35579 37080 35624 37108
rect 34793 37071 34851 37077
rect 35618 37068 35624 37080
rect 35676 37068 35682 37120
rect 35802 37117 35808 37120
rect 35789 37111 35808 37117
rect 35789 37077 35801 37111
rect 35789 37071 35808 37077
rect 35802 37068 35808 37071
rect 35860 37068 35866 37120
rect 40034 37108 40040 37120
rect 39995 37080 40040 37108
rect 40034 37068 40040 37080
rect 40092 37068 40098 37120
rect 40218 37068 40224 37120
rect 40276 37108 40282 37120
rect 40497 37111 40555 37117
rect 40497 37108 40509 37111
rect 40276 37080 40509 37108
rect 40276 37068 40282 37080
rect 40497 37077 40509 37080
rect 40543 37077 40555 37111
rect 40497 37071 40555 37077
rect 47762 37068 47768 37120
rect 47820 37108 47826 37120
rect 48041 37111 48099 37117
rect 48041 37108 48053 37111
rect 47820 37080 48053 37108
rect 47820 37068 47826 37080
rect 48041 37077 48053 37080
rect 48087 37077 48099 37111
rect 48041 37071 48099 37077
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 10962 36904 10968 36916
rect 10923 36876 10968 36904
rect 10962 36864 10968 36876
rect 11020 36864 11026 36916
rect 12434 36864 12440 36916
rect 12492 36904 12498 36916
rect 13538 36904 13544 36916
rect 12492 36876 12537 36904
rect 13499 36876 13544 36904
rect 12492 36864 12498 36876
rect 13538 36864 13544 36876
rect 13596 36864 13602 36916
rect 14277 36907 14335 36913
rect 14277 36873 14289 36907
rect 14323 36904 14335 36907
rect 14642 36904 14648 36916
rect 14323 36876 14648 36904
rect 14323 36873 14335 36876
rect 14277 36867 14335 36873
rect 14642 36864 14648 36876
rect 14700 36864 14706 36916
rect 16850 36904 16856 36916
rect 15212 36876 16856 36904
rect 11882 36836 11888 36848
rect 11795 36808 11888 36836
rect 11882 36796 11888 36808
rect 11940 36836 11946 36848
rect 11940 36808 12434 36836
rect 11940 36796 11946 36808
rect 12406 36700 12434 36808
rect 13170 36796 13176 36848
rect 13228 36836 13234 36848
rect 13228 36808 13676 36836
rect 13228 36796 13234 36808
rect 13446 36768 13452 36780
rect 13407 36740 13452 36768
rect 13446 36728 13452 36740
rect 13504 36728 13510 36780
rect 13538 36728 13544 36780
rect 13596 36768 13602 36780
rect 13648 36777 13676 36808
rect 13906 36796 13912 36848
rect 13964 36836 13970 36848
rect 15212 36836 15240 36876
rect 16850 36864 16856 36876
rect 16908 36864 16914 36916
rect 19061 36907 19119 36913
rect 19061 36873 19073 36907
rect 19107 36904 19119 36907
rect 20530 36904 20536 36916
rect 19107 36876 20536 36904
rect 19107 36873 19119 36876
rect 19061 36867 19119 36873
rect 20530 36864 20536 36876
rect 20588 36864 20594 36916
rect 20714 36904 20720 36916
rect 20675 36876 20720 36904
rect 20714 36864 20720 36876
rect 20772 36864 20778 36916
rect 22094 36904 22100 36916
rect 21192 36876 22100 36904
rect 15378 36836 15384 36848
rect 13964 36808 14320 36836
rect 13964 36796 13970 36808
rect 13633 36771 13691 36777
rect 13633 36768 13645 36771
rect 13596 36740 13645 36768
rect 13596 36728 13602 36740
rect 13633 36737 13645 36740
rect 13679 36737 13691 36771
rect 14090 36768 14096 36780
rect 14051 36740 14096 36768
rect 13633 36731 13691 36737
rect 14090 36728 14096 36740
rect 14148 36728 14154 36780
rect 14292 36777 14320 36808
rect 14384 36808 15240 36836
rect 15339 36808 15384 36836
rect 14277 36771 14335 36777
rect 14277 36737 14289 36771
rect 14323 36737 14335 36771
rect 14277 36731 14335 36737
rect 14384 36700 14412 36808
rect 15378 36796 15384 36808
rect 15436 36796 15442 36848
rect 17954 36836 17960 36848
rect 17420 36808 17960 36836
rect 15102 36768 15108 36780
rect 15063 36740 15108 36768
rect 15102 36728 15108 36740
rect 15160 36728 15166 36780
rect 17420 36777 17448 36808
rect 17954 36796 17960 36808
rect 18012 36796 18018 36848
rect 18690 36836 18696 36848
rect 18248 36808 18696 36836
rect 15197 36771 15255 36777
rect 15197 36737 15209 36771
rect 15243 36737 15255 36771
rect 15197 36731 15255 36737
rect 17405 36771 17463 36777
rect 17405 36737 17417 36771
rect 17451 36737 17463 36771
rect 17405 36731 17463 36737
rect 17497 36771 17555 36777
rect 17497 36737 17509 36771
rect 17543 36737 17555 36771
rect 17497 36731 17555 36737
rect 17681 36771 17739 36777
rect 17681 36737 17693 36771
rect 17727 36768 17739 36771
rect 18248 36768 18276 36808
rect 18690 36796 18696 36808
rect 18748 36796 18754 36848
rect 19797 36839 19855 36845
rect 19797 36805 19809 36839
rect 19843 36836 19855 36839
rect 20622 36836 20628 36848
rect 19843 36808 20628 36836
rect 19843 36805 19855 36808
rect 19797 36799 19855 36805
rect 20622 36796 20628 36808
rect 20680 36796 20686 36848
rect 17727 36740 18276 36768
rect 18325 36771 18383 36777
rect 17727 36737 17739 36740
rect 17681 36731 17739 36737
rect 18325 36737 18337 36771
rect 18371 36737 18383 36771
rect 18506 36768 18512 36780
rect 18467 36740 18512 36768
rect 18325 36731 18383 36737
rect 15212 36700 15240 36731
rect 12406 36672 14412 36700
rect 15120 36672 15240 36700
rect 17512 36700 17540 36731
rect 18340 36700 18368 36731
rect 18506 36728 18512 36740
rect 18564 36728 18570 36780
rect 18598 36728 18604 36780
rect 18656 36768 18662 36780
rect 18874 36768 18880 36780
rect 18656 36740 18701 36768
rect 18835 36740 18880 36768
rect 18656 36728 18662 36740
rect 18874 36728 18880 36740
rect 18932 36728 18938 36780
rect 19334 36728 19340 36780
rect 19392 36728 19398 36780
rect 19702 36768 19708 36780
rect 19663 36740 19708 36768
rect 19702 36728 19708 36740
rect 19760 36728 19766 36780
rect 19886 36768 19892 36780
rect 19847 36740 19892 36768
rect 19886 36728 19892 36740
rect 19944 36728 19950 36780
rect 20349 36771 20407 36777
rect 20349 36737 20361 36771
rect 20395 36737 20407 36771
rect 20530 36768 20536 36780
rect 20491 36740 20536 36768
rect 20349 36731 20407 36737
rect 18690 36700 18696 36712
rect 17512 36672 18460 36700
rect 18651 36672 18696 36700
rect 12526 36592 12532 36644
rect 12584 36632 12590 36644
rect 15120 36632 15148 36672
rect 12584 36604 15148 36632
rect 12584 36592 12590 36604
rect 15286 36592 15292 36644
rect 15344 36632 15350 36644
rect 15381 36635 15439 36641
rect 15381 36632 15393 36635
rect 15344 36604 15393 36632
rect 15344 36592 15350 36604
rect 15381 36601 15393 36604
rect 15427 36601 15439 36635
rect 18432 36632 18460 36672
rect 18690 36660 18696 36672
rect 18748 36660 18754 36712
rect 19352 36700 19380 36728
rect 20364 36700 20392 36731
rect 20530 36728 20536 36740
rect 20588 36728 20594 36780
rect 20622 36700 20628 36712
rect 19352 36672 20628 36700
rect 20622 36660 20628 36672
rect 20680 36700 20686 36712
rect 21192 36709 21220 36876
rect 22094 36864 22100 36876
rect 22152 36864 22158 36916
rect 22646 36864 22652 36916
rect 22704 36904 22710 36916
rect 22925 36907 22983 36913
rect 22925 36904 22937 36907
rect 22704 36876 22937 36904
rect 22704 36864 22710 36876
rect 22925 36873 22937 36876
rect 22971 36873 22983 36907
rect 22925 36867 22983 36873
rect 23842 36864 23848 36916
rect 23900 36904 23906 36916
rect 24397 36907 24455 36913
rect 24397 36904 24409 36907
rect 23900 36876 24409 36904
rect 23900 36864 23906 36876
rect 24397 36873 24409 36876
rect 24443 36873 24455 36907
rect 24397 36867 24455 36873
rect 24670 36864 24676 36916
rect 24728 36904 24734 36916
rect 26053 36907 26111 36913
rect 26053 36904 26065 36907
rect 24728 36876 26065 36904
rect 24728 36864 24734 36876
rect 26053 36873 26065 36876
rect 26099 36904 26111 36907
rect 26234 36904 26240 36916
rect 26099 36876 26240 36904
rect 26099 36873 26111 36876
rect 26053 36867 26111 36873
rect 26234 36864 26240 36876
rect 26292 36864 26298 36916
rect 28258 36904 28264 36916
rect 28219 36876 28264 36904
rect 28258 36864 28264 36876
rect 28316 36864 28322 36916
rect 28626 36864 28632 36916
rect 28684 36904 28690 36916
rect 33042 36904 33048 36916
rect 28684 36876 33048 36904
rect 28684 36864 28690 36876
rect 33042 36864 33048 36876
rect 33100 36904 33106 36916
rect 33597 36907 33655 36913
rect 33597 36904 33609 36907
rect 33100 36876 33609 36904
rect 33100 36864 33106 36876
rect 33597 36873 33609 36876
rect 33643 36873 33655 36907
rect 33597 36867 33655 36873
rect 35713 36907 35771 36913
rect 35713 36873 35725 36907
rect 35759 36904 35771 36907
rect 37274 36904 37280 36916
rect 35759 36876 37280 36904
rect 35759 36873 35771 36876
rect 35713 36867 35771 36873
rect 37274 36864 37280 36876
rect 37332 36864 37338 36916
rect 38102 36864 38108 36916
rect 38160 36904 38166 36916
rect 40218 36904 40224 36916
rect 38160 36876 40080 36904
rect 40179 36876 40224 36904
rect 38160 36864 38166 36876
rect 22462 36836 22468 36848
rect 21284 36808 22468 36836
rect 21177 36703 21235 36709
rect 21177 36700 21189 36703
rect 20680 36672 21189 36700
rect 20680 36660 20686 36672
rect 21177 36669 21189 36672
rect 21223 36669 21235 36703
rect 21177 36663 21235 36669
rect 19334 36632 19340 36644
rect 18432 36604 19340 36632
rect 15381 36595 15439 36601
rect 19334 36592 19340 36604
rect 19392 36592 19398 36644
rect 19702 36592 19708 36644
rect 19760 36632 19766 36644
rect 20254 36632 20260 36644
rect 19760 36604 20260 36632
rect 19760 36592 19766 36604
rect 20254 36592 20260 36604
rect 20312 36592 20318 36644
rect 20530 36592 20536 36644
rect 20588 36632 20594 36644
rect 21284 36632 21312 36808
rect 22462 36796 22468 36808
rect 22520 36796 22526 36848
rect 23661 36839 23719 36845
rect 23661 36836 23673 36839
rect 22664 36808 23673 36836
rect 22664 36777 22692 36808
rect 23661 36805 23673 36808
rect 23707 36805 23719 36839
rect 23661 36799 23719 36805
rect 23934 36796 23940 36848
rect 23992 36836 23998 36848
rect 24762 36836 24768 36848
rect 23992 36808 24768 36836
rect 23992 36796 23998 36808
rect 24762 36796 24768 36808
rect 24820 36796 24826 36848
rect 25130 36836 25136 36848
rect 25091 36808 25136 36836
rect 25130 36796 25136 36808
rect 25188 36796 25194 36848
rect 25222 36796 25228 36848
rect 25280 36836 25286 36848
rect 25333 36839 25391 36845
rect 25333 36836 25345 36839
rect 25280 36808 25345 36836
rect 25280 36796 25286 36808
rect 25333 36805 25345 36808
rect 25379 36805 25391 36839
rect 25333 36799 25391 36805
rect 25866 36796 25872 36848
rect 25924 36836 25930 36848
rect 29822 36836 29828 36848
rect 25924 36808 28764 36836
rect 29783 36808 29828 36836
rect 25924 36796 25930 36808
rect 28736 36780 28764 36808
rect 29822 36796 29828 36808
rect 29880 36796 29886 36848
rect 31110 36796 31116 36848
rect 31168 36836 31174 36848
rect 32766 36836 32772 36848
rect 31168 36808 32352 36836
rect 32727 36808 32772 36836
rect 31168 36796 31174 36808
rect 22649 36771 22707 36777
rect 22649 36737 22661 36771
rect 22695 36737 22707 36771
rect 23382 36768 23388 36780
rect 23343 36740 23388 36768
rect 22649 36731 22707 36737
rect 23382 36728 23388 36740
rect 23440 36728 23446 36780
rect 24118 36728 24124 36780
rect 24176 36768 24182 36780
rect 24305 36771 24363 36777
rect 24305 36768 24317 36771
rect 24176 36740 24317 36768
rect 24176 36728 24182 36740
rect 24305 36737 24317 36740
rect 24351 36737 24363 36771
rect 24305 36731 24363 36737
rect 24489 36771 24547 36777
rect 24489 36737 24501 36771
rect 24535 36768 24547 36771
rect 24578 36768 24584 36780
rect 24535 36740 24584 36768
rect 24535 36737 24547 36740
rect 24489 36731 24547 36737
rect 24578 36728 24584 36740
rect 24636 36728 24642 36780
rect 27433 36771 27491 36777
rect 27433 36737 27445 36771
rect 27479 36768 27491 36771
rect 27798 36768 27804 36780
rect 27479 36740 27804 36768
rect 27479 36737 27491 36740
rect 27433 36731 27491 36737
rect 27798 36728 27804 36740
rect 27856 36728 27862 36780
rect 28442 36768 28448 36780
rect 28403 36740 28448 36768
rect 28442 36728 28448 36740
rect 28500 36728 28506 36780
rect 28534 36728 28540 36780
rect 28592 36768 28598 36780
rect 28629 36771 28687 36777
rect 28629 36768 28641 36771
rect 28592 36740 28641 36768
rect 28592 36728 28598 36740
rect 28629 36737 28641 36740
rect 28675 36737 28687 36771
rect 28629 36731 28687 36737
rect 28718 36728 28724 36780
rect 28776 36768 28782 36780
rect 28905 36771 28963 36777
rect 28776 36740 28869 36768
rect 28776 36728 28782 36740
rect 28905 36737 28917 36771
rect 28951 36737 28963 36771
rect 29546 36768 29552 36780
rect 29507 36740 29552 36768
rect 28905 36731 28963 36737
rect 22278 36700 22284 36712
rect 22239 36672 22284 36700
rect 22278 36660 22284 36672
rect 22336 36660 22342 36712
rect 22370 36660 22376 36712
rect 22428 36700 22434 36712
rect 22741 36703 22799 36709
rect 22428 36672 22473 36700
rect 22428 36660 22434 36672
rect 22741 36669 22753 36703
rect 22787 36700 22799 36703
rect 22830 36700 22836 36712
rect 22787 36672 22836 36700
rect 22787 36669 22799 36672
rect 22741 36663 22799 36669
rect 22830 36660 22836 36672
rect 22888 36660 22894 36712
rect 23014 36660 23020 36712
rect 23072 36700 23078 36712
rect 23477 36703 23535 36709
rect 23477 36700 23489 36703
rect 23072 36672 23489 36700
rect 23072 36660 23078 36672
rect 23477 36669 23489 36672
rect 23523 36669 23535 36703
rect 23477 36663 23535 36669
rect 23566 36660 23572 36712
rect 23624 36700 23630 36712
rect 23661 36703 23719 36709
rect 23661 36700 23673 36703
rect 23624 36672 23673 36700
rect 23624 36660 23630 36672
rect 23661 36669 23673 36672
rect 23707 36669 23719 36703
rect 23661 36663 23719 36669
rect 27341 36703 27399 36709
rect 27341 36669 27353 36703
rect 27387 36700 27399 36703
rect 27522 36700 27528 36712
rect 27387 36672 27528 36700
rect 27387 36669 27399 36672
rect 27341 36663 27399 36669
rect 20588 36604 21312 36632
rect 23676 36632 23704 36663
rect 27522 36660 27528 36672
rect 27580 36700 27586 36712
rect 28920 36700 28948 36731
rect 29546 36728 29552 36740
rect 29604 36728 29610 36780
rect 29641 36771 29699 36777
rect 29641 36737 29653 36771
rect 29687 36768 29699 36771
rect 30098 36768 30104 36780
rect 29687 36740 30104 36768
rect 29687 36737 29699 36740
rect 29641 36731 29699 36737
rect 30098 36728 30104 36740
rect 30156 36728 30162 36780
rect 30374 36768 30380 36780
rect 30335 36740 30380 36768
rect 30374 36728 30380 36740
rect 30432 36728 30438 36780
rect 30558 36768 30564 36780
rect 30519 36740 30564 36768
rect 30558 36728 30564 36740
rect 30616 36728 30622 36780
rect 31205 36771 31263 36777
rect 31205 36737 31217 36771
rect 31251 36737 31263 36771
rect 31205 36731 31263 36737
rect 31110 36700 31116 36712
rect 27580 36672 28580 36700
rect 28920 36672 31116 36700
rect 27580 36660 27586 36672
rect 25130 36632 25136 36644
rect 23676 36604 25136 36632
rect 20588 36592 20594 36604
rect 25130 36592 25136 36604
rect 25188 36592 25194 36644
rect 25501 36635 25559 36641
rect 25501 36601 25513 36635
rect 25547 36632 25559 36635
rect 26142 36632 26148 36644
rect 25547 36604 26148 36632
rect 25547 36601 25559 36604
rect 25501 36595 25559 36601
rect 26142 36592 26148 36604
rect 26200 36592 26206 36644
rect 28442 36632 28448 36644
rect 27724 36604 28448 36632
rect 12989 36567 13047 36573
rect 12989 36533 13001 36567
rect 13035 36564 13047 36567
rect 15838 36564 15844 36576
rect 13035 36536 15844 36564
rect 13035 36533 13047 36536
rect 12989 36527 13047 36533
rect 15838 36524 15844 36536
rect 15896 36524 15902 36576
rect 16114 36564 16120 36576
rect 16075 36536 16120 36564
rect 16114 36524 16120 36536
rect 16172 36524 16178 36576
rect 16942 36564 16948 36576
rect 16903 36536 16948 36564
rect 16942 36524 16948 36536
rect 17000 36524 17006 36576
rect 17865 36567 17923 36573
rect 17865 36533 17877 36567
rect 17911 36564 17923 36567
rect 20070 36564 20076 36576
rect 17911 36536 20076 36564
rect 17911 36533 17923 36536
rect 17865 36527 17923 36533
rect 20070 36524 20076 36536
rect 20128 36524 20134 36576
rect 25314 36564 25320 36576
rect 25227 36536 25320 36564
rect 25314 36524 25320 36536
rect 25372 36564 25378 36576
rect 25682 36564 25688 36576
rect 25372 36536 25688 36564
rect 25372 36524 25378 36536
rect 25682 36524 25688 36536
rect 25740 36524 25746 36576
rect 25958 36524 25964 36576
rect 26016 36564 26022 36576
rect 27724 36564 27752 36604
rect 28442 36592 28448 36604
rect 28500 36592 28506 36644
rect 28552 36641 28580 36672
rect 31110 36660 31116 36672
rect 31168 36660 31174 36712
rect 31220 36700 31248 36731
rect 31294 36728 31300 36780
rect 31352 36768 31358 36780
rect 32324 36768 32352 36808
rect 32766 36796 32772 36808
rect 32824 36796 32830 36848
rect 33502 36796 33508 36848
rect 33560 36836 33566 36848
rect 33749 36839 33807 36845
rect 33749 36836 33761 36839
rect 33560 36808 33761 36836
rect 33560 36796 33566 36808
rect 33749 36805 33761 36808
rect 33795 36805 33807 36839
rect 33749 36799 33807 36805
rect 33965 36839 34023 36845
rect 33965 36805 33977 36839
rect 34011 36805 34023 36839
rect 33965 36799 34023 36805
rect 32490 36768 32496 36780
rect 31352 36740 31397 36768
rect 32324 36740 32496 36768
rect 31352 36728 31358 36740
rect 32490 36728 32496 36740
rect 32548 36728 32554 36780
rect 32641 36771 32699 36777
rect 32641 36737 32653 36771
rect 32687 36768 32699 36771
rect 32858 36771 32916 36777
rect 32687 36737 32720 36768
rect 32641 36731 32720 36737
rect 32858 36737 32870 36771
rect 32904 36737 32916 36771
rect 32858 36731 32916 36737
rect 31478 36700 31484 36712
rect 31220 36672 31484 36700
rect 31478 36660 31484 36672
rect 31536 36660 31542 36712
rect 32306 36660 32312 36712
rect 32364 36700 32370 36712
rect 32692 36700 32720 36731
rect 32364 36672 32720 36700
rect 32364 36660 32370 36672
rect 28537 36635 28595 36641
rect 28537 36601 28549 36635
rect 28583 36601 28595 36635
rect 28537 36595 28595 36601
rect 29638 36592 29644 36644
rect 29696 36632 29702 36644
rect 29825 36635 29883 36641
rect 29825 36632 29837 36635
rect 29696 36604 29837 36632
rect 29696 36592 29702 36604
rect 29825 36601 29837 36604
rect 29871 36601 29883 36635
rect 29825 36595 29883 36601
rect 30392 36604 30696 36632
rect 26016 36536 27752 36564
rect 27801 36567 27859 36573
rect 26016 36524 26022 36536
rect 27801 36533 27813 36567
rect 27847 36564 27859 36567
rect 28166 36564 28172 36576
rect 27847 36536 28172 36564
rect 27847 36533 27859 36536
rect 27801 36527 27859 36533
rect 28166 36524 28172 36536
rect 28224 36524 28230 36576
rect 28994 36524 29000 36576
rect 29052 36564 29058 36576
rect 30392 36564 30420 36604
rect 30558 36564 30564 36576
rect 29052 36536 30420 36564
rect 30519 36536 30564 36564
rect 29052 36524 29058 36536
rect 30558 36524 30564 36536
rect 30616 36524 30622 36576
rect 30668 36564 30696 36604
rect 32398 36592 32404 36644
rect 32456 36632 32462 36644
rect 32876 36632 32904 36731
rect 32950 36728 32956 36780
rect 33008 36777 33014 36780
rect 33008 36768 33016 36777
rect 33008 36740 33053 36768
rect 33008 36731 33016 36740
rect 33008 36728 33014 36731
rect 33594 36728 33600 36780
rect 33652 36768 33658 36780
rect 33980 36768 34008 36799
rect 35526 36796 35532 36848
rect 35584 36836 35590 36848
rect 36081 36839 36139 36845
rect 36081 36836 36093 36839
rect 35584 36808 36093 36836
rect 35584 36796 35590 36808
rect 36081 36805 36093 36808
rect 36127 36836 36139 36839
rect 38289 36839 38347 36845
rect 36127 36808 36768 36836
rect 36127 36805 36139 36808
rect 36081 36799 36139 36805
rect 34514 36768 34520 36780
rect 33652 36740 34008 36768
rect 34475 36740 34520 36768
rect 33652 36728 33658 36740
rect 34514 36728 34520 36740
rect 34572 36728 34578 36780
rect 34793 36771 34851 36777
rect 34793 36737 34805 36771
rect 34839 36768 34851 36771
rect 35434 36768 35440 36780
rect 34839 36740 35440 36768
rect 34839 36737 34851 36740
rect 34793 36731 34851 36737
rect 32456 36604 32904 36632
rect 34517 36635 34575 36641
rect 32456 36592 32462 36604
rect 34517 36601 34529 36635
rect 34563 36632 34575 36635
rect 34698 36632 34704 36644
rect 34563 36604 34704 36632
rect 34563 36601 34575 36604
rect 34517 36595 34575 36601
rect 34698 36592 34704 36604
rect 34756 36592 34762 36644
rect 31294 36564 31300 36576
rect 30668 36536 31300 36564
rect 31294 36524 31300 36536
rect 31352 36524 31358 36576
rect 31938 36524 31944 36576
rect 31996 36564 32002 36576
rect 32490 36564 32496 36576
rect 31996 36536 32496 36564
rect 31996 36524 32002 36536
rect 32490 36524 32496 36536
rect 32548 36524 32554 36576
rect 33137 36567 33195 36573
rect 33137 36533 33149 36567
rect 33183 36564 33195 36567
rect 33318 36564 33324 36576
rect 33183 36536 33324 36564
rect 33183 36533 33195 36536
rect 33137 36527 33195 36533
rect 33318 36524 33324 36536
rect 33376 36524 33382 36576
rect 33781 36567 33839 36573
rect 33781 36533 33793 36567
rect 33827 36564 33839 36567
rect 33870 36564 33876 36576
rect 33827 36536 33876 36564
rect 33827 36533 33839 36536
rect 33781 36527 33839 36533
rect 33870 36524 33876 36536
rect 33928 36524 33934 36576
rect 34238 36524 34244 36576
rect 34296 36564 34302 36576
rect 34422 36564 34428 36576
rect 34296 36536 34428 36564
rect 34296 36524 34302 36536
rect 34422 36524 34428 36536
rect 34480 36564 34486 36576
rect 34808 36564 34836 36731
rect 35434 36728 35440 36740
rect 35492 36728 35498 36780
rect 35802 36768 35808 36780
rect 35763 36740 35808 36768
rect 35802 36728 35808 36740
rect 35860 36728 35866 36780
rect 35897 36771 35955 36777
rect 35897 36737 35909 36771
rect 35943 36768 35955 36771
rect 35986 36768 35992 36780
rect 35943 36740 35992 36768
rect 35943 36737 35955 36740
rect 35897 36731 35955 36737
rect 35986 36728 35992 36740
rect 36044 36768 36050 36780
rect 36740 36777 36768 36808
rect 38289 36805 38301 36839
rect 38335 36836 38347 36839
rect 38470 36836 38476 36848
rect 38335 36808 38476 36836
rect 38335 36805 38347 36808
rect 38289 36799 38347 36805
rect 38470 36796 38476 36808
rect 38528 36836 38534 36848
rect 40052 36836 40080 36876
rect 40218 36864 40224 36876
rect 40276 36864 40282 36916
rect 42521 36907 42579 36913
rect 42521 36873 42533 36907
rect 42567 36904 42579 36907
rect 42610 36904 42616 36916
rect 42567 36876 42616 36904
rect 42567 36873 42579 36876
rect 42521 36867 42579 36873
rect 42610 36864 42616 36876
rect 42668 36864 42674 36916
rect 43073 36907 43131 36913
rect 43073 36873 43085 36907
rect 43119 36904 43131 36907
rect 43346 36904 43352 36916
rect 43119 36876 43352 36904
rect 43119 36873 43131 36876
rect 43073 36867 43131 36873
rect 43346 36864 43352 36876
rect 43404 36864 43410 36916
rect 40402 36836 40408 36848
rect 38528 36808 39804 36836
rect 40052 36808 40408 36836
rect 38528 36796 38534 36808
rect 36541 36771 36599 36777
rect 36541 36768 36553 36771
rect 36044 36740 36553 36768
rect 36044 36728 36050 36740
rect 36541 36737 36553 36740
rect 36587 36737 36599 36771
rect 36541 36731 36599 36737
rect 36725 36771 36783 36777
rect 36725 36737 36737 36771
rect 36771 36737 36783 36771
rect 36725 36731 36783 36737
rect 37921 36771 37979 36777
rect 37921 36737 37933 36771
rect 37967 36737 37979 36771
rect 38378 36768 38384 36780
rect 38339 36740 38384 36768
rect 37921 36731 37979 36737
rect 36630 36700 36636 36712
rect 36591 36672 36636 36700
rect 36630 36660 36636 36672
rect 36688 36700 36694 36712
rect 37936 36700 37964 36731
rect 38378 36728 38384 36740
rect 38436 36728 38442 36780
rect 38562 36728 38568 36780
rect 38620 36768 38626 36780
rect 39117 36771 39175 36777
rect 39117 36768 39129 36771
rect 38620 36740 39129 36768
rect 38620 36728 38626 36740
rect 39117 36737 39129 36740
rect 39163 36737 39175 36771
rect 39117 36731 39175 36737
rect 39301 36771 39359 36777
rect 39301 36737 39313 36771
rect 39347 36768 39359 36771
rect 39482 36768 39488 36780
rect 39347 36740 39488 36768
rect 39347 36737 39359 36740
rect 39301 36731 39359 36737
rect 36688 36672 37964 36700
rect 39132 36700 39160 36731
rect 39482 36728 39488 36740
rect 39540 36728 39546 36780
rect 39776 36777 39804 36808
rect 40402 36796 40408 36808
rect 40460 36796 40466 36848
rect 40862 36796 40868 36848
rect 40920 36836 40926 36848
rect 40920 36808 41460 36836
rect 40920 36796 40926 36808
rect 39761 36771 39819 36777
rect 39761 36737 39773 36771
rect 39807 36737 39819 36771
rect 41230 36768 41236 36780
rect 41191 36740 41236 36768
rect 39761 36731 39819 36737
rect 41230 36728 41236 36740
rect 41288 36728 41294 36780
rect 41432 36777 41460 36808
rect 44174 36796 44180 36848
rect 44232 36836 44238 36848
rect 46661 36839 46719 36845
rect 46661 36836 46673 36839
rect 44232 36808 46673 36836
rect 44232 36796 44238 36808
rect 46661 36805 46673 36808
rect 46707 36805 46719 36839
rect 47578 36836 47584 36848
rect 47539 36808 47584 36836
rect 46661 36799 46719 36805
rect 47578 36796 47584 36808
rect 47636 36796 47642 36848
rect 41417 36771 41475 36777
rect 41417 36737 41429 36771
rect 41463 36737 41475 36771
rect 41417 36731 41475 36737
rect 46845 36771 46903 36777
rect 46845 36737 46857 36771
rect 46891 36768 46903 36771
rect 47762 36768 47768 36780
rect 46891 36740 47624 36768
rect 47723 36740 47768 36768
rect 46891 36737 46903 36740
rect 46845 36731 46903 36737
rect 39942 36700 39948 36712
rect 39132 36672 39948 36700
rect 36688 36660 36694 36672
rect 39942 36660 39948 36672
rect 40000 36660 40006 36712
rect 40773 36703 40831 36709
rect 40773 36700 40785 36703
rect 40512 36672 40785 36700
rect 37274 36632 37280 36644
rect 37235 36604 37280 36632
rect 37274 36592 37280 36604
rect 37332 36592 37338 36644
rect 38059 36635 38117 36641
rect 38059 36601 38071 36635
rect 38105 36632 38117 36635
rect 38654 36632 38660 36644
rect 38105 36604 38660 36632
rect 38105 36601 38117 36604
rect 38059 36595 38117 36601
rect 38654 36592 38660 36604
rect 38712 36592 38718 36644
rect 39301 36635 39359 36641
rect 39301 36601 39313 36635
rect 39347 36632 39359 36635
rect 40310 36632 40316 36644
rect 39347 36604 40316 36632
rect 39347 36601 39359 36604
rect 39301 36595 39359 36601
rect 40310 36592 40316 36604
rect 40368 36592 40374 36644
rect 34480 36536 34836 36564
rect 34480 36524 34486 36536
rect 35342 36524 35348 36576
rect 35400 36564 35406 36576
rect 35529 36567 35587 36573
rect 35529 36564 35541 36567
rect 35400 36536 35541 36564
rect 35400 36524 35406 36536
rect 35529 36533 35541 36536
rect 35575 36533 35587 36567
rect 38194 36564 38200 36576
rect 38155 36536 38200 36564
rect 35529 36527 35587 36533
rect 38194 36524 38200 36536
rect 38252 36524 38258 36576
rect 39114 36524 39120 36576
rect 39172 36564 39178 36576
rect 39850 36564 39856 36576
rect 39172 36536 39856 36564
rect 39172 36524 39178 36536
rect 39850 36524 39856 36536
rect 39908 36564 39914 36576
rect 40512 36564 40540 36672
rect 40773 36669 40785 36672
rect 40819 36669 40831 36703
rect 40773 36663 40831 36669
rect 47029 36703 47087 36709
rect 47029 36669 47041 36703
rect 47075 36669 47087 36703
rect 47596 36700 47624 36740
rect 47762 36728 47768 36740
rect 47820 36728 47826 36780
rect 47946 36768 47952 36780
rect 47907 36740 47952 36768
rect 47946 36728 47952 36740
rect 48004 36728 48010 36780
rect 47964 36700 47992 36728
rect 47596 36672 47992 36700
rect 47029 36663 47087 36669
rect 47044 36632 47072 36663
rect 47210 36632 47216 36644
rect 47044 36604 47216 36632
rect 47210 36592 47216 36604
rect 47268 36632 47274 36644
rect 47762 36632 47768 36644
rect 47268 36604 47768 36632
rect 47268 36592 47274 36604
rect 47762 36592 47768 36604
rect 47820 36592 47826 36644
rect 39908 36536 40540 36564
rect 39908 36524 39914 36536
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 11882 36360 11888 36372
rect 11843 36332 11888 36360
rect 11882 36320 11888 36332
rect 11940 36320 11946 36372
rect 15930 36360 15936 36372
rect 15891 36332 15936 36360
rect 15930 36320 15936 36332
rect 15988 36320 15994 36372
rect 18230 36360 18236 36372
rect 18191 36332 18236 36360
rect 18230 36320 18236 36332
rect 18288 36320 18294 36372
rect 18506 36320 18512 36372
rect 18564 36360 18570 36372
rect 18601 36363 18659 36369
rect 18601 36360 18613 36363
rect 18564 36332 18613 36360
rect 18564 36320 18570 36332
rect 18601 36329 18613 36332
rect 18647 36329 18659 36363
rect 19334 36360 19340 36372
rect 19295 36332 19340 36360
rect 18601 36323 18659 36329
rect 19334 36320 19340 36332
rect 19392 36320 19398 36372
rect 20438 36320 20444 36372
rect 20496 36360 20502 36372
rect 20533 36363 20591 36369
rect 20533 36360 20545 36363
rect 20496 36332 20545 36360
rect 20496 36320 20502 36332
rect 20533 36329 20545 36332
rect 20579 36329 20591 36363
rect 20533 36323 20591 36329
rect 22738 36320 22744 36372
rect 22796 36360 22802 36372
rect 25406 36360 25412 36372
rect 22796 36332 25412 36360
rect 22796 36320 22802 36332
rect 25406 36320 25412 36332
rect 25464 36320 25470 36372
rect 26786 36320 26792 36372
rect 26844 36360 26850 36372
rect 26973 36363 27031 36369
rect 26973 36360 26985 36363
rect 26844 36332 26985 36360
rect 26844 36320 26850 36332
rect 26973 36329 26985 36332
rect 27019 36329 27031 36363
rect 27522 36360 27528 36372
rect 27483 36332 27528 36360
rect 26973 36323 27031 36329
rect 27522 36320 27528 36332
rect 27580 36320 27586 36372
rect 27614 36320 27620 36372
rect 27672 36360 27678 36372
rect 28353 36363 28411 36369
rect 28353 36360 28365 36363
rect 27672 36332 28365 36360
rect 27672 36320 27678 36332
rect 28353 36329 28365 36332
rect 28399 36329 28411 36363
rect 28353 36323 28411 36329
rect 30374 36320 30380 36372
rect 30432 36360 30438 36372
rect 30834 36360 30840 36372
rect 30432 36332 30840 36360
rect 30432 36320 30438 36332
rect 30834 36320 30840 36332
rect 30892 36320 30898 36372
rect 31386 36320 31392 36372
rect 31444 36360 31450 36372
rect 31849 36363 31907 36369
rect 31849 36360 31861 36363
rect 31444 36332 31861 36360
rect 31444 36320 31450 36332
rect 31849 36329 31861 36332
rect 31895 36329 31907 36363
rect 31849 36323 31907 36329
rect 32766 36320 32772 36372
rect 32824 36360 32830 36372
rect 32861 36363 32919 36369
rect 32861 36360 32873 36363
rect 32824 36332 32873 36360
rect 32824 36320 32830 36332
rect 32861 36329 32873 36332
rect 32907 36329 32919 36363
rect 32861 36323 32919 36329
rect 34606 36320 34612 36372
rect 34664 36360 34670 36372
rect 35253 36363 35311 36369
rect 35253 36360 35265 36363
rect 34664 36332 35265 36360
rect 34664 36320 34670 36332
rect 35253 36329 35265 36332
rect 35299 36329 35311 36363
rect 35618 36360 35624 36372
rect 35579 36332 35624 36360
rect 35253 36323 35311 36329
rect 35618 36320 35624 36332
rect 35676 36320 35682 36372
rect 38197 36363 38255 36369
rect 38197 36329 38209 36363
rect 38243 36360 38255 36363
rect 38378 36360 38384 36372
rect 38243 36332 38384 36360
rect 38243 36329 38255 36332
rect 38197 36323 38255 36329
rect 38378 36320 38384 36332
rect 38436 36360 38442 36372
rect 38436 36332 40172 36360
rect 38436 36320 38442 36332
rect 2225 36295 2283 36301
rect 2225 36261 2237 36295
rect 2271 36292 2283 36295
rect 21726 36292 21732 36304
rect 2271 36264 21732 36292
rect 2271 36261 2283 36264
rect 2225 36255 2283 36261
rect 1673 36159 1731 36165
rect 1673 36125 1685 36159
rect 1719 36156 1731 36159
rect 2240 36156 2268 36255
rect 21726 36252 21732 36264
rect 21784 36292 21790 36304
rect 25317 36295 25375 36301
rect 21784 36264 22140 36292
rect 21784 36252 21790 36264
rect 15562 36224 15568 36236
rect 15523 36196 15568 36224
rect 15562 36184 15568 36196
rect 15620 36184 15626 36236
rect 16577 36227 16635 36233
rect 16577 36193 16589 36227
rect 16623 36224 16635 36227
rect 17218 36224 17224 36236
rect 16623 36196 17224 36224
rect 16623 36193 16635 36196
rect 16577 36187 16635 36193
rect 17218 36184 17224 36196
rect 17276 36184 17282 36236
rect 17770 36184 17776 36236
rect 17828 36224 17834 36236
rect 18325 36227 18383 36233
rect 18325 36224 18337 36227
rect 17828 36196 18337 36224
rect 17828 36184 17834 36196
rect 18325 36193 18337 36196
rect 18371 36193 18383 36227
rect 19978 36224 19984 36236
rect 18325 36187 18383 36193
rect 19260 36196 19984 36224
rect 12986 36156 12992 36168
rect 1719 36128 2268 36156
rect 12899 36128 12992 36156
rect 1719 36125 1731 36128
rect 1673 36119 1731 36125
rect 12986 36116 12992 36128
rect 13044 36156 13050 36168
rect 15654 36156 15660 36168
rect 13044 36128 14412 36156
rect 15615 36128 15660 36156
rect 13044 36116 13050 36128
rect 11333 36091 11391 36097
rect 11333 36057 11345 36091
rect 11379 36088 11391 36091
rect 11882 36088 11888 36100
rect 11379 36060 11888 36088
rect 11379 36057 11391 36060
rect 11333 36051 11391 36057
rect 11882 36048 11888 36060
rect 11940 36048 11946 36100
rect 12437 36091 12495 36097
rect 12437 36057 12449 36091
rect 12483 36088 12495 36091
rect 14090 36088 14096 36100
rect 12483 36060 14096 36088
rect 12483 36057 12495 36060
rect 12437 36051 12495 36057
rect 14090 36048 14096 36060
rect 14148 36048 14154 36100
rect 1486 36020 1492 36032
rect 1447 35992 1492 36020
rect 1486 35980 1492 35992
rect 1544 35980 1550 36032
rect 13541 36023 13599 36029
rect 13541 35989 13553 36023
rect 13587 36020 13599 36023
rect 13722 36020 13728 36032
rect 13587 35992 13728 36020
rect 13587 35989 13599 35992
rect 13541 35983 13599 35989
rect 13722 35980 13728 35992
rect 13780 35980 13786 36032
rect 14384 36020 14412 36128
rect 15654 36116 15660 36128
rect 15712 36116 15718 36168
rect 16485 36159 16543 36165
rect 16485 36125 16497 36159
rect 16531 36156 16543 36159
rect 16669 36159 16727 36165
rect 16531 36128 16620 36156
rect 16531 36125 16543 36128
rect 16485 36119 16543 36125
rect 16592 36100 16620 36128
rect 16669 36125 16681 36159
rect 16715 36156 16727 36159
rect 16850 36156 16856 36168
rect 16715 36128 16856 36156
rect 16715 36125 16727 36128
rect 16669 36119 16727 36125
rect 16850 36116 16856 36128
rect 16908 36116 16914 36168
rect 17494 36116 17500 36168
rect 17552 36156 17558 36168
rect 17589 36159 17647 36165
rect 17589 36156 17601 36159
rect 17552 36128 17601 36156
rect 17552 36116 17558 36128
rect 17589 36125 17601 36128
rect 17635 36125 17647 36159
rect 17589 36119 17647 36125
rect 17678 36116 17684 36168
rect 17736 36156 17742 36168
rect 19260 36165 19288 36196
rect 19978 36184 19984 36196
rect 20036 36224 20042 36236
rect 21450 36224 21456 36236
rect 20036 36196 21456 36224
rect 20036 36184 20042 36196
rect 21450 36184 21456 36196
rect 21508 36184 21514 36236
rect 18233 36159 18291 36165
rect 17736 36128 17781 36156
rect 17736 36116 17742 36128
rect 18233 36125 18245 36159
rect 18279 36125 18291 36159
rect 18233 36119 18291 36125
rect 19245 36159 19303 36165
rect 19245 36125 19257 36159
rect 19291 36125 19303 36159
rect 19426 36156 19432 36168
rect 19387 36128 19432 36156
rect 19245 36119 19303 36125
rect 14461 36091 14519 36097
rect 14461 36057 14473 36091
rect 14507 36088 14519 36091
rect 16022 36088 16028 36100
rect 14507 36060 16028 36088
rect 14507 36057 14519 36060
rect 14461 36051 14519 36057
rect 16022 36048 16028 36060
rect 16080 36048 16086 36100
rect 16574 36048 16580 36100
rect 16632 36048 16638 36100
rect 18248 36088 18276 36119
rect 19426 36116 19432 36128
rect 19484 36116 19490 36168
rect 20438 36156 20444 36168
rect 20399 36128 20444 36156
rect 20438 36116 20444 36128
rect 20496 36116 20502 36168
rect 20622 36156 20628 36168
rect 20583 36128 20628 36156
rect 20622 36116 20628 36128
rect 20680 36116 20686 36168
rect 22112 36165 22140 36264
rect 25317 36261 25329 36295
rect 25363 36261 25375 36295
rect 25317 36255 25375 36261
rect 22830 36224 22836 36236
rect 22743 36196 22836 36224
rect 22830 36184 22836 36196
rect 22888 36184 22894 36236
rect 22097 36159 22155 36165
rect 22097 36125 22109 36159
rect 22143 36156 22155 36159
rect 22738 36156 22744 36168
rect 22143 36128 22600 36156
rect 22699 36128 22744 36156
rect 22143 36125 22155 36128
rect 22097 36119 22155 36125
rect 18322 36088 18328 36100
rect 18248 36060 18328 36088
rect 18322 36048 18328 36060
rect 18380 36088 18386 36100
rect 18690 36088 18696 36100
rect 18380 36060 18696 36088
rect 18380 36048 18386 36060
rect 18690 36048 18696 36060
rect 18748 36048 18754 36100
rect 19981 36091 20039 36097
rect 19981 36057 19993 36091
rect 20027 36088 20039 36091
rect 22572 36088 22600 36128
rect 22738 36116 22744 36128
rect 22796 36116 22802 36168
rect 22848 36156 22876 36184
rect 25041 36159 25099 36165
rect 25041 36156 25053 36159
rect 22848 36128 25053 36156
rect 25041 36125 25053 36128
rect 25087 36156 25099 36159
rect 25222 36156 25228 36168
rect 25087 36128 25228 36156
rect 25087 36125 25099 36128
rect 25041 36119 25099 36125
rect 25222 36116 25228 36128
rect 25280 36116 25286 36168
rect 25332 36156 25360 36255
rect 28626 36252 28632 36304
rect 28684 36292 28690 36304
rect 28813 36295 28871 36301
rect 28813 36292 28825 36295
rect 28684 36264 28825 36292
rect 28684 36252 28690 36264
rect 28813 36261 28825 36264
rect 28859 36261 28871 36295
rect 28813 36255 28871 36261
rect 28902 36252 28908 36304
rect 28960 36292 28966 36304
rect 28960 36264 30328 36292
rect 28960 36252 28966 36264
rect 28442 36184 28448 36236
rect 28500 36224 28506 36236
rect 30300 36224 30328 36264
rect 31294 36252 31300 36304
rect 31352 36292 31358 36304
rect 36081 36295 36139 36301
rect 31352 36264 35572 36292
rect 31352 36252 31358 36264
rect 31846 36224 31852 36236
rect 28500 36196 28672 36224
rect 28500 36184 28506 36196
rect 25777 36159 25835 36165
rect 25777 36156 25789 36159
rect 25332 36128 25789 36156
rect 25777 36125 25789 36128
rect 25823 36125 25835 36159
rect 25777 36119 25835 36125
rect 25961 36159 26019 36165
rect 25961 36125 25973 36159
rect 26007 36156 26019 36159
rect 26142 36156 26148 36168
rect 26007 36128 26148 36156
rect 26007 36125 26019 36128
rect 25961 36119 26019 36125
rect 26142 36116 26148 36128
rect 26200 36116 26206 36168
rect 27706 36156 27712 36168
rect 27667 36128 27712 36156
rect 27706 36116 27712 36128
rect 27764 36116 27770 36168
rect 27893 36159 27951 36165
rect 27893 36125 27905 36159
rect 27939 36156 27951 36159
rect 27982 36156 27988 36168
rect 27939 36128 27988 36156
rect 27939 36125 27951 36128
rect 27893 36119 27951 36125
rect 27982 36116 27988 36128
rect 28040 36116 28046 36168
rect 28166 36116 28172 36168
rect 28224 36156 28230 36168
rect 28644 36165 28672 36196
rect 30300 36196 31852 36224
rect 28537 36159 28595 36165
rect 28537 36156 28549 36159
rect 28224 36128 28549 36156
rect 28224 36116 28230 36128
rect 28537 36125 28549 36128
rect 28583 36125 28595 36159
rect 28537 36119 28595 36125
rect 28629 36159 28687 36165
rect 28629 36125 28641 36159
rect 28675 36125 28687 36159
rect 28629 36119 28687 36125
rect 25314 36088 25320 36100
rect 20027 36060 22094 36088
rect 22572 36060 25320 36088
rect 20027 36057 20039 36060
rect 19981 36051 20039 36057
rect 15013 36023 15071 36029
rect 15013 36020 15025 36023
rect 14384 35992 15025 36020
rect 15013 35989 15025 35992
rect 15059 36020 15071 36023
rect 16666 36020 16672 36032
rect 15059 35992 16672 36020
rect 15059 35989 15071 35992
rect 15013 35983 15071 35989
rect 16666 35980 16672 35992
rect 16724 35980 16730 36032
rect 17497 36023 17555 36029
rect 17497 35989 17509 36023
rect 17543 36020 17555 36023
rect 17954 36020 17960 36032
rect 17543 35992 17960 36020
rect 17543 35989 17555 35992
rect 17497 35983 17555 35989
rect 17954 35980 17960 35992
rect 18012 36020 18018 36032
rect 18506 36020 18512 36032
rect 18012 35992 18512 36020
rect 18012 35980 18018 35992
rect 18506 35980 18512 35992
rect 18564 35980 18570 36032
rect 19150 35980 19156 36032
rect 19208 36020 19214 36032
rect 21450 36020 21456 36032
rect 19208 35992 21456 36020
rect 19208 35980 19214 35992
rect 21450 35980 21456 35992
rect 21508 35980 21514 36032
rect 22066 36020 22094 36060
rect 25314 36048 25320 36060
rect 25372 36048 25378 36100
rect 26421 36091 26479 36097
rect 26421 36088 26433 36091
rect 25792 36060 26433 36088
rect 25792 36032 25820 36060
rect 26421 36057 26433 36060
rect 26467 36057 26479 36091
rect 26421 36051 26479 36057
rect 22462 36020 22468 36032
rect 22066 35992 22468 36020
rect 22462 35980 22468 35992
rect 22520 36020 22526 36032
rect 22738 36020 22744 36032
rect 22520 35992 22744 36020
rect 22520 35980 22526 35992
rect 22738 35980 22744 35992
rect 22796 35980 22802 36032
rect 23109 36023 23167 36029
rect 23109 35989 23121 36023
rect 23155 36020 23167 36023
rect 23474 36020 23480 36032
rect 23155 35992 23480 36020
rect 23155 35989 23167 35992
rect 23109 35983 23167 35989
rect 23474 35980 23480 35992
rect 23532 35980 23538 36032
rect 23658 35980 23664 36032
rect 23716 36020 23722 36032
rect 23753 36023 23811 36029
rect 23753 36020 23765 36023
rect 23716 35992 23765 36020
rect 23716 35980 23722 35992
rect 23753 35989 23765 35992
rect 23799 36020 23811 36023
rect 24302 36020 24308 36032
rect 23799 35992 24308 36020
rect 23799 35989 23811 35992
rect 23753 35983 23811 35989
rect 24302 35980 24308 35992
rect 24360 35980 24366 36032
rect 24581 36023 24639 36029
rect 24581 35989 24593 36023
rect 24627 36020 24639 36023
rect 24762 36020 24768 36032
rect 24627 35992 24768 36020
rect 24627 35989 24639 35992
rect 24581 35983 24639 35989
rect 24762 35980 24768 35992
rect 24820 35980 24826 36032
rect 25133 36023 25191 36029
rect 25133 35989 25145 36023
rect 25179 36020 25191 36023
rect 25406 36020 25412 36032
rect 25179 35992 25412 36020
rect 25179 35989 25191 35992
rect 25133 35983 25191 35989
rect 25406 35980 25412 35992
rect 25464 35980 25470 36032
rect 25774 35980 25780 36032
rect 25832 35980 25838 36032
rect 25869 36023 25927 36029
rect 25869 35989 25881 36023
rect 25915 36020 25927 36023
rect 26050 36020 26056 36032
rect 25915 35992 26056 36020
rect 25915 35989 25927 35992
rect 25869 35983 25927 35989
rect 26050 35980 26056 35992
rect 26108 35980 26114 36032
rect 28644 36020 28672 36119
rect 28718 36116 28724 36168
rect 28776 36156 28782 36168
rect 30300 36165 30328 36196
rect 31846 36184 31852 36196
rect 31904 36184 31910 36236
rect 34698 36224 34704 36236
rect 31956 36196 34704 36224
rect 31956 36168 31984 36196
rect 34698 36184 34704 36196
rect 34756 36184 34762 36236
rect 34790 36184 34796 36236
rect 34848 36224 34854 36236
rect 35544 36233 35572 36264
rect 36081 36261 36093 36295
rect 36127 36261 36139 36295
rect 36081 36255 36139 36261
rect 38473 36295 38531 36301
rect 38473 36261 38485 36295
rect 38519 36292 38531 36295
rect 38654 36292 38660 36304
rect 38519 36264 38660 36292
rect 38519 36261 38531 36264
rect 38473 36255 38531 36261
rect 35529 36227 35587 36233
rect 34848 36196 34893 36224
rect 34848 36184 34854 36196
rect 35529 36193 35541 36227
rect 35575 36193 35587 36227
rect 35529 36187 35587 36193
rect 28905 36159 28963 36165
rect 28905 36156 28917 36159
rect 28776 36128 28917 36156
rect 28776 36116 28782 36128
rect 28905 36125 28917 36128
rect 28951 36125 28963 36159
rect 28905 36119 28963 36125
rect 30285 36159 30343 36165
rect 30285 36125 30297 36159
rect 30331 36125 30343 36159
rect 30558 36156 30564 36168
rect 30519 36128 30564 36156
rect 30285 36119 30343 36125
rect 30558 36116 30564 36128
rect 30616 36116 30622 36168
rect 31389 36159 31447 36165
rect 31389 36125 31401 36159
rect 31435 36156 31447 36159
rect 31478 36156 31484 36168
rect 31435 36128 31484 36156
rect 31435 36125 31447 36128
rect 31389 36119 31447 36125
rect 31478 36116 31484 36128
rect 31536 36116 31542 36168
rect 31938 36156 31944 36168
rect 31851 36128 31944 36156
rect 31938 36116 31944 36128
rect 31996 36116 32002 36168
rect 33042 36156 33048 36168
rect 33003 36128 33048 36156
rect 33042 36116 33048 36128
rect 33100 36116 33106 36168
rect 33686 36156 33692 36168
rect 33647 36128 33692 36156
rect 33686 36116 33692 36128
rect 33744 36116 33750 36168
rect 33870 36156 33876 36168
rect 33831 36128 33876 36156
rect 33870 36116 33876 36128
rect 33928 36116 33934 36168
rect 35621 36159 35679 36165
rect 35621 36125 35633 36159
rect 35667 36156 35679 36159
rect 36096 36156 36124 36255
rect 38654 36252 38660 36264
rect 38712 36292 38718 36304
rect 38712 36264 39160 36292
rect 38712 36252 38718 36264
rect 38212 36196 38976 36224
rect 38212 36168 38240 36196
rect 36262 36156 36268 36168
rect 35667 36128 36124 36156
rect 36223 36128 36268 36156
rect 35667 36125 35679 36128
rect 35621 36119 35679 36125
rect 36262 36116 36268 36128
rect 36320 36116 36326 36168
rect 36357 36159 36415 36165
rect 36357 36125 36369 36159
rect 36403 36156 36415 36159
rect 36630 36156 36636 36168
rect 36403 36128 36636 36156
rect 36403 36125 36415 36128
rect 36357 36119 36415 36125
rect 36630 36116 36636 36128
rect 36688 36116 36694 36168
rect 36998 36156 37004 36168
rect 36959 36128 37004 36156
rect 36998 36116 37004 36128
rect 37056 36116 37062 36168
rect 37185 36159 37243 36165
rect 37185 36125 37197 36159
rect 37231 36156 37243 36159
rect 37458 36156 37464 36168
rect 37231 36128 37464 36156
rect 37231 36125 37243 36128
rect 37185 36119 37243 36125
rect 37458 36116 37464 36128
rect 37516 36156 37522 36168
rect 37734 36156 37740 36168
rect 37516 36128 37740 36156
rect 37516 36116 37522 36128
rect 37734 36116 37740 36128
rect 37792 36116 37798 36168
rect 38013 36159 38071 36165
rect 38013 36125 38025 36159
rect 38059 36125 38071 36159
rect 38194 36156 38200 36168
rect 38155 36128 38200 36156
rect 38013 36119 38071 36125
rect 30745 36091 30803 36097
rect 30745 36057 30757 36091
rect 30791 36088 30803 36091
rect 31294 36088 31300 36100
rect 30791 36060 31300 36088
rect 30791 36057 30803 36060
rect 30745 36051 30803 36057
rect 31294 36048 31300 36060
rect 31352 36048 31358 36100
rect 33229 36091 33287 36097
rect 33229 36057 33241 36091
rect 33275 36088 33287 36091
rect 33781 36091 33839 36097
rect 33781 36088 33793 36091
rect 33275 36060 33793 36088
rect 33275 36057 33287 36060
rect 33229 36051 33287 36057
rect 33781 36057 33793 36060
rect 33827 36057 33839 36091
rect 33781 36051 33839 36057
rect 35802 36048 35808 36100
rect 35860 36088 35866 36100
rect 36081 36091 36139 36097
rect 36081 36088 36093 36091
rect 35860 36060 36093 36088
rect 35860 36048 35866 36060
rect 36081 36057 36093 36060
rect 36127 36057 36139 36091
rect 36081 36051 36139 36057
rect 31754 36020 31760 36032
rect 28644 35992 31760 36020
rect 31754 35980 31760 35992
rect 31812 36020 31818 36032
rect 32214 36020 32220 36032
rect 31812 35992 32220 36020
rect 31812 35980 31818 35992
rect 32214 35980 32220 35992
rect 32272 35980 32278 36032
rect 36096 36020 36124 36051
rect 36446 36048 36452 36100
rect 36504 36088 36510 36100
rect 36817 36091 36875 36097
rect 36817 36088 36829 36091
rect 36504 36060 36829 36088
rect 36504 36048 36510 36060
rect 36817 36057 36829 36060
rect 36863 36088 36875 36091
rect 38028 36088 38056 36119
rect 38194 36116 38200 36128
rect 38252 36116 38258 36168
rect 38948 36165 38976 36196
rect 39132 36165 39160 36264
rect 40034 36252 40040 36304
rect 40092 36252 40098 36304
rect 40144 36301 40172 36332
rect 40402 36320 40408 36372
rect 40460 36360 40466 36372
rect 40460 36332 41460 36360
rect 40460 36320 40466 36332
rect 40129 36295 40187 36301
rect 40129 36261 40141 36295
rect 40175 36261 40187 36295
rect 41432 36292 41460 36332
rect 41874 36320 41880 36372
rect 41932 36360 41938 36372
rect 41969 36363 42027 36369
rect 41969 36360 41981 36363
rect 41932 36332 41981 36360
rect 41932 36320 41938 36332
rect 41969 36329 41981 36332
rect 42015 36360 42027 36363
rect 42610 36360 42616 36372
rect 42015 36332 42616 36360
rect 42015 36329 42027 36332
rect 41969 36323 42027 36329
rect 42610 36320 42616 36332
rect 42668 36320 42674 36372
rect 47210 36360 47216 36372
rect 47171 36332 47216 36360
rect 47210 36320 47216 36332
rect 47268 36320 47274 36372
rect 42429 36295 42487 36301
rect 42429 36292 42441 36295
rect 41432 36264 42441 36292
rect 40129 36255 40187 36261
rect 42429 36261 42441 36264
rect 42475 36261 42487 36295
rect 42429 36255 42487 36261
rect 40052 36224 40080 36252
rect 40052 36196 40540 36224
rect 38933 36159 38991 36165
rect 38933 36125 38945 36159
rect 38979 36125 38991 36159
rect 38933 36119 38991 36125
rect 39117 36159 39175 36165
rect 39117 36125 39129 36159
rect 39163 36156 39175 36159
rect 39206 36156 39212 36168
rect 39163 36128 39212 36156
rect 39163 36125 39175 36128
rect 39117 36119 39175 36125
rect 39206 36116 39212 36128
rect 39264 36116 39270 36168
rect 39850 36116 39856 36168
rect 39908 36156 39914 36168
rect 40037 36159 40095 36165
rect 40037 36156 40049 36159
rect 39908 36128 40049 36156
rect 39908 36116 39914 36128
rect 40037 36125 40049 36128
rect 40083 36125 40095 36159
rect 40037 36119 40095 36125
rect 40126 36116 40132 36168
rect 40184 36156 40190 36168
rect 40512 36165 40540 36196
rect 40221 36159 40279 36165
rect 40221 36156 40233 36159
rect 40184 36128 40233 36156
rect 40184 36116 40190 36128
rect 40221 36125 40233 36128
rect 40267 36125 40279 36159
rect 40221 36119 40279 36125
rect 40313 36159 40371 36165
rect 40313 36125 40325 36159
rect 40359 36125 40371 36159
rect 40313 36119 40371 36125
rect 40497 36159 40555 36165
rect 40497 36125 40509 36159
rect 40543 36125 40555 36159
rect 40497 36119 40555 36125
rect 36863 36060 38056 36088
rect 40328 36088 40356 36119
rect 40862 36116 40868 36168
rect 40920 36156 40926 36168
rect 41141 36159 41199 36165
rect 41141 36156 41153 36159
rect 40920 36128 41153 36156
rect 40920 36116 40926 36128
rect 41141 36125 41153 36128
rect 41187 36125 41199 36159
rect 41361 36159 41419 36165
rect 41141 36119 41199 36125
rect 40957 36091 41015 36097
rect 41230 36094 41236 36146
rect 41288 36134 41294 36146
rect 41288 36106 41333 36134
rect 41361 36125 41373 36159
rect 41407 36125 41419 36159
rect 41361 36119 41419 36125
rect 41288 36094 41294 36106
rect 40957 36088 40969 36091
rect 40328 36060 40969 36088
rect 36863 36057 36875 36060
rect 36817 36051 36875 36057
rect 40957 36057 40969 36060
rect 41003 36057 41015 36091
rect 40957 36051 41015 36057
rect 39025 36023 39083 36029
rect 39025 36020 39037 36023
rect 36096 35992 39037 36020
rect 39025 35989 39037 35992
rect 39071 35989 39083 36023
rect 39850 36020 39856 36032
rect 39811 35992 39856 36020
rect 39025 35983 39083 35989
rect 39850 35980 39856 35992
rect 39908 35980 39914 36032
rect 40310 35980 40316 36032
rect 40368 36020 40374 36032
rect 41386 36020 41414 36119
rect 47854 36088 47860 36100
rect 47815 36060 47860 36088
rect 47854 36048 47860 36060
rect 47912 36048 47918 36100
rect 48038 36088 48044 36100
rect 47999 36060 48044 36088
rect 48038 36048 48044 36060
rect 48096 36048 48102 36100
rect 42978 36020 42984 36032
rect 40368 35992 41414 36020
rect 42939 35992 42984 36020
rect 40368 35980 40374 35992
rect 42978 35980 42984 35992
rect 43036 35980 43042 36032
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 10226 35776 10232 35828
rect 10284 35816 10290 35828
rect 10873 35819 10931 35825
rect 10873 35816 10885 35819
rect 10284 35788 10885 35816
rect 10284 35776 10290 35788
rect 10873 35785 10885 35788
rect 10919 35785 10931 35819
rect 10873 35779 10931 35785
rect 12161 35819 12219 35825
rect 12161 35785 12173 35819
rect 12207 35816 12219 35819
rect 12710 35816 12716 35828
rect 12207 35788 12434 35816
rect 12671 35788 12716 35816
rect 12207 35785 12219 35788
rect 12161 35779 12219 35785
rect 12406 35748 12434 35788
rect 12710 35776 12716 35788
rect 12768 35776 12774 35828
rect 13262 35816 13268 35828
rect 13223 35788 13268 35816
rect 13262 35776 13268 35788
rect 13320 35776 13326 35828
rect 15749 35819 15807 35825
rect 15749 35785 15761 35819
rect 15795 35785 15807 35819
rect 15749 35779 15807 35785
rect 17037 35819 17095 35825
rect 17037 35785 17049 35819
rect 17083 35816 17095 35819
rect 17494 35816 17500 35828
rect 17083 35788 17500 35816
rect 17083 35785 17095 35788
rect 17037 35779 17095 35785
rect 12986 35748 12992 35760
rect 12406 35720 12992 35748
rect 12986 35708 12992 35720
rect 13044 35708 13050 35760
rect 15764 35748 15792 35779
rect 17494 35776 17500 35788
rect 17552 35776 17558 35828
rect 17788 35788 18552 35816
rect 17788 35748 17816 35788
rect 15764 35720 17816 35748
rect 17865 35751 17923 35757
rect 17865 35717 17877 35751
rect 17911 35748 17923 35751
rect 18230 35748 18236 35760
rect 17911 35720 18236 35748
rect 17911 35717 17923 35720
rect 17865 35711 17923 35717
rect 18230 35708 18236 35720
rect 18288 35708 18294 35760
rect 18524 35748 18552 35788
rect 19794 35776 19800 35828
rect 19852 35816 19858 35828
rect 20625 35819 20683 35825
rect 20625 35816 20637 35819
rect 19852 35788 20637 35816
rect 19852 35776 19858 35788
rect 20625 35785 20637 35788
rect 20671 35785 20683 35819
rect 20625 35779 20683 35785
rect 20993 35819 21051 35825
rect 20993 35785 21005 35819
rect 21039 35816 21051 35819
rect 21910 35816 21916 35828
rect 21039 35788 21916 35816
rect 21039 35785 21051 35788
rect 20993 35779 21051 35785
rect 21910 35776 21916 35788
rect 21968 35776 21974 35828
rect 24026 35816 24032 35828
rect 23987 35788 24032 35816
rect 24026 35776 24032 35788
rect 24084 35776 24090 35828
rect 24670 35776 24676 35828
rect 24728 35776 24734 35828
rect 25133 35819 25191 35825
rect 25133 35785 25145 35819
rect 25179 35816 25191 35819
rect 25406 35816 25412 35828
rect 25179 35788 25412 35816
rect 25179 35785 25191 35788
rect 25133 35779 25191 35785
rect 25406 35776 25412 35788
rect 25464 35776 25470 35828
rect 25498 35776 25504 35828
rect 25556 35816 25562 35828
rect 30006 35816 30012 35828
rect 25556 35788 30012 35816
rect 25556 35776 25562 35788
rect 30006 35776 30012 35788
rect 30064 35776 30070 35828
rect 30650 35776 30656 35828
rect 30708 35816 30714 35828
rect 31113 35819 31171 35825
rect 31113 35816 31125 35819
rect 30708 35788 31125 35816
rect 30708 35776 30714 35788
rect 31113 35785 31125 35788
rect 31159 35785 31171 35819
rect 31113 35779 31171 35785
rect 31294 35776 31300 35828
rect 31352 35816 31358 35828
rect 32401 35819 32459 35825
rect 32401 35816 32413 35819
rect 31352 35788 32413 35816
rect 31352 35776 31358 35788
rect 32401 35785 32413 35788
rect 32447 35816 32459 35819
rect 33134 35816 33140 35828
rect 32447 35788 33140 35816
rect 32447 35785 32459 35788
rect 32401 35779 32459 35785
rect 33134 35776 33140 35788
rect 33192 35776 33198 35828
rect 33410 35776 33416 35828
rect 33468 35816 33474 35828
rect 33597 35819 33655 35825
rect 33597 35816 33609 35819
rect 33468 35788 33609 35816
rect 33468 35776 33474 35788
rect 33597 35785 33609 35788
rect 33643 35816 33655 35819
rect 33686 35816 33692 35828
rect 33643 35788 33692 35816
rect 33643 35785 33655 35788
rect 33597 35779 33655 35785
rect 33686 35776 33692 35788
rect 33744 35776 33750 35828
rect 35526 35816 35532 35828
rect 35487 35788 35532 35816
rect 35526 35776 35532 35788
rect 35584 35776 35590 35828
rect 36173 35819 36231 35825
rect 36173 35785 36185 35819
rect 36219 35816 36231 35819
rect 36262 35816 36268 35828
rect 36219 35788 36268 35816
rect 36219 35785 36231 35788
rect 36173 35779 36231 35785
rect 36262 35776 36268 35788
rect 36320 35776 36326 35828
rect 38194 35776 38200 35828
rect 38252 35816 38258 35828
rect 38473 35819 38531 35825
rect 38473 35816 38485 35819
rect 38252 35788 38485 35816
rect 38252 35776 38258 35788
rect 38473 35785 38485 35788
rect 38519 35785 38531 35819
rect 38473 35779 38531 35785
rect 38838 35776 38844 35828
rect 38896 35816 38902 35828
rect 48038 35816 48044 35828
rect 38896 35788 39252 35816
rect 47999 35788 48044 35816
rect 38896 35776 38902 35788
rect 24210 35748 24216 35760
rect 18524 35720 24216 35748
rect 24210 35708 24216 35720
rect 24268 35708 24274 35760
rect 24688 35748 24716 35776
rect 24504 35720 24716 35748
rect 14274 35680 14280 35692
rect 14235 35652 14280 35680
rect 14274 35640 14280 35652
rect 14332 35640 14338 35692
rect 14461 35683 14519 35689
rect 14461 35649 14473 35683
rect 14507 35649 14519 35683
rect 15378 35680 15384 35692
rect 15339 35652 15384 35680
rect 14461 35643 14519 35649
rect 13814 35572 13820 35624
rect 13872 35612 13878 35624
rect 14476 35612 14504 35643
rect 15378 35640 15384 35652
rect 15436 35640 15442 35692
rect 16574 35640 16580 35692
rect 16632 35680 16638 35692
rect 16669 35683 16727 35689
rect 16669 35680 16681 35683
rect 16632 35652 16681 35680
rect 16632 35640 16638 35652
rect 16669 35649 16681 35652
rect 16715 35649 16727 35683
rect 16669 35643 16727 35649
rect 15470 35612 15476 35624
rect 13872 35584 14504 35612
rect 15431 35584 15476 35612
rect 13872 35572 13878 35584
rect 15470 35572 15476 35584
rect 15528 35572 15534 35624
rect 16684 35612 16712 35643
rect 16850 35640 16856 35692
rect 16908 35680 16914 35692
rect 17218 35680 17224 35692
rect 16908 35652 17224 35680
rect 16908 35640 16914 35652
rect 17218 35640 17224 35652
rect 17276 35640 17282 35692
rect 18141 35683 18199 35689
rect 18141 35649 18153 35683
rect 18187 35680 18199 35683
rect 18506 35680 18512 35692
rect 18187 35652 18512 35680
rect 18187 35649 18199 35652
rect 18141 35643 18199 35649
rect 18506 35640 18512 35652
rect 18564 35640 18570 35692
rect 18601 35683 18659 35689
rect 18601 35649 18613 35683
rect 18647 35680 18659 35683
rect 18966 35680 18972 35692
rect 18647 35652 18972 35680
rect 18647 35649 18659 35652
rect 18601 35643 18659 35649
rect 18966 35640 18972 35652
rect 19024 35640 19030 35692
rect 19058 35640 19064 35692
rect 19116 35680 19122 35692
rect 19116 35652 19161 35680
rect 19116 35640 19122 35652
rect 19426 35640 19432 35692
rect 19484 35680 19490 35692
rect 19705 35683 19763 35689
rect 19705 35680 19717 35683
rect 19484 35652 19717 35680
rect 19484 35640 19490 35652
rect 19705 35649 19717 35652
rect 19751 35649 19763 35683
rect 19886 35680 19892 35692
rect 19847 35652 19892 35680
rect 19705 35643 19763 35649
rect 19886 35640 19892 35652
rect 19944 35640 19950 35692
rect 19978 35640 19984 35692
rect 20036 35680 20042 35692
rect 20533 35683 20591 35689
rect 20533 35680 20545 35683
rect 20036 35652 20545 35680
rect 20036 35640 20042 35652
rect 20533 35649 20545 35652
rect 20579 35649 20591 35683
rect 20806 35680 20812 35692
rect 20767 35652 20812 35680
rect 20533 35643 20591 35649
rect 20806 35640 20812 35652
rect 20864 35640 20870 35692
rect 21450 35640 21456 35692
rect 21508 35680 21514 35692
rect 22370 35680 22376 35692
rect 21508 35652 22376 35680
rect 21508 35640 21514 35652
rect 22370 35640 22376 35652
rect 22428 35640 22434 35692
rect 22554 35680 22560 35692
rect 22515 35652 22560 35680
rect 22554 35640 22560 35652
rect 22612 35640 22618 35692
rect 24504 35689 24532 35720
rect 25958 35708 25964 35760
rect 26016 35748 26022 35760
rect 26016 35720 26188 35748
rect 26016 35708 26022 35720
rect 24489 35683 24547 35689
rect 24489 35649 24501 35683
rect 24535 35649 24547 35683
rect 24670 35680 24676 35692
rect 24631 35652 24676 35680
rect 24489 35643 24547 35649
rect 24670 35640 24676 35652
rect 24728 35640 24734 35692
rect 24765 35683 24823 35689
rect 24765 35649 24777 35683
rect 24811 35649 24823 35683
rect 24765 35643 24823 35649
rect 24857 35683 24915 35689
rect 24857 35649 24869 35683
rect 24903 35680 24915 35683
rect 24946 35680 24952 35692
rect 24903 35652 24952 35680
rect 24903 35649 24915 35652
rect 24857 35643 24915 35649
rect 17494 35612 17500 35624
rect 16684 35584 17500 35612
rect 17494 35572 17500 35584
rect 17552 35572 17558 35624
rect 18414 35572 18420 35624
rect 18472 35612 18478 35624
rect 18785 35615 18843 35621
rect 18785 35612 18797 35615
rect 18472 35584 18797 35612
rect 18472 35572 18478 35584
rect 18785 35581 18797 35584
rect 18831 35581 18843 35615
rect 18785 35575 18843 35581
rect 18874 35572 18880 35624
rect 18932 35612 18938 35624
rect 19245 35615 19303 35621
rect 18932 35584 18977 35612
rect 18932 35572 18938 35584
rect 19245 35581 19257 35615
rect 19291 35612 19303 35615
rect 24780 35612 24808 35643
rect 24946 35640 24952 35652
rect 25004 35640 25010 35692
rect 25777 35683 25835 35689
rect 25777 35649 25789 35683
rect 25823 35649 25835 35683
rect 25777 35643 25835 35649
rect 25593 35615 25651 35621
rect 25593 35612 25605 35615
rect 19291 35584 22094 35612
rect 24780 35584 25605 35612
rect 19291 35581 19303 35584
rect 19245 35575 19303 35581
rect 13722 35504 13728 35556
rect 13780 35544 13786 35556
rect 17954 35544 17960 35556
rect 13780 35516 17960 35544
rect 13780 35504 13786 35516
rect 17954 35504 17960 35516
rect 18012 35504 18018 35556
rect 18049 35547 18107 35553
rect 18049 35513 18061 35547
rect 18095 35513 18107 35547
rect 18049 35507 18107 35513
rect 18141 35547 18199 35553
rect 18141 35513 18153 35547
rect 18187 35544 18199 35547
rect 18969 35547 19027 35553
rect 18969 35544 18981 35547
rect 18187 35516 18981 35544
rect 18187 35513 18199 35516
rect 18141 35507 18199 35513
rect 18969 35513 18981 35516
rect 19015 35513 19027 35547
rect 22066 35544 22094 35584
rect 25593 35581 25605 35584
rect 25639 35581 25651 35615
rect 25593 35575 25651 35581
rect 23750 35544 23756 35556
rect 22066 35516 23756 35544
rect 18969 35507 19027 35513
rect 9122 35436 9128 35488
rect 9180 35476 9186 35488
rect 10321 35479 10379 35485
rect 10321 35476 10333 35479
rect 9180 35448 10333 35476
rect 9180 35436 9186 35448
rect 10321 35445 10333 35448
rect 10367 35445 10379 35479
rect 10321 35439 10379 35445
rect 11609 35479 11667 35485
rect 11609 35445 11621 35479
rect 11655 35476 11667 35479
rect 11882 35476 11888 35488
rect 11655 35448 11888 35476
rect 11655 35445 11667 35448
rect 11609 35439 11667 35445
rect 11882 35436 11888 35448
rect 11940 35436 11946 35488
rect 13817 35479 13875 35485
rect 13817 35445 13829 35479
rect 13863 35476 13875 35479
rect 14090 35476 14096 35488
rect 13863 35448 14096 35476
rect 13863 35445 13875 35448
rect 13817 35439 13875 35445
rect 14090 35436 14096 35448
rect 14148 35436 14154 35488
rect 14458 35476 14464 35488
rect 14419 35448 14464 35476
rect 14458 35436 14464 35448
rect 14516 35436 14522 35488
rect 18064 35476 18092 35507
rect 23750 35504 23756 35516
rect 23808 35504 23814 35556
rect 24394 35504 24400 35556
rect 24452 35544 24458 35556
rect 25792 35544 25820 35643
rect 25866 35640 25872 35692
rect 25924 35680 25930 35692
rect 26160 35689 26188 35720
rect 26786 35708 26792 35760
rect 26844 35748 26850 35760
rect 27154 35748 27160 35760
rect 26844 35720 27160 35748
rect 26844 35708 26850 35720
rect 27154 35708 27160 35720
rect 27212 35748 27218 35760
rect 28261 35751 28319 35757
rect 28261 35748 28273 35751
rect 27212 35720 28273 35748
rect 27212 35708 27218 35720
rect 28261 35717 28273 35720
rect 28307 35717 28319 35751
rect 28261 35711 28319 35717
rect 29181 35751 29239 35757
rect 29181 35717 29193 35751
rect 29227 35748 29239 35751
rect 30282 35748 30288 35760
rect 29227 35720 30288 35748
rect 29227 35717 29239 35720
rect 29181 35711 29239 35717
rect 30282 35708 30288 35720
rect 30340 35708 30346 35760
rect 34054 35748 34060 35760
rect 34015 35720 34060 35748
rect 30668 35692 30880 35714
rect 34054 35708 34060 35720
rect 34112 35708 34118 35760
rect 38105 35751 38163 35757
rect 35452 35720 36308 35748
rect 26145 35683 26203 35689
rect 25924 35652 25969 35680
rect 25924 35640 25930 35652
rect 26145 35649 26157 35683
rect 26191 35649 26203 35683
rect 26145 35643 26203 35649
rect 26973 35683 27031 35689
rect 26973 35649 26985 35683
rect 27019 35680 27031 35683
rect 27614 35680 27620 35692
rect 27019 35652 27620 35680
rect 27019 35649 27031 35652
rect 26973 35643 27031 35649
rect 27614 35640 27620 35652
rect 27672 35640 27678 35692
rect 29086 35640 29092 35692
rect 29144 35680 29150 35692
rect 29365 35683 29423 35689
rect 29365 35680 29377 35683
rect 29144 35652 29377 35680
rect 29144 35640 29150 35652
rect 29365 35649 29377 35652
rect 29411 35649 29423 35683
rect 29365 35643 29423 35649
rect 30098 35640 30104 35692
rect 30156 35680 30162 35692
rect 30668 35689 30840 35692
rect 30377 35683 30435 35689
rect 30377 35680 30389 35683
rect 30156 35652 30389 35680
rect 30156 35640 30162 35652
rect 30377 35649 30389 35652
rect 30423 35649 30435 35683
rect 30561 35683 30619 35689
rect 30561 35680 30573 35683
rect 30377 35643 30435 35649
rect 30484 35652 30573 35680
rect 26050 35612 26056 35624
rect 26011 35584 26056 35612
rect 26050 35572 26056 35584
rect 26108 35572 26114 35624
rect 27249 35615 27307 35621
rect 27249 35612 27261 35615
rect 26896 35584 27261 35612
rect 24452 35516 25820 35544
rect 24452 35504 24458 35516
rect 18322 35476 18328 35488
rect 18064 35448 18328 35476
rect 18322 35436 18328 35448
rect 18380 35476 18386 35488
rect 19705 35479 19763 35485
rect 19705 35476 19717 35479
rect 18380 35448 19717 35476
rect 18380 35436 18386 35448
rect 19705 35445 19717 35448
rect 19751 35445 19763 35479
rect 19705 35439 19763 35445
rect 22370 35436 22376 35488
rect 22428 35476 22434 35488
rect 22465 35479 22523 35485
rect 22465 35476 22477 35479
rect 22428 35448 22477 35476
rect 22428 35436 22434 35448
rect 22465 35445 22477 35448
rect 22511 35476 22523 35479
rect 22738 35476 22744 35488
rect 22511 35448 22744 35476
rect 22511 35445 22523 35448
rect 22465 35439 22523 35445
rect 22738 35436 22744 35448
rect 22796 35436 22802 35488
rect 23477 35479 23535 35485
rect 23477 35445 23489 35479
rect 23523 35476 23535 35479
rect 23566 35476 23572 35488
rect 23523 35448 23572 35476
rect 23523 35445 23535 35448
rect 23477 35439 23535 35445
rect 23566 35436 23572 35448
rect 23624 35436 23630 35488
rect 25130 35436 25136 35488
rect 25188 35476 25194 35488
rect 26896 35476 26924 35584
rect 27249 35581 27261 35584
rect 27295 35612 27307 35615
rect 27706 35612 27712 35624
rect 27295 35584 27712 35612
rect 27295 35581 27307 35584
rect 27249 35575 27307 35581
rect 27706 35572 27712 35584
rect 27764 35572 27770 35624
rect 27801 35615 27859 35621
rect 27801 35581 27813 35615
rect 27847 35612 27859 35615
rect 29454 35612 29460 35624
rect 27847 35584 29460 35612
rect 27847 35581 27859 35584
rect 27801 35575 27859 35581
rect 26970 35504 26976 35556
rect 27028 35544 27034 35556
rect 27816 35544 27844 35575
rect 29454 35572 29460 35584
rect 29512 35572 29518 35624
rect 29641 35615 29699 35621
rect 29641 35581 29653 35615
rect 29687 35612 29699 35615
rect 29822 35612 29828 35624
rect 29687 35584 29828 35612
rect 29687 35581 29699 35584
rect 29641 35575 29699 35581
rect 29822 35572 29828 35584
rect 29880 35572 29886 35624
rect 30282 35572 30288 35624
rect 30340 35612 30346 35624
rect 30484 35612 30512 35652
rect 30561 35649 30573 35652
rect 30607 35649 30619 35683
rect 30561 35643 30619 35649
rect 30653 35686 30840 35689
rect 30653 35683 30711 35686
rect 30653 35649 30665 35683
rect 30699 35649 30711 35683
rect 30653 35643 30711 35649
rect 30834 35640 30840 35686
rect 30892 35640 30898 35692
rect 30929 35683 30987 35689
rect 30929 35649 30941 35683
rect 30975 35680 30987 35683
rect 31478 35680 31484 35692
rect 30975 35652 31484 35680
rect 30975 35649 30987 35652
rect 30929 35643 30987 35649
rect 31478 35640 31484 35652
rect 31536 35640 31542 35692
rect 32214 35680 32220 35692
rect 32175 35652 32220 35680
rect 32214 35640 32220 35652
rect 32272 35640 32278 35692
rect 32398 35680 32404 35692
rect 32359 35652 32404 35680
rect 32398 35640 32404 35652
rect 32456 35640 32462 35692
rect 33413 35683 33471 35689
rect 33413 35649 33425 35683
rect 33459 35680 33471 35683
rect 33502 35680 33508 35692
rect 33459 35652 33508 35680
rect 33459 35649 33471 35652
rect 33413 35643 33471 35649
rect 33502 35640 33508 35652
rect 33560 35640 33566 35692
rect 34238 35640 34244 35692
rect 34296 35680 34302 35692
rect 34333 35683 34391 35689
rect 34333 35680 34345 35683
rect 34296 35652 34345 35680
rect 34296 35640 34302 35652
rect 34333 35649 34345 35652
rect 34379 35680 34391 35683
rect 34422 35680 34428 35692
rect 34379 35652 34428 35680
rect 34379 35649 34391 35652
rect 34333 35643 34391 35649
rect 34422 35640 34428 35652
rect 34480 35640 34486 35692
rect 35452 35689 35480 35720
rect 36280 35689 36308 35720
rect 38105 35717 38117 35751
rect 38151 35717 38163 35751
rect 38105 35711 38163 35717
rect 35437 35683 35495 35689
rect 35437 35649 35449 35683
rect 35483 35649 35495 35683
rect 35437 35643 35495 35649
rect 35621 35683 35679 35689
rect 35621 35649 35633 35683
rect 35667 35649 35679 35683
rect 35621 35643 35679 35649
rect 36265 35683 36323 35689
rect 36265 35649 36277 35683
rect 36311 35680 36323 35683
rect 36446 35680 36452 35692
rect 36311 35652 36452 35680
rect 36311 35649 36323 35652
rect 36265 35643 36323 35649
rect 30340 35584 30512 35612
rect 30340 35572 30346 35584
rect 30742 35572 30748 35624
rect 30800 35612 30806 35624
rect 33229 35615 33287 35621
rect 30800 35584 30845 35612
rect 30800 35572 30806 35584
rect 33229 35581 33241 35615
rect 33275 35612 33287 35615
rect 33594 35612 33600 35624
rect 33275 35584 33600 35612
rect 33275 35581 33287 35584
rect 33229 35575 33287 35581
rect 27028 35516 27844 35544
rect 27028 35504 27034 35516
rect 28810 35504 28816 35556
rect 28868 35544 28874 35556
rect 28868 35516 30696 35544
rect 28868 35504 28874 35516
rect 27062 35476 27068 35488
rect 25188 35448 26924 35476
rect 27023 35448 27068 35476
rect 25188 35436 25194 35448
rect 27062 35436 27068 35448
rect 27120 35436 27126 35488
rect 27157 35479 27215 35485
rect 27157 35445 27169 35479
rect 27203 35476 27215 35479
rect 27246 35476 27252 35488
rect 27203 35448 27252 35476
rect 27203 35445 27215 35448
rect 27157 35439 27215 35445
rect 27246 35436 27252 35448
rect 27304 35436 27310 35488
rect 29546 35476 29552 35488
rect 29507 35448 29552 35476
rect 29546 35436 29552 35448
rect 29604 35436 29610 35488
rect 30668 35476 30696 35516
rect 33244 35476 33272 35575
rect 33594 35572 33600 35584
rect 33652 35572 33658 35624
rect 35636 35612 35664 35643
rect 36446 35640 36452 35652
rect 36504 35640 36510 35692
rect 36538 35640 36544 35692
rect 36596 35680 36602 35692
rect 36998 35680 37004 35692
rect 36596 35652 37004 35680
rect 36596 35640 36602 35652
rect 36998 35640 37004 35652
rect 37056 35680 37062 35692
rect 37277 35683 37335 35689
rect 37277 35680 37289 35683
rect 37056 35652 37289 35680
rect 37056 35640 37062 35652
rect 37277 35649 37289 35652
rect 37323 35649 37335 35683
rect 37277 35643 37335 35649
rect 37458 35640 37464 35692
rect 37516 35680 37522 35692
rect 38120 35680 38148 35711
rect 38286 35708 38292 35760
rect 38344 35757 38350 35760
rect 39224 35757 39252 35788
rect 48038 35776 48044 35788
rect 48096 35776 48102 35828
rect 38344 35751 38363 35757
rect 38351 35748 38363 35751
rect 39209 35751 39267 35757
rect 38351 35720 38976 35748
rect 38351 35717 38363 35720
rect 38344 35711 38363 35717
rect 38344 35708 38350 35711
rect 38838 35680 38844 35692
rect 37516 35652 37609 35680
rect 38120 35652 38844 35680
rect 37516 35640 37522 35652
rect 38838 35640 38844 35652
rect 38896 35640 38902 35692
rect 38948 35689 38976 35720
rect 39209 35717 39221 35751
rect 39255 35717 39267 35751
rect 39209 35711 39267 35717
rect 38933 35683 38991 35689
rect 38933 35649 38945 35683
rect 38979 35649 38991 35683
rect 38933 35643 38991 35649
rect 39022 35640 39028 35692
rect 39080 35680 39086 35692
rect 39080 35652 39125 35680
rect 39080 35640 39086 35652
rect 40034 35640 40040 35692
rect 40092 35680 40098 35692
rect 40159 35683 40217 35689
rect 40159 35680 40171 35683
rect 40092 35652 40171 35680
rect 40092 35640 40098 35652
rect 40159 35649 40171 35652
rect 40205 35649 40217 35683
rect 40159 35643 40217 35649
rect 40310 35640 40316 35692
rect 40368 35680 40374 35692
rect 40368 35652 40413 35680
rect 40368 35640 40374 35652
rect 37369 35615 37427 35621
rect 37369 35612 37381 35615
rect 35636 35584 37381 35612
rect 37369 35581 37381 35584
rect 37415 35581 37427 35615
rect 37476 35612 37504 35640
rect 37476 35584 41414 35612
rect 37369 35575 37427 35581
rect 39206 35544 39212 35556
rect 39167 35516 39212 35544
rect 39206 35504 39212 35516
rect 39264 35504 39270 35556
rect 41386 35544 41414 35584
rect 41386 35516 43024 35544
rect 42996 35488 43024 35516
rect 34790 35476 34796 35488
rect 30668 35448 33272 35476
rect 34751 35448 34796 35476
rect 34790 35436 34796 35448
rect 34848 35436 34854 35488
rect 38289 35479 38347 35485
rect 38289 35445 38301 35479
rect 38335 35476 38347 35479
rect 39022 35476 39028 35488
rect 38335 35448 39028 35476
rect 38335 35445 38347 35448
rect 38289 35439 38347 35445
rect 39022 35436 39028 35448
rect 39080 35436 39086 35488
rect 40126 35476 40132 35488
rect 40087 35448 40132 35476
rect 40126 35436 40132 35448
rect 40184 35436 40190 35488
rect 40865 35479 40923 35485
rect 40865 35445 40877 35479
rect 40911 35476 40923 35479
rect 41414 35476 41420 35488
rect 40911 35448 41420 35476
rect 40911 35445 40923 35448
rect 40865 35439 40923 35445
rect 41414 35436 41420 35448
rect 41472 35436 41478 35488
rect 41506 35436 41512 35488
rect 41564 35476 41570 35488
rect 42150 35476 42156 35488
rect 41564 35448 42156 35476
rect 41564 35436 41570 35448
rect 42150 35436 42156 35448
rect 42208 35476 42214 35488
rect 42429 35479 42487 35485
rect 42429 35476 42441 35479
rect 42208 35448 42441 35476
rect 42208 35436 42214 35448
rect 42429 35445 42441 35448
rect 42475 35445 42487 35479
rect 42429 35439 42487 35445
rect 42978 35436 42984 35488
rect 43036 35476 43042 35488
rect 43073 35479 43131 35485
rect 43073 35476 43085 35479
rect 43036 35448 43085 35476
rect 43036 35436 43042 35448
rect 43073 35445 43085 35448
rect 43119 35476 43131 35479
rect 43254 35476 43260 35488
rect 43119 35448 43260 35476
rect 43119 35445 43131 35448
rect 43073 35439 43131 35445
rect 43254 35436 43260 35448
rect 43312 35436 43318 35488
rect 43530 35476 43536 35488
rect 43491 35448 43536 35476
rect 43530 35436 43536 35448
rect 43588 35436 43594 35488
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 10229 35275 10287 35281
rect 10229 35241 10241 35275
rect 10275 35272 10287 35275
rect 10781 35275 10839 35281
rect 10781 35272 10793 35275
rect 10275 35244 10793 35272
rect 10275 35241 10287 35244
rect 10229 35235 10287 35241
rect 10781 35241 10793 35244
rect 10827 35272 10839 35275
rect 10870 35272 10876 35284
rect 10827 35244 10876 35272
rect 10827 35241 10839 35244
rect 10781 35235 10839 35241
rect 10870 35232 10876 35244
rect 10928 35232 10934 35284
rect 11333 35275 11391 35281
rect 11333 35241 11345 35275
rect 11379 35272 11391 35275
rect 13541 35275 13599 35281
rect 11379 35244 13492 35272
rect 11379 35241 11391 35244
rect 11333 35235 11391 35241
rect 12805 35207 12863 35213
rect 12805 35173 12817 35207
rect 12851 35173 12863 35207
rect 13464 35204 13492 35244
rect 13541 35241 13553 35275
rect 13587 35272 13599 35275
rect 15289 35275 15347 35281
rect 13587 35244 15148 35272
rect 13587 35241 13599 35244
rect 13541 35235 13599 35241
rect 14090 35204 14096 35216
rect 13464 35176 14096 35204
rect 12805 35167 12863 35173
rect 12618 35136 12624 35148
rect 6886 35108 12624 35136
rect 1946 34960 1952 35012
rect 2004 35000 2010 35012
rect 6886 35000 6914 35108
rect 12618 35096 12624 35108
rect 12676 35096 12682 35148
rect 12820 35136 12848 35167
rect 14090 35164 14096 35176
rect 14148 35164 14154 35216
rect 15120 35145 15148 35244
rect 15289 35241 15301 35275
rect 15335 35272 15347 35275
rect 15562 35272 15568 35284
rect 15335 35244 15568 35272
rect 15335 35241 15347 35244
rect 15289 35235 15347 35241
rect 15562 35232 15568 35244
rect 15620 35232 15626 35284
rect 17773 35275 17831 35281
rect 17773 35241 17785 35275
rect 17819 35272 17831 35275
rect 18230 35272 18236 35284
rect 17819 35244 18236 35272
rect 17819 35241 17831 35244
rect 17773 35235 17831 35241
rect 18230 35232 18236 35244
rect 18288 35232 18294 35284
rect 18322 35232 18328 35284
rect 18380 35272 18386 35284
rect 18693 35275 18751 35281
rect 18380 35244 18425 35272
rect 18380 35232 18386 35244
rect 18693 35241 18705 35275
rect 18739 35272 18751 35275
rect 18874 35272 18880 35284
rect 18739 35244 18880 35272
rect 18739 35241 18751 35244
rect 18693 35235 18751 35241
rect 18874 35232 18880 35244
rect 18932 35232 18938 35284
rect 19337 35275 19395 35281
rect 19337 35241 19349 35275
rect 19383 35272 19395 35275
rect 19426 35272 19432 35284
rect 19383 35244 19432 35272
rect 19383 35241 19395 35244
rect 19337 35235 19395 35241
rect 19426 35232 19432 35244
rect 19484 35232 19490 35284
rect 19886 35232 19892 35284
rect 19944 35232 19950 35284
rect 19981 35275 20039 35281
rect 19981 35241 19993 35275
rect 20027 35272 20039 35275
rect 20806 35272 20812 35284
rect 20027 35244 20812 35272
rect 20027 35241 20039 35244
rect 19981 35235 20039 35241
rect 20806 35232 20812 35244
rect 20864 35232 20870 35284
rect 21085 35275 21143 35281
rect 21085 35241 21097 35275
rect 21131 35272 21143 35275
rect 22278 35272 22284 35284
rect 21131 35244 22284 35272
rect 21131 35241 21143 35244
rect 21085 35235 21143 35241
rect 22278 35232 22284 35244
rect 22336 35232 22342 35284
rect 24762 35232 24768 35284
rect 24820 35272 24826 35284
rect 26970 35272 26976 35284
rect 24820 35244 26976 35272
rect 24820 35232 24826 35244
rect 26970 35232 26976 35244
rect 27028 35232 27034 35284
rect 28077 35275 28135 35281
rect 28077 35241 28089 35275
rect 28123 35272 28135 35275
rect 28166 35272 28172 35284
rect 28123 35244 28172 35272
rect 28123 35241 28135 35244
rect 28077 35235 28135 35241
rect 28166 35232 28172 35244
rect 28224 35232 28230 35284
rect 28258 35232 28264 35284
rect 28316 35272 28322 35284
rect 28316 35244 29684 35272
rect 28316 35232 28322 35244
rect 15105 35139 15163 35145
rect 12820 35108 13492 35136
rect 11514 35028 11520 35080
rect 11572 35068 11578 35080
rect 11793 35071 11851 35077
rect 11793 35068 11805 35071
rect 11572 35040 11805 35068
rect 11572 35028 11578 35040
rect 11793 35037 11805 35040
rect 11839 35037 11851 35071
rect 11974 35068 11980 35080
rect 11935 35040 11980 35068
rect 11793 35031 11851 35037
rect 11974 35028 11980 35040
rect 12032 35028 12038 35080
rect 12434 35028 12440 35080
rect 12492 35068 12498 35080
rect 12713 35071 12771 35077
rect 12713 35068 12725 35071
rect 12492 35040 12725 35068
rect 12492 35028 12498 35040
rect 12713 35037 12725 35040
rect 12759 35037 12771 35071
rect 12713 35031 12771 35037
rect 12802 35028 12808 35080
rect 12860 35068 12866 35080
rect 13464 35077 13492 35108
rect 13556 35108 14412 35136
rect 13556 35080 13584 35108
rect 13449 35071 13507 35077
rect 12860 35040 12905 35068
rect 12860 35028 12866 35040
rect 13449 35037 13461 35071
rect 13495 35037 13507 35071
rect 13449 35031 13507 35037
rect 2004 34972 6914 35000
rect 11885 35003 11943 35009
rect 2004 34960 2010 34972
rect 11885 34969 11897 35003
rect 11931 35000 11943 35003
rect 12529 35003 12587 35009
rect 12529 35000 12541 35003
rect 11931 34972 12541 35000
rect 11931 34969 11943 34972
rect 11885 34963 11943 34969
rect 12529 34969 12541 34972
rect 12575 34969 12587 35003
rect 13262 35000 13268 35012
rect 13223 34972 13268 35000
rect 12529 34963 12587 34969
rect 12544 34932 12572 34963
rect 13262 34960 13268 34972
rect 13320 34960 13326 35012
rect 13464 35000 13492 35031
rect 13538 35028 13544 35080
rect 13596 35068 13602 35080
rect 14384 35077 14412 35108
rect 15105 35105 15117 35139
rect 15151 35136 15163 35139
rect 15838 35136 15844 35148
rect 15151 35108 15844 35136
rect 15151 35105 15163 35108
rect 15105 35099 15163 35105
rect 15838 35096 15844 35108
rect 15896 35136 15902 35148
rect 17034 35136 17040 35148
rect 15896 35108 17040 35136
rect 15896 35096 15902 35108
rect 14093 35071 14151 35077
rect 13596 35040 13641 35068
rect 13596 35028 13602 35040
rect 14093 35037 14105 35071
rect 14139 35068 14151 35071
rect 14369 35071 14427 35077
rect 14139 35040 14320 35068
rect 14139 35037 14151 35040
rect 14093 35031 14151 35037
rect 14185 35003 14243 35009
rect 14185 35000 14197 35003
rect 13464 34972 14197 35000
rect 14185 34969 14197 34972
rect 14231 34969 14243 35003
rect 14185 34963 14243 34969
rect 12710 34932 12716 34944
rect 12544 34904 12716 34932
rect 12710 34892 12716 34904
rect 12768 34892 12774 34944
rect 13280 34932 13308 34960
rect 14292 34932 14320 35040
rect 14369 35037 14381 35071
rect 14415 35037 14427 35071
rect 15562 35068 15568 35080
rect 15523 35040 15568 35068
rect 14369 35031 14427 35037
rect 15562 35028 15568 35040
rect 15620 35028 15626 35080
rect 16224 35077 16252 35108
rect 17034 35096 17040 35108
rect 17092 35096 17098 35148
rect 18248 35145 18276 35232
rect 19904 35204 19932 35232
rect 22554 35204 22560 35216
rect 18340 35176 19932 35204
rect 20088 35176 22560 35204
rect 17405 35139 17463 35145
rect 17405 35105 17417 35139
rect 17451 35136 17463 35139
rect 18233 35139 18291 35145
rect 17451 35108 17724 35136
rect 17451 35105 17463 35108
rect 17405 35099 17463 35105
rect 16209 35071 16267 35077
rect 16209 35037 16221 35071
rect 16255 35037 16267 35071
rect 16209 35031 16267 35037
rect 16301 35071 16359 35077
rect 16301 35037 16313 35071
rect 16347 35037 16359 35071
rect 16301 35031 16359 35037
rect 16316 35000 16344 35031
rect 16666 35028 16672 35080
rect 16724 35068 16730 35080
rect 17126 35068 17132 35080
rect 16724 35040 17132 35068
rect 16724 35028 16730 35040
rect 17126 35028 17132 35040
rect 17184 35068 17190 35080
rect 17589 35071 17647 35077
rect 17589 35068 17601 35071
rect 17184 35040 17601 35068
rect 17184 35028 17190 35040
rect 17589 35037 17601 35040
rect 17635 35037 17647 35071
rect 17696 35068 17724 35108
rect 18233 35105 18245 35139
rect 18279 35105 18291 35139
rect 18233 35099 18291 35105
rect 18138 35068 18144 35080
rect 17696 35040 18144 35068
rect 17589 35031 17647 35037
rect 14568 34972 16344 35000
rect 17604 35000 17632 35031
rect 18138 35028 18144 35040
rect 18196 35068 18202 35080
rect 18340 35068 18368 35176
rect 19889 35139 19947 35145
rect 19889 35105 19901 35139
rect 19935 35136 19947 35139
rect 19978 35136 19984 35148
rect 19935 35108 19984 35136
rect 19935 35105 19947 35108
rect 19889 35099 19947 35105
rect 19978 35096 19984 35108
rect 20036 35096 20042 35148
rect 20088 35145 20116 35176
rect 22554 35164 22560 35176
rect 22612 35204 22618 35216
rect 24489 35207 24547 35213
rect 24489 35204 24501 35207
rect 22612 35176 24501 35204
rect 22612 35164 22618 35176
rect 24489 35173 24501 35176
rect 24535 35173 24547 35207
rect 24489 35167 24547 35173
rect 25317 35207 25375 35213
rect 25317 35173 25329 35207
rect 25363 35204 25375 35207
rect 25363 35176 26188 35204
rect 25363 35173 25375 35176
rect 25317 35167 25375 35173
rect 20073 35139 20131 35145
rect 20073 35105 20085 35139
rect 20119 35105 20131 35139
rect 20073 35099 20131 35105
rect 20809 35139 20867 35145
rect 20809 35105 20821 35139
rect 20855 35136 20867 35139
rect 21082 35136 21088 35148
rect 20855 35108 21088 35136
rect 20855 35105 20867 35108
rect 20809 35099 20867 35105
rect 21082 35096 21088 35108
rect 21140 35096 21146 35148
rect 21450 35096 21456 35148
rect 21508 35136 21514 35148
rect 21821 35139 21879 35145
rect 21821 35136 21833 35139
rect 21508 35108 21833 35136
rect 21508 35096 21514 35108
rect 21821 35105 21833 35108
rect 21867 35105 21879 35139
rect 22738 35136 22744 35148
rect 22699 35108 22744 35136
rect 21821 35099 21879 35105
rect 22738 35096 22744 35108
rect 22796 35096 22802 35148
rect 23014 35136 23020 35148
rect 22975 35108 23020 35136
rect 23014 35096 23020 35108
rect 23072 35096 23078 35148
rect 23845 35139 23903 35145
rect 23845 35105 23857 35139
rect 23891 35136 23903 35139
rect 23891 35108 25084 35136
rect 23891 35105 23903 35108
rect 23845 35099 23903 35105
rect 18506 35068 18512 35080
rect 18196 35040 18368 35068
rect 18467 35040 18512 35068
rect 18196 35028 18202 35040
rect 18506 35028 18512 35040
rect 18564 35028 18570 35080
rect 19794 35068 19800 35080
rect 19755 35040 19800 35068
rect 19794 35028 19800 35040
rect 19852 35028 19858 35080
rect 20714 35068 20720 35080
rect 20675 35040 20720 35068
rect 20714 35028 20720 35040
rect 20772 35028 20778 35080
rect 21542 35068 21548 35080
rect 21503 35040 21548 35068
rect 21542 35028 21548 35040
rect 21600 35028 21606 35080
rect 21634 35028 21640 35080
rect 21692 35068 21698 35080
rect 22373 35071 22431 35077
rect 22373 35068 22385 35071
rect 21692 35040 21737 35068
rect 22066 35040 22385 35068
rect 21692 35028 21698 35040
rect 19426 35000 19432 35012
rect 17604 34972 19432 35000
rect 14568 34944 14596 34972
rect 19426 34960 19432 34972
rect 19484 34960 19490 35012
rect 19812 35000 19840 35028
rect 20070 35000 20076 35012
rect 19812 34972 20076 35000
rect 20070 34960 20076 34972
rect 20128 34960 20134 35012
rect 21821 35003 21879 35009
rect 21821 34969 21833 35003
rect 21867 35000 21879 35003
rect 22066 35000 22094 35040
rect 22373 35037 22385 35040
rect 22419 35037 22431 35071
rect 22554 35068 22560 35080
rect 22515 35040 22560 35068
rect 22373 35031 22431 35037
rect 22554 35028 22560 35040
rect 22612 35028 22618 35080
rect 23106 35068 23112 35080
rect 23067 35040 23112 35068
rect 23106 35028 23112 35040
rect 23164 35028 23170 35080
rect 24486 35068 24492 35080
rect 24447 35040 24492 35068
rect 24486 35028 24492 35040
rect 24544 35028 24550 35080
rect 24673 35071 24731 35077
rect 24673 35037 24685 35071
rect 24719 35068 24731 35071
rect 24946 35068 24952 35080
rect 24719 35040 24952 35068
rect 24719 35037 24731 35040
rect 24673 35031 24731 35037
rect 24946 35028 24952 35040
rect 25004 35028 25010 35080
rect 25056 35068 25084 35108
rect 25130 35096 25136 35148
rect 25188 35136 25194 35148
rect 25501 35139 25559 35145
rect 25501 35136 25513 35139
rect 25188 35108 25513 35136
rect 25188 35096 25194 35108
rect 25501 35105 25513 35108
rect 25547 35105 25559 35139
rect 25501 35099 25559 35105
rect 26160 35080 26188 35176
rect 27706 35164 27712 35216
rect 27764 35204 27770 35216
rect 29656 35213 29684 35244
rect 30282 35232 30288 35284
rect 30340 35272 30346 35284
rect 30377 35275 30435 35281
rect 30377 35272 30389 35275
rect 30340 35244 30389 35272
rect 30340 35232 30346 35244
rect 30377 35241 30389 35244
rect 30423 35241 30435 35275
rect 30377 35235 30435 35241
rect 30834 35232 30840 35284
rect 30892 35272 30898 35284
rect 31294 35272 31300 35284
rect 30892 35244 31300 35272
rect 30892 35232 30898 35244
rect 31294 35232 31300 35244
rect 31352 35232 31358 35284
rect 32030 35232 32036 35284
rect 32088 35272 32094 35284
rect 32493 35275 32551 35281
rect 32493 35272 32505 35275
rect 32088 35244 32505 35272
rect 32088 35232 32094 35244
rect 32493 35241 32505 35244
rect 32539 35241 32551 35275
rect 33226 35272 33232 35284
rect 33187 35244 33232 35272
rect 32493 35235 32551 35241
rect 33226 35232 33232 35244
rect 33284 35232 33290 35284
rect 33502 35232 33508 35284
rect 33560 35272 33566 35284
rect 34885 35275 34943 35281
rect 34885 35272 34897 35275
rect 33560 35244 34897 35272
rect 33560 35232 33566 35244
rect 34885 35241 34897 35244
rect 34931 35241 34943 35275
rect 39945 35275 40003 35281
rect 39945 35272 39957 35275
rect 34885 35235 34943 35241
rect 38764 35244 39957 35272
rect 29641 35207 29699 35213
rect 27764 35176 29592 35204
rect 27764 35164 27770 35176
rect 29012 35145 29040 35176
rect 28993 35139 29051 35145
rect 28736 35108 28948 35136
rect 25225 35071 25283 35077
rect 25225 35068 25237 35071
rect 25056 35040 25237 35068
rect 25225 35037 25237 35040
rect 25271 35068 25283 35071
rect 25961 35071 26019 35077
rect 25961 35068 25973 35071
rect 25271 35040 25973 35068
rect 25271 35037 25283 35040
rect 25225 35031 25283 35037
rect 25961 35037 25973 35040
rect 26007 35037 26019 35071
rect 26142 35068 26148 35080
rect 26103 35040 26148 35068
rect 25961 35031 26019 35037
rect 24854 35000 24860 35012
rect 21867 34972 22094 35000
rect 23676 34972 24860 35000
rect 21867 34969 21879 34972
rect 21821 34963 21879 34969
rect 14550 34932 14556 34944
rect 13280 34904 14320 34932
rect 14511 34904 14556 34932
rect 14550 34892 14556 34904
rect 14608 34892 14614 34944
rect 15378 34892 15384 34944
rect 15436 34932 15442 34944
rect 15473 34935 15531 34941
rect 15473 34932 15485 34935
rect 15436 34904 15485 34932
rect 15436 34892 15442 34904
rect 15473 34901 15485 34904
rect 15519 34932 15531 34935
rect 15930 34932 15936 34944
rect 15519 34904 15936 34932
rect 15519 34901 15531 34904
rect 15473 34895 15531 34901
rect 15930 34892 15936 34904
rect 15988 34932 15994 34944
rect 16025 34935 16083 34941
rect 16025 34932 16037 34935
rect 15988 34904 16037 34932
rect 15988 34892 15994 34904
rect 16025 34901 16037 34904
rect 16071 34901 16083 34935
rect 16025 34895 16083 34901
rect 16945 34935 17003 34941
rect 16945 34901 16957 34935
rect 16991 34932 17003 34935
rect 18046 34932 18052 34944
rect 16991 34904 18052 34932
rect 16991 34901 17003 34904
rect 16945 34895 17003 34901
rect 18046 34892 18052 34904
rect 18104 34932 18110 34944
rect 18782 34932 18788 34944
rect 18104 34904 18788 34932
rect 18104 34892 18110 34904
rect 18782 34892 18788 34904
rect 18840 34892 18846 34944
rect 19334 34892 19340 34944
rect 19392 34932 19398 34944
rect 23676 34932 23704 34972
rect 24854 34960 24860 34972
rect 24912 34960 24918 35012
rect 25866 34960 25872 35012
rect 25924 35000 25930 35012
rect 25976 35000 26004 35031
rect 26142 35028 26148 35040
rect 26200 35028 26206 35080
rect 26234 35028 26240 35080
rect 26292 35068 26298 35080
rect 26329 35071 26387 35077
rect 26329 35068 26341 35071
rect 26292 35040 26341 35068
rect 26292 35028 26298 35040
rect 26329 35037 26341 35040
rect 26375 35068 26387 35071
rect 26973 35071 27031 35077
rect 26973 35068 26985 35071
rect 26375 35040 26985 35068
rect 26375 35037 26387 35040
rect 26329 35031 26387 35037
rect 26973 35037 26985 35040
rect 27019 35068 27031 35071
rect 27062 35068 27068 35080
rect 27019 35040 27068 35068
rect 27019 35037 27031 35040
rect 26973 35031 27031 35037
rect 26786 35000 26792 35012
rect 25924 34972 26792 35000
rect 25924 34960 25930 34972
rect 26786 34960 26792 34972
rect 26844 34960 26850 35012
rect 26988 35000 27016 35031
rect 27062 35028 27068 35040
rect 27120 35028 27126 35080
rect 27246 35068 27252 35080
rect 27207 35040 27252 35068
rect 27246 35028 27252 35040
rect 27304 35028 27310 35080
rect 28258 35068 28264 35080
rect 27908 35040 28264 35068
rect 26988 34972 27568 35000
rect 19392 34904 23704 34932
rect 25501 34935 25559 34941
rect 19392 34892 19398 34904
rect 25501 34901 25513 34935
rect 25547 34932 25559 34935
rect 26050 34932 26056 34944
rect 25547 34904 26056 34932
rect 25547 34901 25559 34904
rect 25501 34895 25559 34901
rect 26050 34892 26056 34904
rect 26108 34892 26114 34944
rect 27065 34935 27123 34941
rect 27065 34901 27077 34935
rect 27111 34932 27123 34935
rect 27246 34932 27252 34944
rect 27111 34904 27252 34932
rect 27111 34901 27123 34904
rect 27065 34895 27123 34901
rect 27246 34892 27252 34904
rect 27304 34892 27310 34944
rect 27338 34892 27344 34944
rect 27396 34932 27402 34944
rect 27433 34935 27491 34941
rect 27433 34932 27445 34935
rect 27396 34904 27445 34932
rect 27396 34892 27402 34904
rect 27433 34901 27445 34904
rect 27479 34901 27491 34935
rect 27540 34932 27568 34972
rect 27614 34960 27620 35012
rect 27672 35000 27678 35012
rect 27908 35009 27936 35040
rect 28258 35028 28264 35040
rect 28316 35028 28322 35080
rect 28736 35077 28764 35108
rect 28721 35071 28779 35077
rect 28721 35037 28733 35071
rect 28767 35037 28779 35071
rect 28721 35031 28779 35037
rect 28813 35071 28871 35077
rect 28813 35037 28825 35071
rect 28859 35037 28871 35071
rect 28920 35068 28948 35108
rect 28993 35105 29005 35139
rect 29039 35105 29051 35139
rect 29564 35136 29592 35176
rect 29641 35173 29653 35207
rect 29687 35204 29699 35207
rect 31570 35204 31576 35216
rect 29687 35176 31576 35204
rect 29687 35173 29699 35176
rect 29641 35167 29699 35173
rect 31570 35164 31576 35176
rect 31628 35164 31634 35216
rect 33594 35164 33600 35216
rect 33652 35204 33658 35216
rect 36538 35204 36544 35216
rect 33652 35176 35020 35204
rect 36499 35176 36544 35204
rect 33652 35164 33658 35176
rect 30834 35136 30840 35148
rect 29564 35108 30840 35136
rect 28993 35099 29051 35105
rect 30834 35096 30840 35108
rect 30892 35096 30898 35148
rect 31938 35136 31944 35148
rect 30944 35108 31944 35136
rect 29914 35068 29920 35080
rect 28920 35040 29920 35068
rect 28813 35031 28871 35037
rect 27893 35003 27951 35009
rect 27893 35000 27905 35003
rect 27672 34972 27905 35000
rect 27672 34960 27678 34972
rect 27893 34969 27905 34972
rect 27939 34969 27951 35003
rect 28828 35000 28856 35031
rect 29914 35028 29920 35040
rect 29972 35028 29978 35080
rect 30558 35077 30564 35080
rect 30556 35068 30564 35077
rect 30519 35040 30564 35068
rect 30556 35031 30564 35040
rect 30558 35028 30564 35031
rect 30616 35028 30622 35080
rect 30944 35077 30972 35108
rect 31938 35096 31944 35108
rect 31996 35096 32002 35148
rect 33689 35139 33747 35145
rect 33689 35105 33701 35139
rect 33735 35136 33747 35139
rect 34146 35136 34152 35148
rect 33735 35108 34152 35136
rect 33735 35105 33747 35108
rect 33689 35099 33747 35105
rect 34146 35096 34152 35108
rect 34204 35096 34210 35148
rect 34698 35136 34704 35148
rect 34659 35108 34704 35136
rect 34698 35096 34704 35108
rect 34756 35096 34762 35148
rect 30928 35071 30986 35077
rect 30928 35037 30940 35071
rect 30974 35037 30986 35071
rect 30928 35031 30986 35037
rect 31021 35071 31079 35077
rect 31021 35037 31033 35071
rect 31067 35068 31079 35071
rect 32030 35068 32036 35080
rect 31067 35040 32036 35068
rect 31067 35037 31079 35040
rect 31021 35031 31079 35037
rect 32030 35028 32036 35040
rect 32088 35028 32094 35080
rect 33410 35068 33416 35080
rect 33371 35040 33416 35068
rect 33410 35028 33416 35040
rect 33468 35028 33474 35080
rect 33505 35071 33563 35077
rect 33505 35037 33517 35071
rect 33551 35037 33563 35071
rect 33778 35068 33784 35080
rect 33739 35040 33784 35068
rect 33505 35031 33563 35037
rect 27893 34963 27951 34969
rect 28276 34972 28856 35000
rect 28276 34944 28304 34972
rect 30466 34960 30472 35012
rect 30524 35000 30530 35012
rect 30653 35003 30711 35009
rect 30653 35000 30665 35003
rect 30524 34972 30665 35000
rect 30524 34960 30530 34972
rect 30653 34969 30665 34972
rect 30699 34969 30711 35003
rect 30653 34963 30711 34969
rect 28093 34935 28151 34941
rect 28093 34932 28105 34935
rect 27540 34904 28105 34932
rect 27433 34895 27491 34901
rect 28093 34901 28105 34904
rect 28139 34901 28151 34935
rect 28258 34932 28264 34944
rect 28219 34904 28264 34932
rect 28093 34895 28151 34901
rect 28258 34892 28264 34904
rect 28316 34892 28322 34944
rect 28902 34892 28908 34944
rect 28960 34932 28966 34944
rect 28997 34935 29055 34941
rect 28997 34932 29009 34935
rect 28960 34904 29009 34932
rect 28960 34892 28966 34904
rect 28997 34901 29009 34904
rect 29043 34901 29055 34935
rect 30668 34932 30696 34963
rect 30742 34960 30748 35012
rect 30800 35000 30806 35012
rect 31481 35003 31539 35009
rect 30800 34972 30845 35000
rect 30800 34960 30806 34972
rect 31481 34969 31493 35003
rect 31527 34969 31539 35003
rect 31481 34963 31539 34969
rect 31665 35003 31723 35009
rect 31665 34969 31677 35003
rect 31711 34969 31723 35003
rect 31665 34963 31723 34969
rect 31849 35003 31907 35009
rect 31849 34969 31861 35003
rect 31895 35000 31907 35003
rect 31938 35000 31944 35012
rect 31895 34972 31944 35000
rect 31895 34969 31907 34972
rect 31849 34963 31907 34969
rect 31496 34932 31524 34963
rect 30668 34904 31524 34932
rect 31680 34932 31708 34963
rect 31938 34960 31944 34972
rect 31996 35000 32002 35012
rect 32122 35000 32128 35012
rect 31996 34972 32128 35000
rect 31996 34960 32002 34972
rect 32122 34960 32128 34972
rect 32180 34960 32186 35012
rect 32398 35000 32404 35012
rect 32359 34972 32404 35000
rect 32398 34960 32404 34972
rect 32456 34960 32462 35012
rect 33520 35000 33548 35031
rect 33778 35028 33784 35040
rect 33836 35028 33842 35080
rect 34882 35028 34888 35080
rect 34940 35068 34946 35080
rect 34992 35077 35020 35176
rect 36538 35164 36544 35176
rect 36596 35164 36602 35216
rect 38102 35164 38108 35216
rect 38160 35204 38166 35216
rect 38562 35204 38568 35216
rect 38160 35176 38568 35204
rect 38160 35164 38166 35176
rect 38562 35164 38568 35176
rect 38620 35164 38626 35216
rect 36262 35136 36268 35148
rect 36223 35108 36268 35136
rect 36262 35096 36268 35108
rect 36320 35096 36326 35148
rect 34977 35071 35035 35077
rect 34977 35068 34989 35071
rect 34940 35040 34989 35068
rect 34940 35028 34946 35040
rect 34977 35037 34989 35040
rect 35023 35037 35035 35071
rect 34977 35031 35035 35037
rect 36173 35071 36231 35077
rect 36173 35037 36185 35071
rect 36219 35068 36231 35071
rect 37366 35068 37372 35080
rect 36219 35040 37372 35068
rect 36219 35037 36231 35040
rect 36173 35031 36231 35037
rect 37366 35028 37372 35040
rect 37424 35028 37430 35080
rect 37918 35068 37924 35080
rect 37879 35040 37924 35068
rect 37918 35028 37924 35040
rect 37976 35028 37982 35080
rect 38105 35071 38163 35077
rect 38105 35037 38117 35071
rect 38151 35068 38163 35071
rect 38194 35068 38200 35080
rect 38151 35040 38200 35068
rect 38151 35037 38163 35040
rect 38105 35031 38163 35037
rect 38194 35028 38200 35040
rect 38252 35068 38258 35080
rect 38764 35077 38792 35244
rect 39945 35241 39957 35244
rect 39991 35241 40003 35275
rect 41506 35272 41512 35284
rect 41467 35244 41512 35272
rect 39945 35235 40003 35241
rect 41506 35232 41512 35244
rect 41564 35232 41570 35284
rect 42613 35275 42671 35281
rect 42613 35241 42625 35275
rect 42659 35272 42671 35275
rect 43530 35272 43536 35284
rect 42659 35244 43536 35272
rect 42659 35241 42671 35244
rect 42613 35235 42671 35241
rect 38838 35164 38844 35216
rect 38896 35204 38902 35216
rect 42628 35204 42656 35235
rect 43530 35232 43536 35244
rect 43588 35232 43594 35284
rect 38896 35176 42656 35204
rect 38896 35164 38902 35176
rect 40126 35136 40132 35148
rect 40087 35108 40132 35136
rect 40126 35096 40132 35108
rect 40184 35096 40190 35148
rect 38749 35071 38807 35077
rect 38749 35068 38761 35071
rect 38252 35040 38761 35068
rect 38252 35028 38258 35040
rect 38749 35037 38761 35040
rect 38795 35037 38807 35071
rect 38749 35031 38807 35037
rect 39758 35028 39764 35080
rect 39816 35068 39822 35080
rect 40221 35071 40279 35077
rect 40221 35068 40233 35071
rect 39816 35040 40233 35068
rect 39816 35028 39822 35040
rect 40221 35037 40233 35040
rect 40267 35068 40279 35071
rect 40862 35068 40868 35080
rect 40267 35040 40868 35068
rect 40267 35037 40279 35040
rect 40221 35031 40279 35037
rect 40862 35028 40868 35040
rect 40920 35028 40926 35080
rect 40957 35071 41015 35077
rect 40957 35037 40969 35071
rect 41003 35068 41015 35071
rect 41414 35068 41420 35080
rect 41003 35040 41420 35068
rect 41003 35037 41015 35040
rect 40957 35031 41015 35037
rect 34701 35003 34759 35009
rect 34701 35000 34713 35003
rect 33520 34972 34713 35000
rect 34701 34969 34713 34972
rect 34747 34969 34759 35003
rect 34701 34963 34759 34969
rect 38013 35003 38071 35009
rect 38013 34969 38025 35003
rect 38059 35000 38071 35003
rect 39114 35000 39120 35012
rect 38059 34972 39120 35000
rect 38059 34969 38071 34972
rect 38013 34963 38071 34969
rect 39114 34960 39120 34972
rect 39172 34960 39178 35012
rect 39942 34960 39948 35012
rect 40000 35000 40006 35012
rect 40972 35000 41000 35031
rect 41414 35028 41420 35040
rect 41472 35068 41478 35080
rect 41966 35068 41972 35080
rect 41472 35040 41972 35068
rect 41472 35028 41478 35040
rect 41966 35028 41972 35040
rect 42024 35028 42030 35080
rect 40000 34972 41000 35000
rect 40000 34960 40006 34972
rect 41506 34960 41512 35012
rect 41564 35000 41570 35012
rect 41874 35000 41880 35012
rect 41564 34972 41880 35000
rect 41564 34960 41570 34972
rect 41874 34960 41880 34972
rect 41932 35000 41938 35012
rect 42061 35003 42119 35009
rect 42061 35000 42073 35003
rect 41932 34972 42073 35000
rect 41932 34960 41938 34972
rect 42061 34969 42073 34972
rect 42107 34969 42119 35003
rect 42061 34963 42119 34969
rect 31754 34932 31760 34944
rect 31680 34904 31760 34932
rect 28997 34895 29055 34901
rect 31754 34892 31760 34904
rect 31812 34932 31818 34944
rect 32416 34932 32444 34960
rect 31812 34904 32444 34932
rect 31812 34892 31818 34904
rect 34514 34892 34520 34944
rect 34572 34932 34578 34944
rect 35437 34935 35495 34941
rect 35437 34932 35449 34935
rect 34572 34904 35449 34932
rect 34572 34892 34578 34904
rect 35437 34901 35449 34904
rect 35483 34901 35495 34935
rect 36998 34932 37004 34944
rect 36959 34904 37004 34932
rect 35437 34895 35495 34901
rect 36998 34892 37004 34904
rect 37056 34892 37062 34944
rect 38102 34892 38108 34944
rect 38160 34932 38166 34944
rect 38657 34935 38715 34941
rect 38657 34932 38669 34935
rect 38160 34904 38669 34932
rect 38160 34892 38166 34904
rect 38657 34901 38669 34904
rect 38703 34901 38715 34935
rect 39298 34932 39304 34944
rect 39211 34904 39304 34932
rect 38657 34895 38715 34901
rect 39298 34892 39304 34904
rect 39356 34932 39362 34944
rect 39758 34932 39764 34944
rect 39356 34904 39764 34932
rect 39356 34892 39362 34904
rect 39758 34892 39764 34904
rect 39816 34932 39822 34944
rect 41690 34932 41696 34944
rect 39816 34904 41696 34932
rect 39816 34892 39822 34904
rect 41690 34892 41696 34904
rect 41748 34892 41754 34944
rect 43070 34932 43076 34944
rect 43031 34904 43076 34932
rect 43070 34892 43076 34904
rect 43128 34892 43134 34944
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 1946 34728 1952 34740
rect 1907 34700 1952 34728
rect 1946 34688 1952 34700
rect 2004 34688 2010 34740
rect 9122 34728 9128 34740
rect 9083 34700 9128 34728
rect 9122 34688 9128 34700
rect 9180 34688 9186 34740
rect 10226 34728 10232 34740
rect 10187 34700 10232 34728
rect 10226 34688 10232 34700
rect 10284 34688 10290 34740
rect 10965 34731 11023 34737
rect 10965 34697 10977 34731
rect 11011 34728 11023 34731
rect 11974 34728 11980 34740
rect 11011 34700 11980 34728
rect 11011 34697 11023 34700
rect 10965 34691 11023 34697
rect 11974 34688 11980 34700
rect 12032 34688 12038 34740
rect 12066 34688 12072 34740
rect 12124 34728 12130 34740
rect 12529 34731 12587 34737
rect 12529 34728 12541 34731
rect 12124 34700 12541 34728
rect 12124 34688 12130 34700
rect 12529 34697 12541 34700
rect 12575 34728 12587 34731
rect 12802 34728 12808 34740
rect 12575 34700 12808 34728
rect 12575 34697 12587 34700
rect 12529 34691 12587 34697
rect 12802 34688 12808 34700
rect 12860 34688 12866 34740
rect 12897 34731 12955 34737
rect 12897 34697 12909 34731
rect 12943 34728 12955 34731
rect 13262 34728 13268 34740
rect 12943 34700 13268 34728
rect 12943 34697 12955 34700
rect 12897 34691 12955 34697
rect 13262 34688 13268 34700
rect 13320 34688 13326 34740
rect 14550 34688 14556 34740
rect 14608 34728 14614 34740
rect 15565 34731 15623 34737
rect 15565 34728 15577 34731
rect 14608 34700 15577 34728
rect 14608 34688 14614 34700
rect 15565 34697 15577 34700
rect 15611 34697 15623 34731
rect 15565 34691 15623 34697
rect 15654 34688 15660 34740
rect 15712 34728 15718 34740
rect 15749 34731 15807 34737
rect 15749 34728 15761 34731
rect 15712 34700 15761 34728
rect 15712 34688 15718 34700
rect 15749 34697 15761 34700
rect 15795 34697 15807 34731
rect 15749 34691 15807 34697
rect 16850 34688 16856 34740
rect 16908 34728 16914 34740
rect 18065 34731 18123 34737
rect 18065 34728 18077 34731
rect 16908 34700 18077 34728
rect 16908 34688 16914 34700
rect 18065 34697 18077 34700
rect 18111 34697 18123 34731
rect 18065 34691 18123 34697
rect 18233 34731 18291 34737
rect 18233 34697 18245 34731
rect 18279 34728 18291 34731
rect 19334 34728 19340 34740
rect 18279 34700 19340 34728
rect 18279 34697 18291 34700
rect 18233 34691 18291 34697
rect 19334 34688 19340 34700
rect 19392 34688 19398 34740
rect 19705 34731 19763 34737
rect 19705 34697 19717 34731
rect 19751 34728 19763 34731
rect 19978 34728 19984 34740
rect 19751 34700 19984 34728
rect 19751 34697 19763 34700
rect 19705 34691 19763 34697
rect 19978 34688 19984 34700
rect 20036 34688 20042 34740
rect 21177 34731 21235 34737
rect 21177 34697 21189 34731
rect 21223 34728 21235 34731
rect 21634 34728 21640 34740
rect 21223 34700 21640 34728
rect 21223 34697 21235 34700
rect 21177 34691 21235 34697
rect 21634 34688 21640 34700
rect 21692 34688 21698 34740
rect 23106 34728 23112 34740
rect 23067 34700 23112 34728
rect 23106 34688 23112 34700
rect 23164 34688 23170 34740
rect 24397 34731 24455 34737
rect 24397 34697 24409 34731
rect 24443 34728 24455 34731
rect 24670 34728 24676 34740
rect 24443 34700 24676 34728
rect 24443 34697 24455 34700
rect 24397 34691 24455 34697
rect 24670 34688 24676 34700
rect 24728 34688 24734 34740
rect 25038 34688 25044 34740
rect 25096 34688 25102 34740
rect 26142 34688 26148 34740
rect 26200 34728 26206 34740
rect 30377 34731 30435 34737
rect 26200 34700 27384 34728
rect 26200 34688 26206 34700
rect 1578 34552 1584 34604
rect 1636 34592 1642 34604
rect 1857 34595 1915 34601
rect 1857 34592 1869 34595
rect 1636 34564 1869 34592
rect 1636 34552 1642 34564
rect 1857 34561 1869 34564
rect 1903 34561 1915 34595
rect 9140 34592 9168 34688
rect 11517 34663 11575 34669
rect 11517 34660 11529 34663
rect 10796 34632 11529 34660
rect 10796 34601 10824 34632
rect 11517 34629 11529 34632
rect 11563 34629 11575 34663
rect 11517 34623 11575 34629
rect 12618 34620 12624 34672
rect 12676 34660 12682 34672
rect 14921 34663 14979 34669
rect 12676 34632 14872 34660
rect 12676 34620 12682 34632
rect 10781 34595 10839 34601
rect 10781 34592 10793 34595
rect 9140 34564 10793 34592
rect 1857 34555 1915 34561
rect 10781 34561 10793 34564
rect 10827 34561 10839 34595
rect 10781 34555 10839 34561
rect 10965 34595 11023 34601
rect 10965 34561 10977 34595
rect 11011 34592 11023 34595
rect 11701 34595 11759 34601
rect 11701 34592 11713 34595
rect 11011 34564 11713 34592
rect 11011 34561 11023 34564
rect 10965 34555 11023 34561
rect 11701 34561 11713 34564
rect 11747 34561 11759 34595
rect 11701 34555 11759 34561
rect 10318 34524 10324 34536
rect 9784 34496 10324 34524
rect 9784 34400 9812 34496
rect 10318 34484 10324 34496
rect 10376 34524 10382 34536
rect 10980 34524 11008 34555
rect 12434 34552 12440 34604
rect 12492 34592 12498 34604
rect 12710 34592 12716 34604
rect 12492 34564 12537 34592
rect 12671 34564 12716 34592
rect 12492 34552 12498 34564
rect 12710 34552 12716 34564
rect 12768 34552 12774 34604
rect 13814 34592 13820 34604
rect 13775 34564 13820 34592
rect 13814 34552 13820 34564
rect 13872 34552 13878 34604
rect 13909 34595 13967 34601
rect 13909 34561 13921 34595
rect 13955 34561 13967 34595
rect 13909 34555 13967 34561
rect 14093 34595 14151 34601
rect 14093 34561 14105 34595
rect 14139 34592 14151 34595
rect 14139 34564 14412 34592
rect 14139 34561 14151 34564
rect 14093 34555 14151 34561
rect 13924 34524 13952 34555
rect 14274 34524 14280 34536
rect 10376 34496 11008 34524
rect 11072 34496 14280 34524
rect 10376 34484 10382 34496
rect 10226 34416 10232 34468
rect 10284 34456 10290 34468
rect 11072 34456 11100 34496
rect 14274 34484 14280 34496
rect 14332 34484 14338 34536
rect 14384 34524 14412 34564
rect 14458 34552 14464 34604
rect 14516 34592 14522 34604
rect 14553 34595 14611 34601
rect 14553 34592 14565 34595
rect 14516 34564 14565 34592
rect 14516 34552 14522 34564
rect 14553 34561 14565 34564
rect 14599 34561 14611 34595
rect 14734 34592 14740 34604
rect 14695 34564 14740 34592
rect 14553 34555 14611 34561
rect 14734 34552 14740 34564
rect 14792 34552 14798 34604
rect 14844 34592 14872 34632
rect 14921 34629 14933 34663
rect 14967 34660 14979 34663
rect 16574 34660 16580 34672
rect 14967 34632 16580 34660
rect 14967 34629 14979 34632
rect 14921 34623 14979 34629
rect 16574 34620 16580 34632
rect 16632 34660 16638 34672
rect 17865 34663 17923 34669
rect 16632 34632 16896 34660
rect 16632 34620 16638 34632
rect 15657 34595 15715 34601
rect 14844 34564 15424 34592
rect 15286 34524 15292 34536
rect 14384 34496 15292 34524
rect 15286 34484 15292 34496
rect 15344 34484 15350 34536
rect 15396 34524 15424 34564
rect 15657 34561 15669 34595
rect 15703 34592 15715 34595
rect 15838 34592 15844 34604
rect 15703 34564 15844 34592
rect 15703 34561 15715 34564
rect 15657 34555 15715 34561
rect 15838 34552 15844 34564
rect 15896 34552 15902 34604
rect 16868 34601 16896 34632
rect 17865 34629 17877 34663
rect 17911 34660 17923 34663
rect 17954 34660 17960 34672
rect 17911 34632 17960 34660
rect 17911 34629 17923 34632
rect 17865 34623 17923 34629
rect 17954 34620 17960 34632
rect 18012 34620 18018 34672
rect 18782 34660 18788 34672
rect 18743 34632 18788 34660
rect 18782 34620 18788 34632
rect 18840 34620 18846 34672
rect 21266 34660 21272 34672
rect 18892 34632 21272 34660
rect 16853 34595 16911 34601
rect 16853 34561 16865 34595
rect 16899 34561 16911 34595
rect 16853 34555 16911 34561
rect 15933 34527 15991 34533
rect 15396 34496 15884 34524
rect 15378 34456 15384 34468
rect 10284 34428 11100 34456
rect 15339 34428 15384 34456
rect 10284 34416 10290 34428
rect 15378 34416 15384 34428
rect 15436 34416 15442 34468
rect 15856 34456 15884 34496
rect 15933 34493 15945 34527
rect 15979 34524 15991 34527
rect 16666 34524 16672 34536
rect 15979 34496 16672 34524
rect 15979 34493 15991 34496
rect 15933 34487 15991 34493
rect 16666 34484 16672 34496
rect 16724 34484 16730 34536
rect 16758 34484 16764 34536
rect 16816 34524 16822 34536
rect 18892 34524 18920 34632
rect 21266 34620 21272 34632
rect 21324 34620 21330 34672
rect 23474 34660 23480 34672
rect 23435 34632 23480 34660
rect 23474 34620 23480 34632
rect 23532 34620 23538 34672
rect 19242 34592 19248 34604
rect 19203 34564 19248 34592
rect 19242 34552 19248 34564
rect 19300 34552 19306 34604
rect 19334 34552 19340 34604
rect 19392 34592 19398 34604
rect 19521 34595 19579 34601
rect 19392 34564 19437 34592
rect 19392 34552 19398 34564
rect 19521 34561 19533 34595
rect 19567 34561 19579 34595
rect 19521 34555 19579 34561
rect 20993 34595 21051 34601
rect 20993 34561 21005 34595
rect 21039 34592 21051 34595
rect 21082 34592 21088 34604
rect 21039 34564 21088 34592
rect 21039 34561 21051 34564
rect 20993 34555 21051 34561
rect 16816 34496 16861 34524
rect 16960 34496 18920 34524
rect 16816 34484 16822 34496
rect 16960 34456 16988 34496
rect 19426 34484 19432 34536
rect 19484 34524 19490 34536
rect 19536 34524 19564 34555
rect 21082 34552 21088 34564
rect 21140 34552 21146 34604
rect 22281 34595 22339 34601
rect 22281 34561 22293 34595
rect 22327 34592 22339 34595
rect 22370 34592 22376 34604
rect 22327 34564 22376 34592
rect 22327 34561 22339 34564
rect 22281 34555 22339 34561
rect 22370 34552 22376 34564
rect 22428 34552 22434 34604
rect 23247 34595 23305 34601
rect 23247 34592 23259 34595
rect 22664 34564 23259 34592
rect 19484 34496 19564 34524
rect 19484 34484 19490 34496
rect 20714 34484 20720 34536
rect 20772 34524 20778 34536
rect 20809 34527 20867 34533
rect 20809 34524 20821 34527
rect 20772 34496 20821 34524
rect 20772 34484 20778 34496
rect 20809 34493 20821 34496
rect 20855 34493 20867 34527
rect 22186 34524 22192 34536
rect 22147 34496 22192 34524
rect 20809 34487 20867 34493
rect 22186 34484 22192 34496
rect 22244 34484 22250 34536
rect 15856 34428 16988 34456
rect 17221 34459 17279 34465
rect 17221 34425 17233 34459
rect 17267 34456 17279 34459
rect 17310 34456 17316 34468
rect 17267 34428 17316 34456
rect 17267 34425 17279 34428
rect 17221 34419 17279 34425
rect 17310 34416 17316 34428
rect 17368 34416 17374 34468
rect 22664 34465 22692 34564
rect 23247 34561 23259 34564
rect 23293 34561 23305 34595
rect 23247 34555 23305 34561
rect 23385 34595 23443 34601
rect 23385 34561 23397 34595
rect 23431 34592 23443 34595
rect 23658 34592 23664 34604
rect 23431 34564 23520 34592
rect 23619 34564 23664 34592
rect 23431 34561 23443 34564
rect 23385 34555 23443 34561
rect 23492 34536 23520 34564
rect 23658 34552 23664 34564
rect 23716 34552 23722 34604
rect 23753 34595 23811 34601
rect 23753 34561 23765 34595
rect 23799 34592 23811 34595
rect 24026 34592 24032 34604
rect 23799 34564 24032 34592
rect 23799 34561 23811 34564
rect 23753 34555 23811 34561
rect 24026 34552 24032 34564
rect 24084 34552 24090 34604
rect 24210 34592 24216 34604
rect 24171 34564 24216 34592
rect 24210 34552 24216 34564
rect 24268 34552 24274 34604
rect 24397 34595 24455 34601
rect 24397 34561 24409 34595
rect 24443 34592 24455 34595
rect 24762 34592 24768 34604
rect 24443 34564 24768 34592
rect 24443 34561 24455 34564
rect 24397 34555 24455 34561
rect 24762 34552 24768 34564
rect 24820 34552 24826 34604
rect 25056 34601 25084 34688
rect 26329 34663 26387 34669
rect 26329 34660 26341 34663
rect 25332 34632 26341 34660
rect 25041 34595 25099 34601
rect 25041 34561 25053 34595
rect 25087 34561 25099 34595
rect 25222 34592 25228 34604
rect 25183 34564 25228 34592
rect 25041 34555 25099 34561
rect 23474 34484 23480 34536
rect 23532 34484 23538 34536
rect 25056 34524 25084 34555
rect 25222 34552 25228 34564
rect 25280 34552 25286 34604
rect 25332 34601 25360 34632
rect 26329 34629 26341 34632
rect 26375 34629 26387 34663
rect 26329 34623 26387 34629
rect 25317 34595 25375 34601
rect 25317 34561 25329 34595
rect 25363 34561 25375 34595
rect 25774 34592 25780 34604
rect 25735 34564 25780 34592
rect 25317 34555 25375 34561
rect 25774 34552 25780 34564
rect 25832 34552 25838 34604
rect 26050 34592 26056 34604
rect 26011 34564 26056 34592
rect 26050 34552 26056 34564
rect 26108 34552 26114 34604
rect 26145 34595 26203 34601
rect 26145 34561 26157 34595
rect 26191 34592 26203 34595
rect 26234 34592 26240 34604
rect 26191 34564 26240 34592
rect 26191 34561 26203 34564
rect 26145 34555 26203 34561
rect 26234 34552 26240 34564
rect 26292 34552 26298 34604
rect 27154 34592 27160 34604
rect 27115 34564 27160 34592
rect 27154 34552 27160 34564
rect 27212 34552 27218 34604
rect 27356 34601 27384 34700
rect 30377 34697 30389 34731
rect 30423 34728 30435 34731
rect 30742 34728 30748 34740
rect 30423 34700 30748 34728
rect 30423 34697 30435 34700
rect 30377 34691 30435 34697
rect 30742 34688 30748 34700
rect 30800 34688 30806 34740
rect 31478 34728 31484 34740
rect 31439 34700 31484 34728
rect 31478 34688 31484 34700
rect 31536 34688 31542 34740
rect 31570 34688 31576 34740
rect 31628 34688 31634 34740
rect 32214 34728 32220 34740
rect 32175 34700 32220 34728
rect 32214 34688 32220 34700
rect 32272 34688 32278 34740
rect 33410 34728 33416 34740
rect 33371 34700 33416 34728
rect 33410 34688 33416 34700
rect 33468 34688 33474 34740
rect 34146 34728 34152 34740
rect 34107 34700 34152 34728
rect 34146 34688 34152 34700
rect 34204 34688 34210 34740
rect 36262 34688 36268 34740
rect 36320 34728 36326 34740
rect 36455 34731 36513 34737
rect 36455 34728 36467 34731
rect 36320 34700 36467 34728
rect 36320 34688 36326 34700
rect 36455 34697 36467 34700
rect 36501 34697 36513 34731
rect 36455 34691 36513 34697
rect 38197 34731 38255 34737
rect 38197 34697 38209 34731
rect 38243 34728 38255 34731
rect 38286 34728 38292 34740
rect 38243 34700 38292 34728
rect 38243 34697 38255 34700
rect 38197 34691 38255 34697
rect 38286 34688 38292 34700
rect 38344 34688 38350 34740
rect 38565 34731 38623 34737
rect 38565 34697 38577 34731
rect 38611 34728 38623 34731
rect 38654 34728 38660 34740
rect 38611 34700 38660 34728
rect 38611 34697 38623 34700
rect 38565 34691 38623 34697
rect 38654 34688 38660 34700
rect 38712 34688 38718 34740
rect 39022 34688 39028 34740
rect 39080 34728 39086 34740
rect 39209 34731 39267 34737
rect 39209 34728 39221 34731
rect 39080 34700 39221 34728
rect 39080 34688 39086 34700
rect 39209 34697 39221 34700
rect 39255 34697 39267 34731
rect 39209 34691 39267 34697
rect 39853 34731 39911 34737
rect 39853 34697 39865 34731
rect 39899 34728 39911 34731
rect 39942 34728 39948 34740
rect 39899 34700 39948 34728
rect 39899 34697 39911 34700
rect 39853 34691 39911 34697
rect 39942 34688 39948 34700
rect 40000 34688 40006 34740
rect 41230 34688 41236 34740
rect 41288 34728 41294 34740
rect 41417 34731 41475 34737
rect 41417 34728 41429 34731
rect 41288 34700 41429 34728
rect 41288 34688 41294 34700
rect 41417 34697 41429 34700
rect 41463 34697 41475 34731
rect 41417 34691 41475 34697
rect 27614 34620 27620 34672
rect 27672 34620 27678 34672
rect 28258 34620 28264 34672
rect 28316 34660 28322 34672
rect 31294 34660 31300 34672
rect 28316 34632 29776 34660
rect 28316 34620 28322 34632
rect 27341 34595 27399 34601
rect 27341 34561 27353 34595
rect 27387 34561 27399 34595
rect 27632 34592 27660 34620
rect 27341 34555 27399 34561
rect 27448 34564 27660 34592
rect 25406 34524 25412 34536
rect 25056 34496 25412 34524
rect 25406 34484 25412 34496
rect 25464 34484 25470 34536
rect 25682 34484 25688 34536
rect 25740 34524 25746 34536
rect 25869 34527 25927 34533
rect 25869 34524 25881 34527
rect 25740 34496 25881 34524
rect 25740 34484 25746 34496
rect 25869 34493 25881 34496
rect 25915 34493 25927 34527
rect 27062 34524 27068 34536
rect 27023 34496 27068 34524
rect 25869 34487 25927 34493
rect 27062 34484 27068 34496
rect 27120 34484 27126 34536
rect 27246 34484 27252 34536
rect 27304 34524 27310 34536
rect 27448 34524 27476 34564
rect 28166 34552 28172 34604
rect 28224 34592 28230 34604
rect 28629 34595 28687 34601
rect 28629 34592 28641 34595
rect 28224 34564 28641 34592
rect 28224 34552 28230 34564
rect 28629 34561 28641 34564
rect 28675 34592 28687 34595
rect 28718 34592 28724 34604
rect 28675 34564 28724 34592
rect 28675 34561 28687 34564
rect 28629 34555 28687 34561
rect 28718 34552 28724 34564
rect 28776 34552 28782 34604
rect 28902 34592 28908 34604
rect 28863 34564 28908 34592
rect 28902 34552 28908 34564
rect 28960 34552 28966 34604
rect 29748 34601 29776 34632
rect 29840 34632 31300 34660
rect 29089 34595 29147 34601
rect 29089 34561 29101 34595
rect 29135 34592 29147 34595
rect 29549 34595 29607 34601
rect 29549 34592 29561 34595
rect 29135 34564 29561 34592
rect 29135 34561 29147 34564
rect 29089 34555 29147 34561
rect 29549 34561 29561 34564
rect 29595 34561 29607 34595
rect 29549 34555 29607 34561
rect 29733 34595 29791 34601
rect 29733 34561 29745 34595
rect 29779 34561 29791 34595
rect 29733 34555 29791 34561
rect 27304 34496 27476 34524
rect 27525 34527 27583 34533
rect 27304 34484 27310 34496
rect 27525 34493 27537 34527
rect 27571 34524 27583 34527
rect 27614 34524 27620 34536
rect 27571 34496 27620 34524
rect 27571 34493 27583 34496
rect 27525 34487 27583 34493
rect 27614 34484 27620 34496
rect 27672 34484 27678 34536
rect 28810 34524 28816 34536
rect 28771 34496 28816 34524
rect 28810 34484 28816 34496
rect 28868 34484 28874 34536
rect 29564 34524 29592 34555
rect 29840 34524 29868 34632
rect 31294 34620 31300 34632
rect 31352 34620 31358 34672
rect 31588 34660 31616 34688
rect 32677 34663 32735 34669
rect 32677 34660 32689 34663
rect 31588 34632 32689 34660
rect 32677 34629 32689 34632
rect 32723 34629 32735 34663
rect 35894 34660 35900 34672
rect 32677 34623 32735 34629
rect 34440 34632 35900 34660
rect 29914 34552 29920 34604
rect 29972 34592 29978 34604
rect 30742 34592 30748 34604
rect 29972 34564 30017 34592
rect 30703 34564 30748 34592
rect 29972 34552 29978 34564
rect 30742 34552 30748 34564
rect 30800 34552 30806 34604
rect 31573 34595 31631 34601
rect 31573 34561 31585 34595
rect 31619 34592 31631 34595
rect 31754 34592 31760 34604
rect 31619 34564 31760 34592
rect 31619 34561 31631 34564
rect 31573 34555 31631 34561
rect 31754 34552 31760 34564
rect 31812 34552 31818 34604
rect 33318 34592 33324 34604
rect 33279 34564 33324 34592
rect 33318 34552 33324 34564
rect 33376 34552 33382 34604
rect 33594 34592 33600 34604
rect 33555 34564 33600 34592
rect 33594 34552 33600 34564
rect 33652 34552 33658 34604
rect 34440 34601 34468 34632
rect 35894 34620 35900 34632
rect 35952 34620 35958 34672
rect 36541 34663 36599 34669
rect 36541 34660 36553 34663
rect 36280 34632 36553 34660
rect 33689 34595 33747 34601
rect 33689 34561 33701 34595
rect 33735 34592 33747 34595
rect 34425 34595 34483 34601
rect 33735 34564 34376 34592
rect 33735 34561 33747 34564
rect 33689 34555 33747 34561
rect 30834 34524 30840 34536
rect 29564 34496 29868 34524
rect 30795 34496 30840 34524
rect 30834 34484 30840 34496
rect 30892 34484 30898 34536
rect 33505 34527 33563 34533
rect 33505 34493 33517 34527
rect 33551 34524 33563 34527
rect 33962 34524 33968 34536
rect 33551 34496 33968 34524
rect 33551 34493 33563 34496
rect 33505 34487 33563 34493
rect 22649 34459 22707 34465
rect 22649 34425 22661 34459
rect 22695 34425 22707 34459
rect 23492 34456 23520 34484
rect 28350 34456 28356 34468
rect 23492 34428 28356 34456
rect 22649 34419 22707 34425
rect 28350 34416 28356 34428
rect 28408 34416 28414 34468
rect 28718 34456 28724 34468
rect 28679 34428 28724 34456
rect 28718 34416 28724 34428
rect 28776 34416 28782 34468
rect 30098 34416 30104 34468
rect 30156 34456 30162 34468
rect 33520 34456 33548 34487
rect 33962 34484 33968 34496
rect 34020 34484 34026 34536
rect 34149 34527 34207 34533
rect 34149 34493 34161 34527
rect 34195 34524 34207 34527
rect 34238 34524 34244 34536
rect 34195 34496 34244 34524
rect 34195 34493 34207 34496
rect 34149 34487 34207 34493
rect 34238 34484 34244 34496
rect 34296 34484 34302 34536
rect 34348 34524 34376 34564
rect 34425 34561 34437 34595
rect 34471 34561 34483 34595
rect 35526 34592 35532 34604
rect 35487 34564 35532 34592
rect 34425 34555 34483 34561
rect 35526 34552 35532 34564
rect 35584 34592 35590 34604
rect 36280 34592 36308 34632
rect 36541 34629 36553 34632
rect 36587 34660 36599 34663
rect 36722 34660 36728 34672
rect 36587 34632 36728 34660
rect 36587 34629 36599 34632
rect 36541 34623 36599 34629
rect 36722 34620 36728 34632
rect 36780 34660 36786 34672
rect 37369 34663 37427 34669
rect 37369 34660 37381 34663
rect 36780 34632 37381 34660
rect 36780 34620 36786 34632
rect 37369 34629 37381 34632
rect 37415 34660 37427 34663
rect 37415 34632 42104 34660
rect 37415 34629 37427 34632
rect 37369 34623 37427 34629
rect 35584 34564 36308 34592
rect 36357 34595 36415 34601
rect 35584 34552 35590 34564
rect 36357 34561 36369 34595
rect 36403 34592 36415 34595
rect 36446 34592 36452 34604
rect 36403 34564 36452 34592
rect 36403 34561 36415 34564
rect 36357 34555 36415 34561
rect 36446 34552 36452 34564
rect 36504 34552 36510 34604
rect 36633 34595 36691 34601
rect 36633 34561 36645 34595
rect 36679 34592 36691 34595
rect 37277 34595 37335 34601
rect 37277 34592 37289 34595
rect 36679 34564 37289 34592
rect 36679 34561 36691 34564
rect 36633 34555 36691 34561
rect 37277 34561 37289 34564
rect 37323 34561 37335 34595
rect 37550 34592 37556 34604
rect 37511 34564 37556 34592
rect 37277 34555 37335 34561
rect 35434 34524 35440 34536
rect 34348 34496 35440 34524
rect 35434 34484 35440 34496
rect 35492 34484 35498 34536
rect 35621 34527 35679 34533
rect 35621 34493 35633 34527
rect 35667 34524 35679 34527
rect 36262 34524 36268 34536
rect 35667 34496 36268 34524
rect 35667 34493 35679 34496
rect 35621 34487 35679 34493
rect 36262 34484 36268 34496
rect 36320 34524 36326 34536
rect 36648 34524 36676 34555
rect 37550 34552 37556 34564
rect 37608 34552 37614 34604
rect 38102 34552 38108 34604
rect 38160 34592 38166 34604
rect 38381 34595 38439 34601
rect 38381 34592 38393 34595
rect 38160 34564 38393 34592
rect 38160 34552 38166 34564
rect 38381 34561 38393 34564
rect 38427 34561 38439 34595
rect 38381 34555 38439 34561
rect 38657 34595 38715 34601
rect 38657 34561 38669 34595
rect 38703 34592 38715 34595
rect 39114 34592 39120 34604
rect 38703 34564 38737 34592
rect 39075 34564 39120 34592
rect 38703 34561 38715 34564
rect 38657 34555 38715 34561
rect 36320 34496 36676 34524
rect 37737 34527 37795 34533
rect 36320 34484 36326 34496
rect 37737 34493 37749 34527
rect 37783 34524 37795 34527
rect 38672 34524 38700 34555
rect 39114 34552 39120 34564
rect 39172 34552 39178 34604
rect 39298 34592 39304 34604
rect 39224 34564 39304 34592
rect 39224 34524 39252 34564
rect 39298 34552 39304 34564
rect 39356 34552 39362 34604
rect 40402 34592 40408 34604
rect 40363 34564 40408 34592
rect 40402 34552 40408 34564
rect 40460 34552 40466 34604
rect 40586 34592 40592 34604
rect 40547 34564 40592 34592
rect 40586 34552 40592 34564
rect 40644 34552 40650 34604
rect 42076 34536 42104 34632
rect 37783 34496 39252 34524
rect 37783 34493 37795 34496
rect 37737 34487 37795 34493
rect 42058 34484 42064 34536
rect 42116 34524 42122 34536
rect 42521 34527 42579 34533
rect 42521 34524 42533 34527
rect 42116 34496 42533 34524
rect 42116 34484 42122 34496
rect 42521 34493 42533 34496
rect 42567 34524 42579 34527
rect 42981 34527 43039 34533
rect 42981 34524 42993 34527
rect 42567 34496 42993 34524
rect 42567 34493 42579 34496
rect 42521 34487 42579 34493
rect 42981 34493 42993 34496
rect 43027 34493 43039 34527
rect 42981 34487 43039 34493
rect 30156 34428 33548 34456
rect 30156 34416 30162 34428
rect 33686 34416 33692 34468
rect 33744 34456 33750 34468
rect 33744 34428 34468 34456
rect 33744 34416 33750 34428
rect 9766 34388 9772 34400
rect 9727 34360 9772 34388
rect 9766 34348 9772 34360
rect 9824 34348 9830 34400
rect 11514 34348 11520 34400
rect 11572 34388 11578 34400
rect 11885 34391 11943 34397
rect 11885 34388 11897 34391
rect 11572 34360 11897 34388
rect 11572 34348 11578 34360
rect 11885 34357 11897 34360
rect 11931 34357 11943 34391
rect 11885 34351 11943 34357
rect 14093 34391 14151 34397
rect 14093 34357 14105 34391
rect 14139 34388 14151 34391
rect 14826 34388 14832 34400
rect 14139 34360 14832 34388
rect 14139 34357 14151 34360
rect 14093 34351 14151 34357
rect 14826 34348 14832 34360
rect 14884 34348 14890 34400
rect 17954 34348 17960 34400
rect 18012 34388 18018 34400
rect 18049 34391 18107 34397
rect 18049 34388 18061 34391
rect 18012 34360 18061 34388
rect 18012 34348 18018 34360
rect 18049 34357 18061 34360
rect 18095 34357 18107 34391
rect 18049 34351 18107 34357
rect 20349 34391 20407 34397
rect 20349 34357 20361 34391
rect 20395 34388 20407 34391
rect 22002 34388 22008 34400
rect 20395 34360 22008 34388
rect 20395 34357 20407 34360
rect 20349 34351 20407 34357
rect 22002 34348 22008 34360
rect 22060 34348 22066 34400
rect 25038 34388 25044 34400
rect 24999 34360 25044 34388
rect 25038 34348 25044 34360
rect 25096 34348 25102 34400
rect 28442 34388 28448 34400
rect 28403 34360 28448 34388
rect 28442 34348 28448 34360
rect 28500 34348 28506 34400
rect 33962 34348 33968 34400
rect 34020 34388 34026 34400
rect 34333 34391 34391 34397
rect 34333 34388 34345 34391
rect 34020 34360 34345 34388
rect 34020 34348 34026 34360
rect 34333 34357 34345 34360
rect 34379 34357 34391 34391
rect 34440 34388 34468 34428
rect 35710 34416 35716 34468
rect 35768 34456 35774 34468
rect 35897 34459 35955 34465
rect 35897 34456 35909 34459
rect 35768 34428 35909 34456
rect 35768 34416 35774 34428
rect 35897 34425 35909 34428
rect 35943 34425 35955 34459
rect 35897 34419 35955 34425
rect 39850 34388 39856 34400
rect 34440 34360 39856 34388
rect 34333 34351 34391 34357
rect 39850 34348 39856 34360
rect 39908 34348 39914 34400
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 10226 34144 10232 34196
rect 10284 34184 10290 34196
rect 10321 34187 10379 34193
rect 10321 34184 10333 34187
rect 10284 34156 10333 34184
rect 10284 34144 10290 34156
rect 10321 34153 10333 34156
rect 10367 34153 10379 34187
rect 10321 34147 10379 34153
rect 14645 34187 14703 34193
rect 14645 34153 14657 34187
rect 14691 34184 14703 34187
rect 14734 34184 14740 34196
rect 14691 34156 14740 34184
rect 14691 34153 14703 34156
rect 14645 34147 14703 34153
rect 14734 34144 14740 34156
rect 14792 34144 14798 34196
rect 15381 34187 15439 34193
rect 15381 34153 15393 34187
rect 15427 34184 15439 34187
rect 15562 34184 15568 34196
rect 15427 34156 15568 34184
rect 15427 34153 15439 34156
rect 15381 34147 15439 34153
rect 15562 34144 15568 34156
rect 15620 34144 15626 34196
rect 16117 34187 16175 34193
rect 16117 34153 16129 34187
rect 16163 34184 16175 34187
rect 16850 34184 16856 34196
rect 16163 34156 16856 34184
rect 16163 34153 16175 34156
rect 16117 34147 16175 34153
rect 1578 34116 1584 34128
rect 1539 34088 1584 34116
rect 1578 34076 1584 34088
rect 1636 34076 1642 34128
rect 13541 34119 13599 34125
rect 13541 34085 13553 34119
rect 13587 34085 13599 34119
rect 16132 34116 16160 34147
rect 16850 34144 16856 34156
rect 16908 34144 16914 34196
rect 17954 34184 17960 34196
rect 17915 34156 17960 34184
rect 17954 34144 17960 34156
rect 18012 34144 18018 34196
rect 21634 34184 21640 34196
rect 21595 34156 21640 34184
rect 21634 34144 21640 34156
rect 21692 34144 21698 34196
rect 21821 34187 21879 34193
rect 21821 34153 21833 34187
rect 21867 34184 21879 34187
rect 22554 34184 22560 34196
rect 21867 34156 22560 34184
rect 21867 34153 21879 34156
rect 21821 34147 21879 34153
rect 22554 34144 22560 34156
rect 22612 34144 22618 34196
rect 25130 34184 25136 34196
rect 25091 34156 25136 34184
rect 25130 34144 25136 34156
rect 25188 34144 25194 34196
rect 25222 34144 25228 34196
rect 25280 34184 25286 34196
rect 25317 34187 25375 34193
rect 25317 34184 25329 34187
rect 25280 34156 25329 34184
rect 25280 34144 25286 34156
rect 25317 34153 25329 34156
rect 25363 34153 25375 34187
rect 25317 34147 25375 34153
rect 25498 34144 25504 34196
rect 25556 34184 25562 34196
rect 25866 34184 25872 34196
rect 25556 34156 25872 34184
rect 25556 34144 25562 34156
rect 25866 34144 25872 34156
rect 25924 34144 25930 34196
rect 27614 34184 27620 34196
rect 27575 34156 27620 34184
rect 27614 34144 27620 34156
rect 27672 34144 27678 34196
rect 28721 34187 28779 34193
rect 28721 34153 28733 34187
rect 28767 34184 28779 34187
rect 29270 34184 29276 34196
rect 28767 34156 29276 34184
rect 28767 34153 28779 34156
rect 28721 34147 28779 34153
rect 29270 34144 29276 34156
rect 29328 34144 29334 34196
rect 29546 34144 29552 34196
rect 29604 34184 29610 34196
rect 29825 34187 29883 34193
rect 29825 34184 29837 34187
rect 29604 34156 29837 34184
rect 29604 34144 29610 34156
rect 29825 34153 29837 34156
rect 29871 34153 29883 34187
rect 29825 34147 29883 34153
rect 31386 34144 31392 34196
rect 31444 34184 31450 34196
rect 31849 34187 31907 34193
rect 31849 34184 31861 34187
rect 31444 34156 31861 34184
rect 31444 34144 31450 34156
rect 31849 34153 31861 34156
rect 31895 34184 31907 34187
rect 32398 34184 32404 34196
rect 31895 34156 32404 34184
rect 31895 34153 31907 34156
rect 31849 34147 31907 34153
rect 32398 34144 32404 34156
rect 32456 34144 32462 34196
rect 33689 34187 33747 34193
rect 33689 34153 33701 34187
rect 33735 34153 33747 34187
rect 33689 34147 33747 34153
rect 13541 34079 13599 34085
rect 15396 34088 16160 34116
rect 11514 34048 11520 34060
rect 11475 34020 11520 34048
rect 11514 34008 11520 34020
rect 11572 34008 11578 34060
rect 11974 34048 11980 34060
rect 11935 34020 11980 34048
rect 11974 34008 11980 34020
rect 12032 34008 12038 34060
rect 13262 34048 13268 34060
rect 13223 34020 13268 34048
rect 13262 34008 13268 34020
rect 13320 34008 13326 34060
rect 13556 34048 13584 34079
rect 13814 34048 13820 34060
rect 13556 34020 13820 34048
rect 13814 34008 13820 34020
rect 13872 34048 13878 34060
rect 13872 34020 14504 34048
rect 13872 34008 13878 34020
rect 10870 33980 10876 33992
rect 10831 33952 10876 33980
rect 10870 33940 10876 33952
rect 10928 33940 10934 33992
rect 11057 33983 11115 33989
rect 11057 33949 11069 33983
rect 11103 33980 11115 33983
rect 11606 33980 11612 33992
rect 11103 33952 11612 33980
rect 11103 33949 11115 33952
rect 11057 33943 11115 33949
rect 11606 33940 11612 33952
rect 11664 33980 11670 33992
rect 11885 33983 11943 33989
rect 11885 33980 11897 33983
rect 11664 33952 11897 33980
rect 11664 33940 11670 33952
rect 11885 33949 11897 33952
rect 11931 33980 11943 33983
rect 12066 33980 12072 33992
rect 11931 33952 12072 33980
rect 11931 33949 11943 33952
rect 11885 33943 11943 33949
rect 12066 33940 12072 33952
rect 12124 33940 12130 33992
rect 12894 33980 12900 33992
rect 12406 33952 12900 33980
rect 10965 33915 11023 33921
rect 10965 33881 10977 33915
rect 11011 33912 11023 33915
rect 12406 33912 12434 33952
rect 12894 33940 12900 33952
rect 12952 33980 12958 33992
rect 13173 33983 13231 33989
rect 13173 33980 13185 33983
rect 12952 33952 13185 33980
rect 12952 33940 12958 33952
rect 13173 33949 13185 33952
rect 13219 33949 13231 33983
rect 14274 33980 14280 33992
rect 14235 33952 14280 33980
rect 13173 33943 13231 33949
rect 14274 33940 14280 33952
rect 14332 33940 14338 33992
rect 14476 33989 14504 34020
rect 14461 33983 14519 33989
rect 14461 33949 14473 33983
rect 14507 33949 14519 33983
rect 14461 33943 14519 33949
rect 14826 33940 14832 33992
rect 14884 33980 14890 33992
rect 15010 33980 15016 33992
rect 14884 33952 15016 33980
rect 14884 33940 14890 33952
rect 15010 33940 15016 33952
rect 15068 33980 15074 33992
rect 15105 33983 15163 33989
rect 15105 33980 15117 33983
rect 15068 33952 15117 33980
rect 15068 33940 15074 33952
rect 15105 33949 15117 33952
rect 15151 33949 15163 33983
rect 15105 33943 15163 33949
rect 15197 33983 15255 33989
rect 15197 33949 15209 33983
rect 15243 33980 15255 33983
rect 15396 33980 15424 34088
rect 16666 34076 16672 34128
rect 16724 34116 16730 34128
rect 16945 34119 17003 34125
rect 16945 34116 16957 34119
rect 16724 34088 16957 34116
rect 16724 34076 16730 34088
rect 16945 34085 16957 34088
rect 16991 34085 17003 34119
rect 16945 34079 17003 34085
rect 19058 34076 19064 34128
rect 19116 34116 19122 34128
rect 23201 34119 23259 34125
rect 19116 34088 23152 34116
rect 19116 34076 19122 34088
rect 16040 34020 17816 34048
rect 15243 33952 15424 33980
rect 15243 33949 15255 33952
rect 15197 33943 15255 33949
rect 15470 33940 15476 33992
rect 15528 33980 15534 33992
rect 16040 33989 16068 34020
rect 16025 33983 16083 33989
rect 16025 33980 16037 33983
rect 15528 33952 16037 33980
rect 15528 33940 15534 33952
rect 16025 33949 16037 33952
rect 16071 33949 16083 33983
rect 16025 33943 16083 33949
rect 16209 33983 16267 33989
rect 16209 33949 16221 33983
rect 16255 33949 16267 33983
rect 16209 33943 16267 33949
rect 15381 33915 15439 33921
rect 15381 33912 15393 33915
rect 11011 33884 12434 33912
rect 14476 33884 15393 33912
rect 11011 33881 11023 33884
rect 10965 33875 11023 33881
rect 14476 33856 14504 33884
rect 15381 33881 15393 33884
rect 15427 33881 15439 33915
rect 16224 33912 16252 33943
rect 16574 33940 16580 33992
rect 16632 33980 16638 33992
rect 17788 33989 17816 34020
rect 19242 34008 19248 34060
rect 19300 34048 19306 34060
rect 19521 34051 19579 34057
rect 19521 34048 19533 34051
rect 19300 34020 19533 34048
rect 19300 34008 19306 34020
rect 19521 34017 19533 34020
rect 19567 34017 19579 34051
rect 19521 34011 19579 34017
rect 20438 34008 20444 34060
rect 20496 34048 20502 34060
rect 20625 34051 20683 34057
rect 20625 34048 20637 34051
rect 20496 34020 20637 34048
rect 20496 34008 20502 34020
rect 20625 34017 20637 34020
rect 20671 34017 20683 34051
rect 22922 34048 22928 34060
rect 22883 34020 22928 34048
rect 20625 34011 20683 34017
rect 22922 34008 22928 34020
rect 22980 34008 22986 34060
rect 23124 34048 23152 34088
rect 23201 34085 23213 34119
rect 23247 34116 23259 34119
rect 24210 34116 24216 34128
rect 23247 34088 24216 34116
rect 23247 34085 23259 34088
rect 23201 34079 23259 34085
rect 24210 34076 24216 34088
rect 24268 34076 24274 34128
rect 27433 34119 27491 34125
rect 27433 34085 27445 34119
rect 27479 34116 27491 34119
rect 27982 34116 27988 34128
rect 27479 34088 27988 34116
rect 27479 34085 27491 34088
rect 27433 34079 27491 34085
rect 27982 34076 27988 34088
rect 28040 34076 28046 34128
rect 30834 34116 30840 34128
rect 30024 34088 30840 34116
rect 23753 34051 23811 34057
rect 23753 34048 23765 34051
rect 23124 34020 23765 34048
rect 23753 34017 23765 34020
rect 23799 34048 23811 34051
rect 25041 34051 25099 34057
rect 25041 34048 25053 34051
rect 23799 34020 25053 34048
rect 23799 34017 23811 34020
rect 23753 34011 23811 34017
rect 25041 34017 25053 34020
rect 25087 34048 25099 34051
rect 27522 34048 27528 34060
rect 25087 34020 27528 34048
rect 25087 34017 25099 34020
rect 25041 34011 25099 34017
rect 27522 34008 27528 34020
rect 27580 34008 27586 34060
rect 16669 33983 16727 33989
rect 16669 33980 16681 33983
rect 16632 33952 16681 33980
rect 16632 33940 16638 33952
rect 16669 33949 16681 33952
rect 16715 33949 16727 33983
rect 16669 33943 16727 33949
rect 17773 33983 17831 33989
rect 17773 33949 17785 33983
rect 17819 33949 17831 33983
rect 17773 33943 17831 33949
rect 18414 33940 18420 33992
rect 18472 33980 18478 33992
rect 18601 33983 18659 33989
rect 18601 33980 18613 33983
rect 18472 33952 18613 33980
rect 18472 33940 18478 33952
rect 18601 33949 18613 33952
rect 18647 33949 18659 33983
rect 18601 33943 18659 33949
rect 19334 33940 19340 33992
rect 19392 33980 19398 33992
rect 19613 33983 19671 33989
rect 19613 33980 19625 33983
rect 19392 33952 19625 33980
rect 19392 33940 19398 33952
rect 19613 33949 19625 33952
rect 19659 33949 19671 33983
rect 19613 33943 19671 33949
rect 20533 33983 20591 33989
rect 20533 33949 20545 33983
rect 20579 33980 20591 33983
rect 21450 33980 21456 33992
rect 20579 33952 21456 33980
rect 20579 33949 20591 33952
rect 20533 33943 20591 33949
rect 21450 33940 21456 33952
rect 21508 33940 21514 33992
rect 21542 33940 21548 33992
rect 21600 33980 21606 33992
rect 22830 33980 22836 33992
rect 21600 33952 21693 33980
rect 22791 33952 22836 33980
rect 21600 33940 21606 33952
rect 22830 33940 22836 33952
rect 22888 33940 22894 33992
rect 24762 33980 24768 33992
rect 24723 33952 24768 33980
rect 24762 33940 24768 33952
rect 24820 33940 24826 33992
rect 26786 33980 26792 33992
rect 26747 33952 26792 33980
rect 26786 33940 26792 33952
rect 26844 33940 26850 33992
rect 26970 33980 26976 33992
rect 26931 33952 26976 33980
rect 26970 33940 26976 33952
rect 27028 33940 27034 33992
rect 27985 33983 28043 33989
rect 27985 33949 27997 33983
rect 28031 33980 28043 33983
rect 28258 33980 28264 33992
rect 28031 33952 28264 33980
rect 28031 33949 28043 33952
rect 27985 33943 28043 33949
rect 28258 33940 28264 33952
rect 28316 33940 28322 33992
rect 28442 33980 28448 33992
rect 28403 33952 28448 33980
rect 28442 33940 28448 33952
rect 28500 33940 28506 33992
rect 30024 33989 30052 34088
rect 30834 34076 30840 34088
rect 30892 34076 30898 34128
rect 32306 34048 32312 34060
rect 30208 34020 32312 34048
rect 30208 33989 30236 34020
rect 32306 34008 32312 34020
rect 32364 34048 32370 34060
rect 32364 34020 32996 34048
rect 32364 34008 32370 34020
rect 30009 33983 30067 33989
rect 30009 33949 30021 33983
rect 30055 33949 30067 33983
rect 30009 33943 30067 33949
rect 30193 33983 30251 33989
rect 30193 33949 30205 33983
rect 30239 33949 30251 33983
rect 30193 33943 30251 33949
rect 30469 33983 30527 33989
rect 30469 33949 30481 33983
rect 30515 33980 30527 33983
rect 30926 33980 30932 33992
rect 30515 33952 30932 33980
rect 30515 33949 30527 33952
rect 30469 33943 30527 33949
rect 30926 33940 30932 33952
rect 30984 33940 30990 33992
rect 31294 33980 31300 33992
rect 31255 33952 31300 33980
rect 31294 33940 31300 33952
rect 31352 33940 31358 33992
rect 17589 33915 17647 33921
rect 17589 33912 17601 33915
rect 16224 33884 17601 33912
rect 15381 33875 15439 33881
rect 17589 33881 17601 33884
rect 17635 33912 17647 33915
rect 18690 33912 18696 33924
rect 17635 33884 18696 33912
rect 17635 33881 17647 33884
rect 17589 33875 17647 33881
rect 18690 33872 18696 33884
rect 18748 33872 18754 33924
rect 20809 33915 20867 33921
rect 20809 33881 20821 33915
rect 20855 33912 20867 33915
rect 20990 33912 20996 33924
rect 20855 33884 20996 33912
rect 20855 33881 20867 33884
rect 20809 33875 20867 33881
rect 20990 33872 20996 33884
rect 21048 33912 21054 33924
rect 21560 33912 21588 33940
rect 21048 33884 21588 33912
rect 21048 33872 21054 33884
rect 25406 33872 25412 33924
rect 25464 33912 25470 33924
rect 27706 33912 27712 33924
rect 25464 33884 27712 33912
rect 25464 33872 25470 33884
rect 27706 33872 27712 33884
rect 27764 33912 27770 33924
rect 28721 33915 28779 33921
rect 28721 33912 28733 33915
rect 27764 33884 28733 33912
rect 27764 33872 27770 33884
rect 28721 33881 28733 33884
rect 28767 33881 28779 33915
rect 28721 33875 28779 33881
rect 30101 33915 30159 33921
rect 30101 33881 30113 33915
rect 30147 33881 30159 33915
rect 30101 33875 30159 33881
rect 9766 33844 9772 33856
rect 9727 33816 9772 33844
rect 9766 33804 9772 33816
rect 9824 33804 9830 33856
rect 12161 33847 12219 33853
rect 12161 33813 12173 33847
rect 12207 33844 12219 33847
rect 12618 33844 12624 33856
rect 12207 33816 12624 33844
rect 12207 33813 12219 33816
rect 12161 33807 12219 33813
rect 12618 33804 12624 33816
rect 12676 33804 12682 33856
rect 14458 33804 14464 33856
rect 14516 33804 14522 33856
rect 17129 33847 17187 33853
rect 17129 33813 17141 33847
rect 17175 33844 17187 33847
rect 18506 33844 18512 33856
rect 17175 33816 18512 33844
rect 17175 33813 17187 33816
rect 17129 33807 17187 33813
rect 18506 33804 18512 33816
rect 18564 33804 18570 33856
rect 18966 33804 18972 33856
rect 19024 33844 19030 33856
rect 19245 33847 19303 33853
rect 19245 33844 19257 33847
rect 19024 33816 19257 33844
rect 19024 33804 19030 33816
rect 19245 33813 19257 33816
rect 19291 33813 19303 33847
rect 20530 33844 20536 33856
rect 20491 33816 20536 33844
rect 19245 33807 19303 33813
rect 20530 33804 20536 33816
rect 20588 33804 20594 33856
rect 26970 33844 26976 33856
rect 26931 33816 26976 33844
rect 26970 33804 26976 33816
rect 27028 33804 27034 33856
rect 27614 33844 27620 33856
rect 27575 33816 27620 33844
rect 27614 33804 27620 33816
rect 27672 33804 27678 33856
rect 28534 33844 28540 33856
rect 28495 33816 28540 33844
rect 28534 33804 28540 33816
rect 28592 33804 28598 33856
rect 30116 33844 30144 33875
rect 30282 33872 30288 33924
rect 30340 33921 30346 33924
rect 30340 33915 30369 33921
rect 30357 33881 30369 33915
rect 30340 33875 30369 33881
rect 31113 33915 31171 33921
rect 31113 33881 31125 33915
rect 31159 33912 31171 33915
rect 31386 33912 31392 33924
rect 31159 33884 31392 33912
rect 31159 33881 31171 33884
rect 31113 33875 31171 33881
rect 30340 33872 30346 33875
rect 31386 33872 31392 33884
rect 31444 33872 31450 33924
rect 30929 33847 30987 33853
rect 30929 33844 30941 33847
rect 30116 33816 30941 33844
rect 30929 33813 30941 33816
rect 30975 33813 30987 33847
rect 30929 33807 30987 33813
rect 31570 33804 31576 33856
rect 31628 33844 31634 33856
rect 32861 33847 32919 33853
rect 32861 33844 32873 33847
rect 31628 33816 32873 33844
rect 31628 33804 31634 33816
rect 32861 33813 32873 33816
rect 32907 33813 32919 33847
rect 32968 33844 32996 34020
rect 33134 34008 33140 34060
rect 33192 34048 33198 34060
rect 33704 34048 33732 34147
rect 33778 34144 33784 34196
rect 33836 34184 33842 34196
rect 34422 34184 34428 34196
rect 33836 34156 34428 34184
rect 33836 34144 33842 34156
rect 34422 34144 34428 34156
rect 34480 34184 34486 34196
rect 34701 34187 34759 34193
rect 34701 34184 34713 34187
rect 34480 34156 34713 34184
rect 34480 34144 34486 34156
rect 34701 34153 34713 34156
rect 34747 34153 34759 34187
rect 34701 34147 34759 34153
rect 34716 34116 34744 34147
rect 35434 34144 35440 34196
rect 35492 34184 35498 34196
rect 35621 34187 35679 34193
rect 35621 34184 35633 34187
rect 35492 34156 35633 34184
rect 35492 34144 35498 34156
rect 35621 34153 35633 34156
rect 35667 34153 35679 34187
rect 35621 34147 35679 34153
rect 36262 34144 36268 34196
rect 36320 34184 36326 34196
rect 36449 34187 36507 34193
rect 36449 34184 36461 34187
rect 36320 34156 36461 34184
rect 36320 34144 36326 34156
rect 36449 34153 36461 34156
rect 36495 34184 36507 34187
rect 36495 34156 37228 34184
rect 36495 34153 36507 34156
rect 36449 34147 36507 34153
rect 37200 34125 37228 34156
rect 39666 34144 39672 34196
rect 39724 34184 39730 34196
rect 39853 34187 39911 34193
rect 39853 34184 39865 34187
rect 39724 34156 39865 34184
rect 39724 34144 39730 34156
rect 39853 34153 39865 34156
rect 39899 34153 39911 34187
rect 42058 34184 42064 34196
rect 42019 34156 42064 34184
rect 39853 34147 39911 34153
rect 42058 34144 42064 34156
rect 42116 34144 42122 34196
rect 35713 34119 35771 34125
rect 35713 34116 35725 34119
rect 34716 34088 35725 34116
rect 35713 34085 35725 34088
rect 35759 34085 35771 34119
rect 35713 34079 35771 34085
rect 37185 34119 37243 34125
rect 37185 34085 37197 34119
rect 37231 34085 37243 34119
rect 37185 34079 37243 34085
rect 37550 34076 37556 34128
rect 37608 34116 37614 34128
rect 38841 34119 38899 34125
rect 37608 34088 38516 34116
rect 37608 34076 37614 34088
rect 35342 34048 35348 34060
rect 33192 34020 35348 34048
rect 33192 34008 33198 34020
rect 35342 34008 35348 34020
rect 35400 34008 35406 34060
rect 35526 34048 35532 34060
rect 35487 34020 35532 34048
rect 35526 34008 35532 34020
rect 35584 34008 35590 34060
rect 38194 34048 38200 34060
rect 38155 34020 38200 34048
rect 38194 34008 38200 34020
rect 38252 34008 38258 34060
rect 38488 34057 38516 34088
rect 38841 34085 38853 34119
rect 38887 34116 38899 34119
rect 40310 34116 40316 34128
rect 38887 34088 40316 34116
rect 38887 34085 38899 34088
rect 38841 34079 38899 34085
rect 40310 34076 40316 34088
rect 40368 34076 40374 34128
rect 40770 34076 40776 34128
rect 40828 34116 40834 34128
rect 42518 34116 42524 34128
rect 40828 34088 42524 34116
rect 40828 34076 40834 34088
rect 42518 34076 42524 34088
rect 42576 34076 42582 34128
rect 38473 34051 38531 34057
rect 38473 34017 38485 34051
rect 38519 34017 38531 34051
rect 38473 34011 38531 34017
rect 38654 34008 38660 34060
rect 38712 34057 38718 34060
rect 38712 34051 38740 34057
rect 38728 34017 38740 34051
rect 38712 34011 38740 34017
rect 40497 34051 40555 34057
rect 40497 34017 40509 34051
rect 40543 34048 40555 34051
rect 40586 34048 40592 34060
rect 40543 34020 40592 34048
rect 40543 34017 40555 34020
rect 40497 34011 40555 34017
rect 38712 34008 38718 34011
rect 33318 33940 33324 33992
rect 33376 33980 33382 33992
rect 33505 33983 33563 33989
rect 33505 33980 33517 33983
rect 33376 33952 33517 33980
rect 33376 33940 33382 33952
rect 33505 33949 33517 33952
rect 33551 33980 33563 33983
rect 33686 33980 33692 33992
rect 33551 33952 33692 33980
rect 33551 33949 33563 33952
rect 33505 33943 33563 33949
rect 33686 33940 33692 33952
rect 33744 33940 33750 33992
rect 33962 33940 33968 33992
rect 34020 33980 34026 33992
rect 34885 33983 34943 33989
rect 34885 33980 34897 33983
rect 34020 33952 34897 33980
rect 34020 33940 34026 33952
rect 34885 33949 34897 33952
rect 34931 33949 34943 33983
rect 34885 33943 34943 33949
rect 35069 33983 35127 33989
rect 35069 33949 35081 33983
rect 35115 33949 35127 33983
rect 35802 33980 35808 33992
rect 35763 33952 35808 33980
rect 35069 33943 35127 33949
rect 33042 33872 33048 33924
rect 33100 33912 33106 33924
rect 35084 33912 35112 33943
rect 35802 33940 35808 33952
rect 35860 33940 35866 33992
rect 36170 33940 36176 33992
rect 36228 33980 36234 33992
rect 36265 33983 36323 33989
rect 36265 33980 36277 33983
rect 36228 33952 36277 33980
rect 36228 33940 36234 33952
rect 36265 33949 36277 33952
rect 36311 33949 36323 33983
rect 36446 33980 36452 33992
rect 36407 33952 36452 33980
rect 36265 33943 36323 33949
rect 36446 33940 36452 33952
rect 36504 33940 36510 33992
rect 37366 33980 37372 33992
rect 37327 33952 37372 33980
rect 37366 33940 37372 33952
rect 37424 33940 37430 33992
rect 37461 33983 37519 33989
rect 37461 33949 37473 33983
rect 37507 33980 37519 33983
rect 38102 33980 38108 33992
rect 37507 33952 38108 33980
rect 37507 33949 37519 33952
rect 37461 33943 37519 33949
rect 38102 33940 38108 33952
rect 38160 33940 38166 33992
rect 38565 33983 38623 33989
rect 38565 33949 38577 33983
rect 38611 33980 38623 33983
rect 40512 33980 40540 34011
rect 40586 34008 40592 34020
rect 40644 34008 40650 34060
rect 48130 34048 48136 34060
rect 48091 34020 48136 34048
rect 48130 34008 48136 34020
rect 48188 34008 48194 34060
rect 38611 33952 40540 33980
rect 40776 33992 40828 33998
rect 38611 33949 38623 33952
rect 38565 33943 38623 33949
rect 35894 33912 35900 33924
rect 33100 33884 35020 33912
rect 35084 33884 35900 33912
rect 33100 33872 33106 33884
rect 33778 33844 33784 33856
rect 32968 33816 33784 33844
rect 32861 33807 32919 33813
rect 33778 33804 33784 33816
rect 33836 33804 33842 33856
rect 33962 33844 33968 33856
rect 33923 33816 33968 33844
rect 33962 33804 33968 33816
rect 34020 33804 34026 33856
rect 34992 33844 35020 33884
rect 35894 33872 35900 33884
rect 35952 33872 35958 33924
rect 37553 33915 37611 33921
rect 37553 33881 37565 33915
rect 37599 33912 37611 33915
rect 38580 33912 38608 33943
rect 41417 33983 41475 33989
rect 41417 33949 41429 33983
rect 41463 33980 41475 33983
rect 47854 33980 47860 33992
rect 41463 33952 43208 33980
rect 47815 33952 47860 33980
rect 41463 33949 41475 33952
rect 41417 33943 41475 33949
rect 40776 33934 40828 33940
rect 41432 33912 41460 33943
rect 37599 33884 38608 33912
rect 41386 33884 41460 33912
rect 37599 33881 37611 33884
rect 37553 33875 37611 33881
rect 36078 33844 36084 33856
rect 34992 33816 36084 33844
rect 36078 33804 36084 33816
rect 36136 33804 36142 33856
rect 37737 33847 37795 33853
rect 37737 33813 37749 33847
rect 37783 33844 37795 33847
rect 37826 33844 37832 33856
rect 37783 33816 37832 33844
rect 37783 33813 37795 33816
rect 37737 33807 37795 33813
rect 37826 33804 37832 33816
rect 37884 33804 37890 33856
rect 40678 33804 40684 33856
rect 40736 33844 40742 33856
rect 41386 33844 41414 33884
rect 43180 33856 43208 33952
rect 47854 33940 47860 33952
rect 47912 33940 47918 33992
rect 43162 33844 43168 33856
rect 40736 33816 41414 33844
rect 43123 33816 43168 33844
rect 40736 33804 40742 33816
rect 43162 33804 43168 33816
rect 43220 33804 43226 33856
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 2038 33600 2044 33652
rect 2096 33640 2102 33652
rect 2096 33612 6914 33640
rect 2096 33600 2102 33612
rect 6886 33368 6914 33612
rect 10870 33600 10876 33652
rect 10928 33640 10934 33652
rect 11885 33643 11943 33649
rect 11885 33640 11897 33643
rect 10928 33612 11897 33640
rect 10928 33600 10934 33612
rect 11885 33609 11897 33612
rect 11931 33609 11943 33643
rect 11885 33603 11943 33609
rect 13262 33600 13268 33652
rect 13320 33640 13326 33652
rect 13718 33643 13776 33649
rect 13718 33640 13730 33643
rect 13320 33612 13730 33640
rect 13320 33600 13326 33612
rect 13718 33609 13730 33612
rect 13764 33609 13776 33643
rect 13718 33603 13776 33609
rect 15378 33600 15384 33652
rect 15436 33640 15442 33652
rect 15565 33643 15623 33649
rect 15565 33640 15577 33643
rect 15436 33612 15577 33640
rect 15436 33600 15442 33612
rect 15565 33609 15577 33612
rect 15611 33640 15623 33643
rect 16853 33643 16911 33649
rect 16853 33640 16865 33643
rect 15611 33612 16865 33640
rect 15611 33609 15623 33612
rect 15565 33603 15623 33609
rect 16853 33609 16865 33612
rect 16899 33609 16911 33643
rect 16853 33603 16911 33609
rect 17497 33643 17555 33649
rect 17497 33609 17509 33643
rect 17543 33640 17555 33643
rect 18138 33640 18144 33652
rect 17543 33612 18144 33640
rect 17543 33609 17555 33612
rect 17497 33603 17555 33609
rect 10413 33575 10471 33581
rect 10413 33541 10425 33575
rect 10459 33572 10471 33575
rect 11146 33572 11152 33584
rect 10459 33544 11152 33572
rect 10459 33541 10471 33544
rect 10413 33535 10471 33541
rect 11146 33532 11152 33544
rect 11204 33572 11210 33584
rect 11698 33572 11704 33584
rect 11204 33544 11704 33572
rect 11204 33532 11210 33544
rect 11698 33532 11704 33544
rect 11756 33532 11762 33584
rect 12710 33572 12716 33584
rect 12671 33544 12716 33572
rect 12710 33532 12716 33544
rect 12768 33532 12774 33584
rect 12894 33572 12900 33584
rect 12855 33544 12900 33572
rect 12894 33532 12900 33544
rect 12952 33532 12958 33584
rect 13446 33532 13452 33584
rect 13504 33572 13510 33584
rect 13633 33575 13691 33581
rect 13633 33572 13645 33575
rect 13504 33544 13645 33572
rect 13504 33532 13510 33544
rect 13633 33541 13645 33544
rect 13679 33541 13691 33575
rect 16669 33575 16727 33581
rect 16669 33572 16681 33575
rect 13633 33535 13691 33541
rect 15488 33544 16681 33572
rect 9861 33507 9919 33513
rect 9861 33473 9873 33507
rect 9907 33504 9919 33507
rect 10965 33507 11023 33513
rect 10965 33504 10977 33507
rect 9907 33476 10977 33504
rect 9907 33473 9919 33476
rect 9861 33467 9919 33473
rect 10965 33473 10977 33476
rect 11011 33504 11023 33507
rect 11514 33504 11520 33516
rect 11011 33476 11520 33504
rect 11011 33473 11023 33476
rect 10965 33467 11023 33473
rect 11514 33464 11520 33476
rect 11572 33464 11578 33516
rect 12802 33464 12808 33516
rect 12860 33504 12866 33516
rect 13541 33507 13599 33513
rect 13541 33504 13553 33507
rect 12860 33476 13553 33504
rect 12860 33464 12866 33476
rect 13541 33473 13553 33476
rect 13587 33473 13599 33507
rect 13814 33504 13820 33516
rect 13775 33476 13820 33504
rect 13541 33467 13599 33473
rect 13814 33464 13820 33476
rect 13872 33464 13878 33516
rect 14458 33464 14464 33516
rect 14516 33504 14522 33516
rect 14829 33507 14887 33513
rect 14829 33504 14841 33507
rect 14516 33476 14841 33504
rect 14516 33464 14522 33476
rect 14829 33473 14841 33476
rect 14875 33473 14887 33507
rect 15010 33504 15016 33516
rect 14971 33476 15016 33504
rect 14829 33467 14887 33473
rect 15010 33464 15016 33476
rect 15068 33464 15074 33516
rect 15286 33464 15292 33516
rect 15344 33504 15350 33516
rect 15488 33513 15516 33544
rect 16669 33541 16681 33544
rect 16715 33541 16727 33575
rect 17512 33572 17540 33603
rect 18138 33600 18144 33612
rect 18196 33600 18202 33652
rect 19242 33640 19248 33652
rect 19203 33612 19248 33640
rect 19242 33600 19248 33612
rect 19300 33600 19306 33652
rect 20993 33643 21051 33649
rect 20993 33640 21005 33643
rect 20180 33612 21005 33640
rect 18690 33572 18696 33584
rect 16669 33535 16727 33541
rect 16868 33544 17540 33572
rect 17880 33544 18696 33572
rect 15473 33507 15531 33513
rect 15473 33504 15485 33507
rect 15344 33476 15485 33504
rect 15344 33464 15350 33476
rect 15473 33473 15485 33476
rect 15519 33473 15531 33507
rect 15654 33504 15660 33516
rect 15615 33476 15660 33504
rect 15473 33467 15531 33473
rect 15654 33464 15660 33476
rect 15712 33464 15718 33516
rect 16868 33504 16896 33544
rect 16500 33476 16896 33504
rect 16945 33507 17003 33513
rect 14090 33396 14096 33448
rect 14148 33436 14154 33448
rect 14369 33439 14427 33445
rect 14369 33436 14381 33439
rect 14148 33408 14381 33436
rect 14148 33396 14154 33408
rect 14369 33405 14381 33408
rect 14415 33436 14427 33439
rect 16500 33436 16528 33476
rect 16945 33473 16957 33507
rect 16991 33504 17003 33507
rect 17880 33504 17908 33544
rect 18690 33532 18696 33544
rect 18748 33532 18754 33584
rect 19705 33575 19763 33581
rect 19705 33541 19717 33575
rect 19751 33572 19763 33575
rect 20070 33572 20076 33584
rect 19751 33544 20076 33572
rect 19751 33541 19763 33544
rect 19705 33535 19763 33541
rect 20070 33532 20076 33544
rect 20128 33532 20134 33584
rect 16991 33476 17908 33504
rect 17957 33507 18015 33513
rect 16991 33473 17003 33476
rect 16945 33467 17003 33473
rect 17957 33473 17969 33507
rect 18003 33504 18015 33507
rect 18046 33504 18052 33516
rect 18003 33476 18052 33504
rect 18003 33473 18015 33476
rect 17957 33467 18015 33473
rect 18046 33464 18052 33476
rect 18104 33464 18110 33516
rect 18138 33464 18144 33516
rect 18196 33504 18202 33516
rect 18322 33504 18328 33516
rect 18196 33476 18328 33504
rect 18196 33464 18202 33476
rect 18322 33464 18328 33476
rect 18380 33464 18386 33516
rect 18506 33464 18512 33516
rect 18564 33504 18570 33516
rect 19061 33507 19119 33513
rect 19061 33504 19073 33507
rect 18564 33476 19073 33504
rect 18564 33464 18570 33476
rect 19061 33473 19073 33476
rect 19107 33504 19119 33507
rect 20180 33504 20208 33612
rect 20993 33609 21005 33612
rect 21039 33609 21051 33643
rect 20993 33603 21051 33609
rect 21177 33643 21235 33649
rect 21177 33609 21189 33643
rect 21223 33640 21235 33643
rect 24118 33640 24124 33652
rect 21223 33612 24124 33640
rect 21223 33609 21235 33612
rect 21177 33603 21235 33609
rect 24118 33600 24124 33612
rect 24176 33600 24182 33652
rect 24305 33643 24363 33649
rect 24305 33609 24317 33643
rect 24351 33640 24363 33643
rect 24762 33640 24768 33652
rect 24351 33612 24768 33640
rect 24351 33609 24363 33612
rect 24305 33603 24363 33609
rect 24762 33600 24768 33612
rect 24820 33640 24826 33652
rect 24820 33612 25636 33640
rect 24820 33600 24826 33612
rect 20349 33575 20407 33581
rect 20349 33541 20361 33575
rect 20395 33572 20407 33575
rect 21082 33572 21088 33584
rect 20395 33544 21088 33572
rect 20395 33541 20407 33544
rect 20349 33535 20407 33541
rect 21082 33532 21088 33544
rect 21140 33532 21146 33584
rect 22278 33532 22284 33584
rect 22336 33572 22342 33584
rect 22373 33575 22431 33581
rect 22373 33572 22385 33575
rect 22336 33544 22385 33572
rect 22336 33532 22342 33544
rect 22373 33541 22385 33544
rect 22419 33572 22431 33575
rect 22462 33572 22468 33584
rect 22419 33544 22468 33572
rect 22419 33541 22431 33544
rect 22373 33535 22431 33541
rect 22462 33532 22468 33544
rect 22520 33532 22526 33584
rect 22925 33575 22983 33581
rect 22925 33541 22937 33575
rect 22971 33572 22983 33575
rect 24213 33575 24271 33581
rect 24213 33572 24225 33575
rect 22971 33544 24225 33572
rect 22971 33541 22983 33544
rect 22925 33535 22983 33541
rect 24213 33541 24225 33544
rect 24259 33572 24271 33575
rect 24259 33544 24900 33572
rect 24259 33541 24271 33544
rect 24213 33535 24271 33541
rect 19107 33476 20208 33504
rect 19107 33473 19119 33476
rect 19061 33467 19119 33473
rect 20530 33464 20536 33516
rect 20588 33504 20594 33516
rect 20809 33507 20867 33513
rect 20809 33504 20821 33507
rect 20588 33476 20821 33504
rect 20588 33464 20594 33476
rect 20809 33473 20821 33476
rect 20855 33473 20867 33507
rect 20809 33467 20867 33473
rect 20901 33507 20959 33513
rect 20901 33473 20913 33507
rect 20947 33473 20959 33507
rect 22830 33504 22836 33516
rect 22791 33476 22836 33504
rect 20901 33467 20959 33473
rect 18414 33436 18420 33448
rect 14415 33408 16528 33436
rect 16592 33408 18420 33436
rect 14415 33405 14427 33408
rect 14369 33399 14427 33405
rect 16592 33380 16620 33408
rect 18414 33396 18420 33408
rect 18472 33396 18478 33448
rect 18601 33439 18659 33445
rect 18601 33405 18613 33439
rect 18647 33405 18659 33439
rect 18601 33399 18659 33405
rect 16574 33368 16580 33380
rect 6886 33340 16580 33368
rect 16574 33328 16580 33340
rect 16632 33328 16638 33380
rect 16669 33371 16727 33377
rect 16669 33337 16681 33371
rect 16715 33368 16727 33371
rect 16758 33368 16764 33380
rect 16715 33340 16764 33368
rect 16715 33337 16727 33340
rect 16669 33331 16727 33337
rect 16758 33328 16764 33340
rect 16816 33328 16822 33380
rect 18616 33368 18644 33399
rect 18690 33396 18696 33448
rect 18748 33436 18754 33448
rect 18969 33439 19027 33445
rect 18969 33436 18981 33439
rect 18748 33408 18981 33436
rect 18748 33396 18754 33408
rect 18969 33405 18981 33408
rect 19015 33405 19027 33439
rect 18969 33399 19027 33405
rect 18874 33368 18880 33380
rect 18616 33340 18880 33368
rect 18874 33328 18880 33340
rect 18932 33328 18938 33380
rect 18984 33368 19012 33399
rect 19242 33396 19248 33448
rect 19300 33436 19306 33448
rect 20073 33439 20131 33445
rect 20073 33436 20085 33439
rect 19300 33408 20085 33436
rect 19300 33396 19306 33408
rect 20073 33405 20085 33408
rect 20119 33405 20131 33439
rect 20073 33399 20131 33405
rect 20162 33396 20168 33448
rect 20220 33436 20226 33448
rect 20916 33436 20944 33467
rect 22830 33464 22836 33476
rect 22888 33464 22894 33516
rect 23017 33507 23075 33513
rect 23017 33473 23029 33507
rect 23063 33504 23075 33507
rect 23106 33504 23112 33516
rect 23063 33476 23112 33504
rect 23063 33473 23075 33476
rect 23017 33467 23075 33473
rect 23106 33464 23112 33476
rect 23164 33464 23170 33516
rect 23474 33464 23480 33516
rect 23532 33504 23538 33516
rect 24121 33507 24179 33513
rect 24121 33504 24133 33507
rect 23532 33476 24133 33504
rect 23532 33464 23538 33476
rect 24121 33473 24133 33476
rect 24167 33473 24179 33507
rect 24121 33467 24179 33473
rect 24397 33507 24455 33513
rect 24397 33473 24409 33507
rect 24443 33504 24455 33507
rect 24762 33504 24768 33516
rect 24443 33476 24768 33504
rect 24443 33473 24455 33476
rect 24397 33467 24455 33473
rect 20220 33408 20944 33436
rect 21177 33439 21235 33445
rect 20220 33396 20226 33408
rect 21177 33405 21189 33439
rect 21223 33436 21235 33439
rect 23290 33436 23296 33448
rect 21223 33408 23296 33436
rect 21223 33405 21235 33408
rect 21177 33399 21235 33405
rect 21192 33368 21220 33399
rect 23290 33396 23296 33408
rect 23348 33396 23354 33448
rect 24136 33436 24164 33467
rect 24762 33464 24768 33476
rect 24820 33464 24826 33516
rect 24872 33513 24900 33544
rect 24857 33507 24915 33513
rect 24857 33473 24869 33507
rect 24903 33473 24915 33507
rect 24857 33467 24915 33473
rect 24949 33507 25007 33513
rect 24949 33473 24961 33507
rect 24995 33473 25007 33507
rect 24949 33467 25007 33473
rect 24964 33436 24992 33467
rect 25038 33464 25044 33516
rect 25096 33504 25102 33516
rect 25133 33507 25191 33513
rect 25133 33504 25145 33507
rect 25096 33476 25145 33504
rect 25096 33464 25102 33476
rect 25133 33473 25145 33476
rect 25179 33504 25191 33507
rect 25222 33504 25228 33516
rect 25179 33476 25228 33504
rect 25179 33473 25191 33476
rect 25133 33467 25191 33473
rect 25222 33464 25228 33476
rect 25280 33464 25286 33516
rect 25608 33513 25636 33612
rect 27614 33600 27620 33652
rect 27672 33640 27678 33652
rect 27890 33640 27896 33652
rect 27672 33612 27896 33640
rect 27672 33600 27678 33612
rect 27890 33600 27896 33612
rect 27948 33640 27954 33652
rect 28169 33643 28227 33649
rect 28169 33640 28181 33643
rect 27948 33612 28181 33640
rect 27948 33600 27954 33612
rect 28169 33609 28181 33612
rect 28215 33609 28227 33643
rect 28169 33603 28227 33609
rect 25593 33507 25651 33513
rect 25593 33473 25605 33507
rect 25639 33473 25651 33507
rect 25774 33504 25780 33516
rect 25735 33476 25780 33504
rect 25593 33467 25651 33473
rect 25774 33464 25780 33476
rect 25832 33464 25838 33516
rect 27338 33504 27344 33516
rect 27299 33476 27344 33504
rect 27338 33464 27344 33476
rect 27396 33464 27402 33516
rect 27430 33464 27436 33516
rect 27488 33504 27494 33516
rect 27706 33504 27712 33516
rect 27488 33476 27533 33504
rect 27667 33476 27712 33504
rect 27488 33464 27494 33476
rect 27706 33464 27712 33476
rect 27764 33464 27770 33516
rect 28184 33504 28212 33603
rect 28350 33600 28356 33652
rect 28408 33640 28414 33652
rect 28721 33643 28779 33649
rect 28721 33640 28733 33643
rect 28408 33612 28733 33640
rect 28408 33600 28414 33612
rect 28721 33609 28733 33612
rect 28767 33609 28779 33643
rect 28721 33603 28779 33609
rect 29733 33643 29791 33649
rect 29733 33609 29745 33643
rect 29779 33640 29791 33643
rect 29914 33640 29920 33652
rect 29779 33612 29920 33640
rect 29779 33609 29791 33612
rect 29733 33603 29791 33609
rect 28736 33572 28764 33603
rect 29914 33600 29920 33612
rect 29972 33600 29978 33652
rect 30834 33600 30840 33652
rect 30892 33640 30898 33652
rect 31297 33643 31355 33649
rect 31297 33640 31309 33643
rect 30892 33612 31309 33640
rect 30892 33600 30898 33612
rect 31297 33609 31309 33612
rect 31343 33609 31355 33643
rect 31297 33603 31355 33609
rect 31478 33600 31484 33652
rect 31536 33640 31542 33652
rect 31536 33612 33548 33640
rect 31536 33600 31542 33612
rect 31938 33572 31944 33584
rect 28736 33544 31944 33572
rect 31938 33532 31944 33544
rect 31996 33532 32002 33584
rect 33520 33572 33548 33612
rect 33594 33600 33600 33652
rect 33652 33640 33658 33652
rect 34241 33643 34299 33649
rect 34241 33640 34253 33643
rect 33652 33612 34253 33640
rect 33652 33600 33658 33612
rect 34241 33609 34253 33612
rect 34287 33609 34299 33643
rect 36170 33640 36176 33652
rect 36131 33612 36176 33640
rect 34241 33603 34299 33609
rect 36170 33600 36176 33612
rect 36228 33600 36234 33652
rect 36262 33600 36268 33652
rect 36320 33640 36326 33652
rect 37277 33643 37335 33649
rect 36320 33612 36584 33640
rect 36320 33600 36326 33612
rect 33689 33575 33747 33581
rect 33689 33572 33701 33575
rect 33520 33544 33701 33572
rect 33689 33541 33701 33544
rect 33735 33572 33747 33575
rect 34514 33572 34520 33584
rect 33735 33544 34520 33572
rect 33735 33541 33747 33544
rect 33689 33535 33747 33541
rect 34514 33532 34520 33544
rect 34572 33532 34578 33584
rect 35526 33572 35532 33584
rect 34624 33544 35532 33572
rect 29178 33504 29184 33516
rect 28184 33476 29184 33504
rect 29178 33464 29184 33476
rect 29236 33464 29242 33516
rect 30374 33504 30380 33516
rect 30335 33476 30380 33504
rect 30374 33464 30380 33476
rect 30432 33464 30438 33516
rect 31205 33507 31263 33513
rect 31205 33473 31217 33507
rect 31251 33504 31263 33507
rect 31294 33504 31300 33516
rect 31251 33476 31300 33504
rect 31251 33473 31263 33476
rect 31205 33467 31263 33473
rect 31294 33464 31300 33476
rect 31352 33464 31358 33516
rect 31386 33464 31392 33516
rect 31444 33504 31450 33516
rect 32309 33507 32367 33513
rect 31444 33476 31489 33504
rect 31444 33464 31450 33476
rect 32309 33473 32321 33507
rect 32355 33473 32367 33507
rect 32309 33467 32367 33473
rect 24136 33408 24992 33436
rect 26970 33396 26976 33448
rect 27028 33436 27034 33448
rect 27525 33439 27583 33445
rect 27525 33436 27537 33439
rect 27028 33408 27537 33436
rect 27028 33396 27034 33408
rect 27525 33405 27537 33408
rect 27571 33405 27583 33439
rect 30466 33436 30472 33448
rect 30427 33408 30472 33436
rect 27525 33399 27583 33405
rect 30466 33396 30472 33408
rect 30524 33396 30530 33448
rect 30558 33396 30564 33448
rect 30616 33436 30622 33448
rect 30745 33439 30803 33445
rect 30745 33436 30757 33439
rect 30616 33408 30757 33436
rect 30616 33396 30622 33408
rect 30745 33405 30757 33408
rect 30791 33405 30803 33439
rect 30745 33399 30803 33405
rect 32122 33396 32128 33448
rect 32180 33436 32186 33448
rect 32324 33436 32352 33467
rect 32398 33464 32404 33516
rect 32456 33504 32462 33516
rect 32582 33504 32588 33516
rect 32456 33476 32501 33504
rect 32543 33476 32588 33504
rect 32456 33464 32462 33476
rect 32582 33464 32588 33476
rect 32640 33464 32646 33516
rect 34624 33513 34652 33544
rect 35526 33532 35532 33544
rect 35584 33532 35590 33584
rect 35621 33575 35679 33581
rect 35621 33541 35633 33575
rect 35667 33572 35679 33575
rect 36446 33572 36452 33584
rect 35667 33544 36452 33572
rect 35667 33541 35679 33544
rect 35621 33535 35679 33541
rect 36446 33532 36452 33544
rect 36504 33532 36510 33584
rect 36556 33572 36584 33612
rect 37277 33609 37289 33643
rect 37323 33640 37335 33643
rect 37550 33640 37556 33652
rect 37323 33612 37556 33640
rect 37323 33609 37335 33612
rect 37277 33603 37335 33609
rect 37550 33600 37556 33612
rect 37608 33600 37614 33652
rect 38654 33640 38660 33652
rect 38615 33612 38660 33640
rect 38654 33600 38660 33612
rect 38712 33600 38718 33652
rect 41046 33640 41052 33652
rect 40512 33612 41052 33640
rect 37645 33575 37703 33581
rect 36556 33544 37596 33572
rect 34609 33507 34667 33513
rect 34609 33473 34621 33507
rect 34655 33473 34667 33507
rect 34609 33467 34667 33473
rect 35437 33507 35495 33513
rect 35437 33473 35449 33507
rect 35483 33504 35495 33507
rect 36081 33507 36139 33513
rect 35483 33476 35664 33504
rect 35483 33473 35495 33476
rect 35437 33467 35495 33473
rect 35636 33448 35664 33476
rect 36081 33473 36093 33507
rect 36127 33504 36139 33507
rect 36170 33504 36176 33516
rect 36127 33476 36176 33504
rect 36127 33473 36139 33476
rect 36081 33467 36139 33473
rect 36170 33464 36176 33476
rect 36228 33464 36234 33516
rect 37568 33513 37596 33544
rect 37645 33541 37657 33575
rect 37691 33572 37703 33575
rect 38378 33572 38384 33584
rect 37691 33544 38384 33572
rect 37691 33541 37703 33544
rect 37645 33535 37703 33541
rect 38378 33532 38384 33544
rect 38436 33572 38442 33584
rect 38473 33575 38531 33581
rect 38473 33572 38485 33575
rect 38436 33544 38485 33572
rect 38436 33532 38442 33544
rect 38473 33541 38485 33544
rect 38519 33541 38531 33575
rect 38473 33535 38531 33541
rect 39485 33575 39543 33581
rect 39485 33541 39497 33575
rect 39531 33572 39543 33575
rect 40402 33572 40408 33584
rect 39531 33544 40408 33572
rect 39531 33541 39543 33544
rect 39485 33535 39543 33541
rect 40402 33532 40408 33544
rect 40460 33532 40466 33584
rect 36265 33507 36323 33513
rect 36265 33473 36277 33507
rect 36311 33504 36323 33507
rect 37461 33507 37519 33513
rect 37461 33504 37473 33507
rect 36311 33476 37473 33504
rect 36311 33473 36323 33476
rect 36265 33467 36323 33473
rect 37461 33473 37473 33476
rect 37507 33473 37519 33507
rect 37461 33467 37519 33473
rect 37553 33507 37611 33513
rect 37553 33473 37565 33507
rect 37599 33473 37611 33507
rect 37553 33467 37611 33473
rect 32950 33436 32956 33448
rect 32180 33408 32956 33436
rect 32180 33396 32186 33408
rect 32950 33396 32956 33408
rect 33008 33396 33014 33448
rect 34514 33436 34520 33448
rect 34475 33408 34520 33436
rect 34514 33396 34520 33408
rect 34572 33396 34578 33448
rect 35253 33439 35311 33445
rect 35253 33405 35265 33439
rect 35299 33405 35311 33439
rect 35253 33399 35311 33405
rect 18984 33340 21220 33368
rect 21266 33328 21272 33380
rect 21324 33368 21330 33380
rect 23569 33371 23627 33377
rect 23569 33368 23581 33371
rect 21324 33340 23581 33368
rect 21324 33328 21330 33340
rect 23569 33337 23581 33340
rect 23615 33368 23627 33371
rect 24210 33368 24216 33380
rect 23615 33340 24216 33368
rect 23615 33337 23627 33340
rect 23569 33331 23627 33337
rect 24210 33328 24216 33340
rect 24268 33368 24274 33380
rect 24762 33368 24768 33380
rect 24268 33340 24768 33368
rect 24268 33328 24274 33340
rect 24762 33328 24768 33340
rect 24820 33328 24826 33380
rect 25130 33368 25136 33380
rect 25091 33340 25136 33368
rect 25130 33328 25136 33340
rect 25188 33328 25194 33380
rect 27709 33371 27767 33377
rect 27709 33337 27721 33371
rect 27755 33368 27767 33371
rect 34330 33368 34336 33380
rect 27755 33340 34336 33368
rect 27755 33337 27767 33340
rect 27709 33331 27767 33337
rect 34330 33328 34336 33340
rect 34388 33328 34394 33380
rect 35268 33368 35296 33399
rect 35618 33396 35624 33448
rect 35676 33436 35682 33448
rect 36280 33436 36308 33467
rect 35676 33408 36308 33436
rect 35676 33396 35682 33408
rect 36170 33368 36176 33380
rect 35268 33340 36176 33368
rect 36170 33328 36176 33340
rect 36228 33328 36234 33380
rect 37476 33368 37504 33467
rect 37568 33436 37596 33467
rect 37734 33464 37740 33516
rect 37792 33504 37798 33516
rect 37829 33507 37887 33513
rect 37829 33504 37841 33507
rect 37792 33476 37841 33504
rect 37792 33464 37798 33476
rect 37829 33473 37841 33476
rect 37875 33504 37887 33507
rect 38102 33504 38108 33516
rect 37875 33476 38108 33504
rect 37875 33473 37887 33476
rect 37829 33467 37887 33473
rect 38102 33464 38108 33476
rect 38160 33504 38166 33516
rect 38289 33507 38347 33513
rect 38289 33504 38301 33507
rect 38160 33476 38301 33504
rect 38160 33464 38166 33476
rect 38289 33473 38301 33476
rect 38335 33473 38347 33507
rect 39114 33504 39120 33516
rect 39075 33476 39120 33504
rect 38289 33467 38347 33473
rect 39114 33464 39120 33476
rect 39172 33464 39178 33516
rect 39298 33504 39304 33516
rect 39259 33476 39304 33504
rect 39298 33464 39304 33476
rect 39356 33464 39362 33516
rect 39574 33504 39580 33516
rect 39535 33476 39580 33504
rect 39574 33464 39580 33476
rect 39632 33464 39638 33516
rect 39945 33507 40003 33513
rect 39945 33473 39957 33507
rect 39991 33504 40003 33507
rect 40126 33504 40132 33516
rect 39991 33476 40132 33504
rect 39991 33473 40003 33476
rect 39945 33467 40003 33473
rect 40126 33464 40132 33476
rect 40184 33504 40190 33516
rect 40512 33504 40540 33612
rect 41046 33600 41052 33612
rect 41104 33600 41110 33652
rect 48130 33640 48136 33652
rect 48091 33612 48136 33640
rect 48130 33600 48136 33612
rect 48188 33600 48194 33652
rect 42981 33575 43039 33581
rect 42981 33572 42993 33575
rect 40972 33544 42993 33572
rect 40678 33504 40684 33516
rect 40184 33476 40540 33504
rect 40639 33476 40684 33504
rect 40184 33464 40190 33476
rect 40678 33464 40684 33476
rect 40736 33464 40742 33516
rect 40770 33507 40828 33513
rect 40770 33473 40782 33507
rect 40816 33473 40828 33507
rect 40770 33467 40828 33473
rect 38010 33436 38016 33448
rect 37568 33408 38016 33436
rect 38010 33396 38016 33408
rect 38068 33436 38074 33448
rect 40034 33436 40040 33448
rect 38068 33408 40040 33436
rect 38068 33396 38074 33408
rect 40034 33396 40040 33408
rect 40092 33396 40098 33448
rect 39850 33368 39856 33380
rect 37476 33340 39856 33368
rect 39850 33328 39856 33340
rect 39908 33328 39914 33380
rect 40785 33312 40813 33467
rect 40862 33464 40868 33516
rect 40920 33504 40926 33516
rect 40972 33504 41000 33544
rect 42981 33541 42993 33544
rect 43027 33572 43039 33575
rect 43070 33572 43076 33584
rect 43027 33544 43076 33572
rect 43027 33541 43039 33544
rect 42981 33535 43039 33541
rect 43070 33532 43076 33544
rect 43128 33532 43134 33584
rect 40920 33476 41000 33504
rect 40920 33464 40926 33476
rect 41046 33464 41052 33516
rect 41104 33504 41110 33516
rect 47854 33504 47860 33516
rect 41104 33476 47860 33504
rect 41104 33464 41110 33476
rect 47854 33464 47860 33476
rect 47912 33464 47918 33516
rect 41414 33328 41420 33380
rect 41472 33368 41478 33380
rect 41509 33371 41567 33377
rect 41509 33368 41521 33371
rect 41472 33340 41521 33368
rect 41472 33328 41478 33340
rect 41509 33337 41521 33340
rect 41555 33337 41567 33371
rect 41509 33331 41567 33337
rect 12710 33260 12716 33312
rect 12768 33300 12774 33312
rect 13081 33303 13139 33309
rect 13081 33300 13093 33303
rect 12768 33272 13093 33300
rect 12768 33260 12774 33272
rect 13081 33269 13093 33272
rect 13127 33269 13139 33303
rect 13081 33263 13139 33269
rect 15013 33303 15071 33309
rect 15013 33269 15025 33303
rect 15059 33300 15071 33303
rect 15562 33300 15568 33312
rect 15059 33272 15568 33300
rect 15059 33269 15071 33272
rect 15013 33263 15071 33269
rect 15562 33260 15568 33272
rect 15620 33260 15626 33312
rect 18049 33303 18107 33309
rect 18049 33269 18061 33303
rect 18095 33300 18107 33303
rect 18138 33300 18144 33312
rect 18095 33272 18144 33300
rect 18095 33269 18107 33272
rect 18049 33263 18107 33269
rect 18138 33260 18144 33272
rect 18196 33260 18202 33312
rect 25682 33300 25688 33312
rect 25643 33272 25688 33300
rect 25682 33260 25688 33272
rect 25740 33260 25746 33312
rect 26421 33303 26479 33309
rect 26421 33269 26433 33303
rect 26467 33300 26479 33303
rect 27154 33300 27160 33312
rect 26467 33272 27160 33300
rect 26467 33269 26479 33272
rect 26421 33263 26479 33269
rect 27154 33260 27160 33272
rect 27212 33260 27218 33312
rect 29914 33260 29920 33312
rect 29972 33300 29978 33312
rect 31478 33300 31484 33312
rect 29972 33272 31484 33300
rect 29972 33260 29978 33272
rect 31478 33260 31484 33272
rect 31536 33260 31542 33312
rect 32214 33260 32220 33312
rect 32272 33300 32278 33312
rect 32585 33303 32643 33309
rect 32585 33300 32597 33303
rect 32272 33272 32597 33300
rect 32272 33260 32278 33272
rect 32585 33269 32597 33272
rect 32631 33269 32643 33303
rect 32585 33263 32643 33269
rect 33137 33303 33195 33309
rect 33137 33269 33149 33303
rect 33183 33300 33195 33303
rect 33226 33300 33232 33312
rect 33183 33272 33232 33300
rect 33183 33269 33195 33272
rect 33137 33263 33195 33269
rect 33226 33260 33232 33272
rect 33284 33260 33290 33312
rect 34422 33260 34428 33312
rect 34480 33300 34486 33312
rect 34517 33303 34575 33309
rect 34517 33300 34529 33303
rect 34480 33272 34529 33300
rect 34480 33260 34486 33272
rect 34517 33269 34529 33272
rect 34563 33269 34575 33303
rect 40402 33300 40408 33312
rect 40363 33272 40408 33300
rect 34517 33263 34575 33269
rect 40402 33260 40408 33272
rect 40460 33260 40466 33312
rect 40770 33260 40776 33312
rect 40828 33260 40834 33312
rect 40862 33260 40868 33312
rect 40920 33300 40926 33312
rect 42429 33303 42487 33309
rect 42429 33300 42441 33303
rect 40920 33272 42441 33300
rect 40920 33260 40926 33272
rect 42429 33269 42441 33272
rect 42475 33269 42487 33303
rect 42429 33263 42487 33269
rect 43162 33260 43168 33312
rect 43220 33300 43226 33312
rect 43625 33303 43683 33309
rect 43625 33300 43637 33303
rect 43220 33272 43637 33300
rect 43220 33260 43226 33272
rect 43625 33269 43637 33272
rect 43671 33300 43683 33303
rect 44174 33300 44180 33312
rect 43671 33272 44180 33300
rect 43671 33269 43683 33272
rect 43625 33263 43683 33269
rect 44174 33260 44180 33272
rect 44232 33260 44238 33312
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 11606 33096 11612 33108
rect 11567 33068 11612 33096
rect 11606 33056 11612 33068
rect 11664 33056 11670 33108
rect 12434 33056 12440 33108
rect 12492 33096 12498 33108
rect 12621 33099 12679 33105
rect 12621 33096 12633 33099
rect 12492 33068 12633 33096
rect 12492 33056 12498 33068
rect 12621 33065 12633 33068
rect 12667 33065 12679 33099
rect 12621 33059 12679 33065
rect 14921 33099 14979 33105
rect 14921 33065 14933 33099
rect 14967 33096 14979 33099
rect 17126 33096 17132 33108
rect 14967 33068 17132 33096
rect 14967 33065 14979 33068
rect 14921 33059 14979 33065
rect 17126 33056 17132 33068
rect 17184 33096 17190 33108
rect 17862 33096 17868 33108
rect 17184 33068 17868 33096
rect 17184 33056 17190 33068
rect 17862 33056 17868 33068
rect 17920 33056 17926 33108
rect 20162 33096 20168 33108
rect 20123 33068 20168 33096
rect 20162 33056 20168 33068
rect 20220 33056 20226 33108
rect 20714 33096 20720 33108
rect 20675 33068 20720 33096
rect 20714 33056 20720 33068
rect 20772 33056 20778 33108
rect 22186 33056 22192 33108
rect 22244 33096 22250 33108
rect 22465 33099 22523 33105
rect 22465 33096 22477 33099
rect 22244 33068 22477 33096
rect 22244 33056 22250 33068
rect 22465 33065 22477 33068
rect 22511 33065 22523 33099
rect 22830 33096 22836 33108
rect 22791 33068 22836 33096
rect 22465 33059 22523 33065
rect 22830 33056 22836 33068
rect 22888 33056 22894 33108
rect 22922 33056 22928 33108
rect 22980 33096 22986 33108
rect 23382 33096 23388 33108
rect 22980 33068 23388 33096
rect 22980 33056 22986 33068
rect 23382 33056 23388 33068
rect 23440 33056 23446 33108
rect 24857 33099 24915 33105
rect 24857 33065 24869 33099
rect 24903 33096 24915 33099
rect 25774 33096 25780 33108
rect 24903 33068 25780 33096
rect 24903 33065 24915 33068
rect 24857 33059 24915 33065
rect 25774 33056 25780 33068
rect 25832 33056 25838 33108
rect 27522 33056 27528 33108
rect 27580 33096 27586 33108
rect 28442 33096 28448 33108
rect 27580 33068 28448 33096
rect 27580 33056 27586 33068
rect 28442 33056 28448 33068
rect 28500 33096 28506 33108
rect 29638 33096 29644 33108
rect 28500 33068 29644 33096
rect 28500 33056 28506 33068
rect 29638 33056 29644 33068
rect 29696 33056 29702 33108
rect 30285 33099 30343 33105
rect 30285 33065 30297 33099
rect 30331 33096 30343 33099
rect 30466 33096 30472 33108
rect 30331 33068 30472 33096
rect 30331 33065 30343 33068
rect 30285 33059 30343 33065
rect 30466 33056 30472 33068
rect 30524 33056 30530 33108
rect 33134 33096 33140 33108
rect 32600 33068 33140 33096
rect 16301 33031 16359 33037
rect 16301 32997 16313 33031
rect 16347 33028 16359 33031
rect 18874 33028 18880 33040
rect 16347 33000 18880 33028
rect 16347 32997 16359 33000
rect 16301 32991 16359 32997
rect 18874 32988 18880 33000
rect 18932 32988 18938 33040
rect 23290 32988 23296 33040
rect 23348 33028 23354 33040
rect 25961 33031 26019 33037
rect 23348 33000 25820 33028
rect 23348 32988 23354 33000
rect 10505 32963 10563 32969
rect 10505 32929 10517 32963
rect 10551 32960 10563 32963
rect 10551 32932 11744 32960
rect 10551 32929 10563 32932
rect 10505 32923 10563 32929
rect 11716 32904 11744 32932
rect 11974 32920 11980 32972
rect 12032 32960 12038 32972
rect 15746 32960 15752 32972
rect 12032 32932 14412 32960
rect 12032 32920 12038 32932
rect 11514 32892 11520 32904
rect 11475 32864 11520 32892
rect 11514 32852 11520 32864
rect 11572 32852 11578 32904
rect 11698 32892 11704 32904
rect 11659 32864 11704 32892
rect 11698 32852 11704 32864
rect 11756 32852 11762 32904
rect 12802 32892 12808 32904
rect 12763 32864 12808 32892
rect 12802 32852 12808 32864
rect 12860 32852 12866 32904
rect 12897 32895 12955 32901
rect 12897 32861 12909 32895
rect 12943 32861 12955 32895
rect 12897 32855 12955 32861
rect 12912 32824 12940 32855
rect 12986 32852 12992 32904
rect 13044 32892 13050 32904
rect 13081 32895 13139 32901
rect 13081 32892 13093 32895
rect 13044 32864 13093 32892
rect 13044 32852 13050 32864
rect 13081 32861 13093 32864
rect 13127 32861 13139 32895
rect 13081 32855 13139 32861
rect 13173 32895 13231 32901
rect 13173 32861 13185 32895
rect 13219 32892 13231 32895
rect 13814 32892 13820 32904
rect 13219 32864 13820 32892
rect 13219 32861 13231 32864
rect 13173 32855 13231 32861
rect 13814 32852 13820 32864
rect 13872 32852 13878 32904
rect 13446 32824 13452 32836
rect 12912 32796 13452 32824
rect 13446 32784 13452 32796
rect 13504 32784 13510 32836
rect 11057 32759 11115 32765
rect 11057 32725 11069 32759
rect 11103 32756 11115 32759
rect 13170 32756 13176 32768
rect 11103 32728 13176 32756
rect 11103 32725 11115 32728
rect 11057 32719 11115 32725
rect 13170 32716 13176 32728
rect 13228 32716 13234 32768
rect 14384 32765 14412 32932
rect 15396 32932 15752 32960
rect 15286 32852 15292 32904
rect 15344 32892 15350 32904
rect 15396 32901 15424 32932
rect 15746 32920 15752 32932
rect 15804 32920 15810 32972
rect 19334 32920 19340 32972
rect 19392 32960 19398 32972
rect 19797 32963 19855 32969
rect 19797 32960 19809 32963
rect 19392 32932 19809 32960
rect 19392 32920 19398 32932
rect 19797 32929 19809 32932
rect 19843 32929 19855 32963
rect 19797 32923 19855 32929
rect 21821 32963 21879 32969
rect 21821 32929 21833 32963
rect 21867 32960 21879 32963
rect 25682 32960 25688 32972
rect 21867 32932 23152 32960
rect 25643 32932 25688 32960
rect 21867 32929 21879 32932
rect 21821 32923 21879 32929
rect 23124 32904 23152 32932
rect 25682 32920 25688 32932
rect 25740 32920 25746 32972
rect 25792 32960 25820 33000
rect 25961 32997 25973 33031
rect 26007 33028 26019 33031
rect 26786 33028 26792 33040
rect 26007 33000 26792 33028
rect 26007 32997 26019 33000
rect 25961 32991 26019 32997
rect 26786 32988 26792 33000
rect 26844 32988 26850 33040
rect 31110 32988 31116 33040
rect 31168 33028 31174 33040
rect 31205 33031 31263 33037
rect 31205 33028 31217 33031
rect 31168 33000 31217 33028
rect 31168 32988 31174 33000
rect 31205 32997 31217 33000
rect 31251 32997 31263 33031
rect 32309 33031 32367 33037
rect 32309 33028 32321 33031
rect 31205 32991 31263 32997
rect 31312 33000 32321 33028
rect 31312 32960 31340 33000
rect 32309 32997 32321 33000
rect 32355 32997 32367 33031
rect 32309 32991 32367 32997
rect 25792 32932 31340 32960
rect 31665 32963 31723 32969
rect 31665 32929 31677 32963
rect 31711 32960 31723 32963
rect 32122 32960 32128 32972
rect 31711 32932 32128 32960
rect 31711 32929 31723 32932
rect 31665 32923 31723 32929
rect 32122 32920 32128 32932
rect 32180 32920 32186 32972
rect 15381 32895 15439 32901
rect 15381 32892 15393 32895
rect 15344 32864 15393 32892
rect 15344 32852 15350 32864
rect 15381 32861 15393 32864
rect 15427 32861 15439 32895
rect 15562 32892 15568 32904
rect 15523 32864 15568 32892
rect 15381 32855 15439 32861
rect 15562 32852 15568 32864
rect 15620 32852 15626 32904
rect 15930 32892 15936 32904
rect 15891 32864 15936 32892
rect 15930 32852 15936 32864
rect 15988 32852 15994 32904
rect 16117 32895 16175 32901
rect 16117 32861 16129 32895
rect 16163 32861 16175 32895
rect 16117 32855 16175 32861
rect 16393 32895 16451 32901
rect 16393 32861 16405 32895
rect 16439 32892 16451 32895
rect 16666 32892 16672 32904
rect 16439 32864 16672 32892
rect 16439 32861 16451 32864
rect 16393 32855 16451 32861
rect 16132 32824 16160 32855
rect 16666 32852 16672 32864
rect 16724 32852 16730 32904
rect 17034 32892 17040 32904
rect 16995 32864 17040 32892
rect 17034 32852 17040 32864
rect 17092 32852 17098 32904
rect 17310 32892 17316 32904
rect 17271 32864 17316 32892
rect 17310 32852 17316 32864
rect 17368 32852 17374 32904
rect 17494 32892 17500 32904
rect 17455 32864 17500 32892
rect 17494 32852 17500 32864
rect 17552 32852 17558 32904
rect 17954 32892 17960 32904
rect 17915 32864 17960 32892
rect 17954 32852 17960 32864
rect 18012 32852 18018 32904
rect 18138 32892 18144 32904
rect 18099 32864 18144 32892
rect 18138 32852 18144 32864
rect 18196 32852 18202 32904
rect 19978 32892 19984 32904
rect 19939 32864 19984 32892
rect 19978 32852 19984 32864
rect 20036 32852 20042 32904
rect 20438 32852 20444 32904
rect 20496 32892 20502 32904
rect 20717 32895 20775 32901
rect 20717 32892 20729 32895
rect 20496 32864 20729 32892
rect 20496 32852 20502 32864
rect 20717 32861 20729 32864
rect 20763 32861 20775 32895
rect 20717 32855 20775 32861
rect 20901 32895 20959 32901
rect 20901 32861 20913 32895
rect 20947 32892 20959 32895
rect 20990 32892 20996 32904
rect 20947 32864 20996 32892
rect 20947 32861 20959 32864
rect 20901 32855 20959 32861
rect 20990 32852 20996 32864
rect 21048 32852 21054 32904
rect 21726 32892 21732 32904
rect 21784 32901 21790 32904
rect 21652 32864 21732 32892
rect 16853 32827 16911 32833
rect 16853 32824 16865 32827
rect 16132 32796 16865 32824
rect 16853 32793 16865 32796
rect 16899 32793 16911 32827
rect 16853 32787 16911 32793
rect 18693 32827 18751 32833
rect 18693 32793 18705 32827
rect 18739 32824 18751 32827
rect 21652 32824 21680 32864
rect 21726 32852 21732 32864
rect 21784 32892 21793 32901
rect 21910 32892 21916 32904
rect 21784 32864 21829 32892
rect 21871 32864 21916 32892
rect 21784 32855 21793 32864
rect 21784 32852 21790 32855
rect 21910 32852 21916 32864
rect 21968 32852 21974 32904
rect 22370 32892 22376 32904
rect 22331 32864 22376 32892
rect 22370 32852 22376 32864
rect 22428 32852 22434 32904
rect 22646 32892 22652 32904
rect 22607 32864 22652 32892
rect 22646 32852 22652 32864
rect 22704 32852 22710 32904
rect 23106 32852 23112 32904
rect 23164 32892 23170 32904
rect 23293 32895 23351 32901
rect 23293 32892 23305 32895
rect 23164 32864 23305 32892
rect 23164 32852 23170 32864
rect 23293 32861 23305 32864
rect 23339 32861 23351 32895
rect 23474 32892 23480 32904
rect 23435 32864 23480 32892
rect 23293 32855 23351 32861
rect 23474 32852 23480 32864
rect 23532 32852 23538 32904
rect 24762 32892 24768 32904
rect 24723 32864 24768 32892
rect 24762 32852 24768 32864
rect 24820 32852 24826 32904
rect 24854 32852 24860 32904
rect 24912 32892 24918 32904
rect 24949 32895 25007 32901
rect 24949 32892 24961 32895
rect 24912 32864 24961 32892
rect 24912 32852 24918 32864
rect 24949 32861 24961 32864
rect 24995 32892 25007 32895
rect 25498 32892 25504 32904
rect 24995 32864 25504 32892
rect 24995 32861 25007 32864
rect 24949 32855 25007 32861
rect 25498 32852 25504 32864
rect 25556 32852 25562 32904
rect 25593 32895 25651 32901
rect 25593 32861 25605 32895
rect 25639 32892 25651 32895
rect 25958 32892 25964 32904
rect 25639 32864 25964 32892
rect 25639 32861 25651 32864
rect 25593 32855 25651 32861
rect 25958 32852 25964 32864
rect 26016 32852 26022 32904
rect 26694 32892 26700 32904
rect 26655 32864 26700 32892
rect 26694 32852 26700 32864
rect 26752 32852 26758 32904
rect 26881 32895 26939 32901
rect 26881 32861 26893 32895
rect 26927 32892 26939 32895
rect 26927 32864 27016 32892
rect 26927 32861 26939 32864
rect 26881 32855 26939 32861
rect 18739 32796 21680 32824
rect 18739 32793 18751 32796
rect 18693 32787 18751 32793
rect 21818 32784 21824 32836
rect 21876 32824 21882 32836
rect 26602 32824 26608 32836
rect 21876 32796 26608 32824
rect 21876 32784 21882 32796
rect 26602 32784 26608 32796
rect 26660 32784 26666 32836
rect 26988 32824 27016 32864
rect 27062 32852 27068 32904
rect 27120 32892 27126 32904
rect 27525 32895 27583 32901
rect 27525 32892 27537 32895
rect 27120 32864 27537 32892
rect 27120 32852 27126 32864
rect 27525 32861 27537 32864
rect 27571 32861 27583 32895
rect 28350 32892 28356 32904
rect 28311 32864 28356 32892
rect 27525 32855 27583 32861
rect 28350 32852 28356 32864
rect 28408 32852 28414 32904
rect 28537 32895 28595 32901
rect 28537 32861 28549 32895
rect 28583 32861 28595 32895
rect 28537 32855 28595 32861
rect 27341 32827 27399 32833
rect 27341 32824 27353 32827
rect 26988 32796 27353 32824
rect 27341 32793 27353 32796
rect 27387 32824 27399 32827
rect 27890 32824 27896 32836
rect 27387 32796 27896 32824
rect 27387 32793 27399 32796
rect 27341 32787 27399 32793
rect 27890 32784 27896 32796
rect 27948 32784 27954 32836
rect 14369 32759 14427 32765
rect 14369 32725 14381 32759
rect 14415 32756 14427 32759
rect 14734 32756 14740 32768
rect 14415 32728 14740 32756
rect 14415 32725 14427 32728
rect 14369 32719 14427 32725
rect 14734 32716 14740 32728
rect 14792 32716 14798 32768
rect 18046 32756 18052 32768
rect 18007 32728 18052 32756
rect 18046 32716 18052 32728
rect 18104 32716 18110 32768
rect 18782 32716 18788 32768
rect 18840 32756 18846 32768
rect 19337 32759 19395 32765
rect 19337 32756 19349 32759
rect 18840 32728 19349 32756
rect 18840 32716 18846 32728
rect 19337 32725 19349 32728
rect 19383 32756 19395 32759
rect 22278 32756 22284 32768
rect 19383 32728 22284 32756
rect 19383 32725 19395 32728
rect 19337 32719 19395 32725
rect 22278 32716 22284 32728
rect 22336 32716 22342 32768
rect 26789 32759 26847 32765
rect 26789 32725 26801 32759
rect 26835 32756 26847 32759
rect 27614 32756 27620 32768
rect 26835 32728 27620 32756
rect 26835 32725 26847 32728
rect 26789 32719 26847 32725
rect 27614 32716 27620 32728
rect 27672 32716 27678 32768
rect 27709 32759 27767 32765
rect 27709 32725 27721 32759
rect 27755 32756 27767 32759
rect 27798 32756 27804 32768
rect 27755 32728 27804 32756
rect 27755 32725 27767 32728
rect 27709 32719 27767 32725
rect 27798 32716 27804 32728
rect 27856 32756 27862 32768
rect 28552 32756 28580 32855
rect 29546 32852 29552 32904
rect 29604 32892 29610 32904
rect 30282 32892 30288 32904
rect 29604 32864 30288 32892
rect 29604 32852 29610 32864
rect 30282 32852 30288 32864
rect 30340 32892 30346 32904
rect 30469 32895 30527 32901
rect 30469 32892 30481 32895
rect 30340 32864 30481 32892
rect 30340 32852 30346 32864
rect 30469 32861 30481 32864
rect 30515 32861 30527 32895
rect 30469 32855 30527 32861
rect 30558 32852 30564 32904
rect 30616 32892 30622 32904
rect 32600 32901 32628 33068
rect 33134 33056 33140 33068
rect 33192 33056 33198 33108
rect 33505 33099 33563 33105
rect 33505 33065 33517 33099
rect 33551 33096 33563 33099
rect 34054 33096 34060 33108
rect 33551 33068 34060 33096
rect 33551 33065 33563 33068
rect 33505 33059 33563 33065
rect 34054 33056 34060 33068
rect 34112 33056 34118 33108
rect 36078 33056 36084 33108
rect 36136 33096 36142 33108
rect 36173 33099 36231 33105
rect 36173 33096 36185 33099
rect 36136 33068 36185 33096
rect 36136 33056 36142 33068
rect 36173 33065 36185 33068
rect 36219 33096 36231 33099
rect 36725 33099 36783 33105
rect 36725 33096 36737 33099
rect 36219 33068 36737 33096
rect 36219 33065 36231 33068
rect 36173 33059 36231 33065
rect 36725 33065 36737 33068
rect 36771 33065 36783 33099
rect 36725 33059 36783 33065
rect 37366 33056 37372 33108
rect 37424 33096 37430 33108
rect 37461 33099 37519 33105
rect 37461 33096 37473 33099
rect 37424 33068 37473 33096
rect 37424 33056 37430 33068
rect 37461 33065 37473 33068
rect 37507 33065 37519 33099
rect 37461 33059 37519 33065
rect 37918 33056 37924 33108
rect 37976 33096 37982 33108
rect 38105 33099 38163 33105
rect 38105 33096 38117 33099
rect 37976 33068 38117 33096
rect 37976 33056 37982 33068
rect 38105 33065 38117 33068
rect 38151 33065 38163 33099
rect 38105 33059 38163 33065
rect 40034 33056 40040 33108
rect 40092 33096 40098 33108
rect 40862 33096 40868 33108
rect 40092 33068 40868 33096
rect 40092 33056 40098 33068
rect 40862 33056 40868 33068
rect 40920 33056 40926 33108
rect 32674 32988 32680 33040
rect 32732 33028 32738 33040
rect 32732 33000 33732 33028
rect 32732 32988 32738 33000
rect 31573 32895 31631 32901
rect 30616 32864 30661 32892
rect 30616 32852 30622 32864
rect 31573 32861 31585 32895
rect 31619 32892 31631 32895
rect 32493 32895 32551 32901
rect 31619 32864 31754 32892
rect 31619 32861 31631 32864
rect 31573 32855 31631 32861
rect 31726 32824 31754 32864
rect 32493 32861 32505 32895
rect 32539 32861 32551 32895
rect 32493 32855 32551 32861
rect 32585 32895 32643 32901
rect 32585 32861 32597 32895
rect 32631 32861 32643 32895
rect 32766 32892 32772 32904
rect 32727 32864 32772 32892
rect 32585 32855 32643 32861
rect 32398 32824 32404 32836
rect 31726 32796 32404 32824
rect 32398 32784 32404 32796
rect 32456 32784 32462 32836
rect 32508 32824 32536 32855
rect 32766 32852 32772 32864
rect 32824 32852 32830 32904
rect 32858 32852 32864 32904
rect 32916 32892 32922 32904
rect 32916 32864 32961 32892
rect 32916 32852 32922 32864
rect 33459 32861 33517 32867
rect 33459 32836 33471 32861
rect 32508 32796 33364 32824
rect 27856 32728 28580 32756
rect 28721 32759 28779 32765
rect 27856 32716 27862 32728
rect 28721 32725 28733 32759
rect 28767 32756 28779 32759
rect 28810 32756 28816 32768
rect 28767 32728 28816 32756
rect 28767 32725 28779 32728
rect 28721 32719 28779 32725
rect 28810 32716 28816 32728
rect 28868 32716 28874 32768
rect 29638 32756 29644 32768
rect 29551 32728 29644 32756
rect 29638 32716 29644 32728
rect 29696 32756 29702 32768
rect 30834 32756 30840 32768
rect 29696 32728 30840 32756
rect 29696 32716 29702 32728
rect 30834 32716 30840 32728
rect 30892 32716 30898 32768
rect 33336 32765 33364 32796
rect 33410 32784 33416 32836
rect 33468 32827 33471 32836
rect 33505 32858 33517 32861
rect 33505 32827 33532 32858
rect 33704 32833 33732 33000
rect 33778 32988 33784 33040
rect 33836 33028 33842 33040
rect 35621 33031 35679 33037
rect 35621 33028 35633 33031
rect 33836 33000 35633 33028
rect 33836 32988 33842 33000
rect 35621 32997 35633 33000
rect 35667 32997 35679 33031
rect 35621 32991 35679 32997
rect 37936 32960 37964 33056
rect 39850 32988 39856 33040
rect 39908 33028 39914 33040
rect 41414 33028 41420 33040
rect 39908 33000 41420 33028
rect 39908 32988 39914 33000
rect 41414 32988 41420 33000
rect 41472 32988 41478 33040
rect 42518 33028 42524 33040
rect 42479 33000 42524 33028
rect 42518 32988 42524 33000
rect 42576 32988 42582 33040
rect 40678 32960 40684 32972
rect 37476 32932 37964 32960
rect 40144 32932 40684 32960
rect 34790 32852 34796 32904
rect 34848 32892 34854 32904
rect 34974 32892 34980 32904
rect 34848 32864 34980 32892
rect 34848 32852 34854 32864
rect 34974 32852 34980 32864
rect 35032 32852 35038 32904
rect 35161 32895 35219 32901
rect 35161 32861 35173 32895
rect 35207 32892 35219 32895
rect 35710 32892 35716 32904
rect 35207 32864 35716 32892
rect 35207 32861 35219 32864
rect 35161 32855 35219 32861
rect 35710 32852 35716 32864
rect 35768 32852 35774 32904
rect 37476 32901 37504 32932
rect 37461 32895 37519 32901
rect 37461 32861 37473 32895
rect 37507 32861 37519 32895
rect 37642 32892 37648 32904
rect 37603 32864 37648 32892
rect 37461 32855 37519 32861
rect 37642 32852 37648 32864
rect 37700 32852 37706 32904
rect 38102 32892 38108 32904
rect 38063 32864 38108 32892
rect 38102 32852 38108 32864
rect 38160 32852 38166 32904
rect 38289 32895 38347 32901
rect 38289 32861 38301 32895
rect 38335 32892 38347 32895
rect 38378 32892 38384 32904
rect 38335 32864 38384 32892
rect 38335 32861 38347 32864
rect 38289 32855 38347 32861
rect 38378 32852 38384 32864
rect 38436 32852 38442 32904
rect 39942 32852 39948 32904
rect 40000 32892 40006 32904
rect 40144 32901 40172 32932
rect 40678 32920 40684 32932
rect 40736 32920 40742 32972
rect 40037 32895 40095 32901
rect 40037 32892 40049 32895
rect 40000 32864 40049 32892
rect 40000 32852 40006 32864
rect 40037 32861 40049 32864
rect 40083 32861 40095 32895
rect 40037 32855 40095 32861
rect 40129 32895 40187 32901
rect 40129 32861 40141 32895
rect 40175 32861 40187 32895
rect 40310 32892 40316 32904
rect 40271 32864 40316 32892
rect 40129 32855 40187 32861
rect 40310 32852 40316 32864
rect 40368 32852 40374 32904
rect 40402 32852 40408 32904
rect 40460 32892 40466 32904
rect 40460 32864 40505 32892
rect 40460 32852 40466 32864
rect 33468 32796 33532 32827
rect 33689 32827 33747 32833
rect 33468 32784 33474 32796
rect 33689 32793 33701 32827
rect 33735 32793 33747 32827
rect 33689 32787 33747 32793
rect 37734 32784 37740 32836
rect 37792 32824 37798 32836
rect 39853 32827 39911 32833
rect 39853 32824 39865 32827
rect 37792 32796 39865 32824
rect 37792 32784 37798 32796
rect 39853 32793 39865 32796
rect 39899 32793 39911 32827
rect 39853 32787 39911 32793
rect 33321 32759 33379 32765
rect 33321 32725 33333 32759
rect 33367 32725 33379 32759
rect 33321 32719 33379 32725
rect 34698 32716 34704 32768
rect 34756 32756 34762 32768
rect 35069 32759 35127 32765
rect 35069 32756 35081 32759
rect 34756 32728 35081 32756
rect 34756 32716 34762 32728
rect 35069 32725 35081 32728
rect 35115 32725 35127 32759
rect 35069 32719 35127 32725
rect 38654 32716 38660 32768
rect 38712 32756 38718 32768
rect 38749 32759 38807 32765
rect 38749 32756 38761 32759
rect 38712 32728 38761 32756
rect 38712 32716 38718 32728
rect 38749 32725 38761 32728
rect 38795 32725 38807 32759
rect 38749 32719 38807 32725
rect 39666 32716 39672 32768
rect 39724 32756 39730 32768
rect 41506 32756 41512 32768
rect 39724 32728 41512 32756
rect 39724 32716 39730 32728
rect 41506 32716 41512 32728
rect 41564 32716 41570 32768
rect 41966 32756 41972 32768
rect 41927 32728 41972 32756
rect 41966 32716 41972 32728
rect 42024 32756 42030 32768
rect 47854 32756 47860 32768
rect 42024 32728 47860 32756
rect 42024 32716 42030 32728
rect 47854 32716 47860 32728
rect 47912 32716 47918 32768
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 10413 32555 10471 32561
rect 10413 32521 10425 32555
rect 10459 32552 10471 32555
rect 10686 32552 10692 32564
rect 10459 32524 10692 32552
rect 10459 32521 10471 32524
rect 10413 32515 10471 32521
rect 10686 32512 10692 32524
rect 10744 32552 10750 32564
rect 14182 32552 14188 32564
rect 10744 32524 14188 32552
rect 10744 32512 10750 32524
rect 14182 32512 14188 32524
rect 14240 32552 14246 32564
rect 16666 32552 16672 32564
rect 14240 32524 14596 32552
rect 14240 32512 14246 32524
rect 13814 32484 13820 32496
rect 12912 32456 13820 32484
rect 1578 32376 1584 32428
rect 1636 32416 1642 32428
rect 1857 32419 1915 32425
rect 1857 32416 1869 32419
rect 1636 32388 1869 32416
rect 1636 32376 1642 32388
rect 1857 32385 1869 32388
rect 1903 32385 1915 32419
rect 12618 32416 12624 32428
rect 12579 32388 12624 32416
rect 1857 32379 1915 32385
rect 12618 32376 12624 32388
rect 12676 32376 12682 32428
rect 12710 32376 12716 32428
rect 12768 32416 12774 32428
rect 12912 32425 12940 32456
rect 13814 32444 13820 32456
rect 13872 32484 13878 32496
rect 14461 32487 14519 32493
rect 14461 32484 14473 32487
rect 13872 32456 14473 32484
rect 13872 32444 13878 32456
rect 14461 32453 14473 32456
rect 14507 32453 14519 32487
rect 14461 32447 14519 32453
rect 12897 32419 12955 32425
rect 12768 32388 12813 32416
rect 12768 32376 12774 32388
rect 12897 32385 12909 32419
rect 12943 32385 12955 32419
rect 12897 32379 12955 32385
rect 13170 32376 13176 32428
rect 13228 32416 13234 32428
rect 14568 32425 14596 32524
rect 14660 32524 15424 32552
rect 16627 32524 16672 32552
rect 13725 32419 13783 32425
rect 13725 32416 13737 32419
rect 13228 32388 13737 32416
rect 13228 32376 13234 32388
rect 13725 32385 13737 32388
rect 13771 32416 13783 32419
rect 14369 32419 14427 32425
rect 14369 32416 14381 32419
rect 13771 32388 14381 32416
rect 13771 32385 13783 32388
rect 13725 32379 13783 32385
rect 14369 32385 14381 32388
rect 14415 32385 14427 32419
rect 14369 32379 14427 32385
rect 14553 32419 14611 32425
rect 14553 32385 14565 32419
rect 14599 32385 14611 32419
rect 14553 32379 14611 32385
rect 12728 32348 12756 32376
rect 13262 32348 13268 32360
rect 12728 32320 13268 32348
rect 13262 32308 13268 32320
rect 13320 32308 13326 32360
rect 13909 32351 13967 32357
rect 13909 32317 13921 32351
rect 13955 32348 13967 32351
rect 14182 32348 14188 32360
rect 13955 32320 14188 32348
rect 13955 32317 13967 32320
rect 13909 32311 13967 32317
rect 14182 32308 14188 32320
rect 14240 32308 14246 32360
rect 14384 32348 14412 32379
rect 14660 32348 14688 32524
rect 15286 32484 15292 32496
rect 15247 32456 15292 32484
rect 15286 32444 15292 32456
rect 15344 32444 15350 32496
rect 15396 32484 15424 32524
rect 16666 32512 16672 32524
rect 16724 32512 16730 32564
rect 17402 32512 17408 32564
rect 17460 32552 17466 32564
rect 18249 32555 18307 32561
rect 18249 32552 18261 32555
rect 17460 32524 18261 32552
rect 17460 32512 17466 32524
rect 18249 32521 18261 32524
rect 18295 32521 18307 32555
rect 18249 32515 18307 32521
rect 18417 32555 18475 32561
rect 18417 32521 18429 32555
rect 18463 32552 18475 32555
rect 19426 32552 19432 32564
rect 18463 32524 19432 32552
rect 18463 32521 18475 32524
rect 18417 32515 18475 32521
rect 19426 32512 19432 32524
rect 19484 32512 19490 32564
rect 22557 32555 22615 32561
rect 22557 32521 22569 32555
rect 22603 32552 22615 32555
rect 22646 32552 22652 32564
rect 22603 32524 22652 32552
rect 22603 32521 22615 32524
rect 22557 32515 22615 32521
rect 22646 32512 22652 32524
rect 22704 32512 22710 32564
rect 24581 32555 24639 32561
rect 24581 32521 24593 32555
rect 24627 32521 24639 32555
rect 25958 32552 25964 32564
rect 25919 32524 25964 32552
rect 24581 32515 24639 32521
rect 15396 32456 17448 32484
rect 16850 32416 16856 32428
rect 15962 32388 16856 32416
rect 16850 32376 16856 32388
rect 16908 32416 16914 32428
rect 17310 32416 17316 32428
rect 16908 32388 17316 32416
rect 16908 32376 16914 32388
rect 17310 32376 17316 32388
rect 17368 32376 17374 32428
rect 17420 32416 17448 32456
rect 17862 32444 17868 32496
rect 17920 32484 17926 32496
rect 18049 32487 18107 32493
rect 18049 32484 18061 32487
rect 17920 32456 18061 32484
rect 17920 32444 17926 32456
rect 18049 32453 18061 32456
rect 18095 32453 18107 32487
rect 21818 32484 21824 32496
rect 18049 32447 18107 32453
rect 18156 32456 21824 32484
rect 18156 32416 18184 32456
rect 21818 32444 21824 32456
rect 21876 32444 21882 32496
rect 22002 32444 22008 32496
rect 22060 32484 22066 32496
rect 23201 32487 23259 32493
rect 22060 32456 22600 32484
rect 22060 32444 22066 32456
rect 17420 32388 18184 32416
rect 18322 32376 18328 32428
rect 18380 32416 18386 32428
rect 19061 32419 19119 32425
rect 19061 32416 19073 32419
rect 18380 32388 19073 32416
rect 18380 32376 18386 32388
rect 19061 32385 19073 32388
rect 19107 32385 19119 32419
rect 19061 32379 19119 32385
rect 19245 32419 19303 32425
rect 19245 32385 19257 32419
rect 19291 32385 19303 32419
rect 19245 32379 19303 32385
rect 14384 32320 14688 32348
rect 14734 32308 14740 32360
rect 14792 32348 14798 32360
rect 15841 32351 15899 32357
rect 15841 32348 15853 32351
rect 14792 32320 15853 32348
rect 14792 32308 14798 32320
rect 15841 32317 15853 32320
rect 15887 32348 15899 32351
rect 17037 32351 17095 32357
rect 17037 32348 17049 32351
rect 15887 32320 17049 32348
rect 15887 32317 15899 32320
rect 15841 32311 15899 32317
rect 17037 32317 17049 32320
rect 17083 32348 17095 32351
rect 17494 32348 17500 32360
rect 17083 32320 17500 32348
rect 17083 32317 17095 32320
rect 17037 32311 17095 32317
rect 17494 32308 17500 32320
rect 17552 32308 17558 32360
rect 18230 32308 18236 32360
rect 18288 32348 18294 32360
rect 19260 32348 19288 32379
rect 19334 32376 19340 32428
rect 19392 32416 19398 32428
rect 19889 32419 19947 32425
rect 19889 32416 19901 32419
rect 19392 32388 19901 32416
rect 19392 32376 19398 32388
rect 19889 32385 19901 32388
rect 19935 32385 19947 32419
rect 19889 32379 19947 32385
rect 19978 32376 19984 32428
rect 20036 32416 20042 32428
rect 20073 32419 20131 32425
rect 20073 32416 20085 32419
rect 20036 32388 20085 32416
rect 20036 32376 20042 32388
rect 20073 32385 20085 32388
rect 20119 32385 20131 32419
rect 20073 32379 20131 32385
rect 20990 32376 20996 32428
rect 21048 32416 21054 32428
rect 21085 32419 21143 32425
rect 21085 32416 21097 32419
rect 21048 32388 21097 32416
rect 21048 32376 21054 32388
rect 21085 32385 21097 32388
rect 21131 32385 21143 32419
rect 21085 32379 21143 32385
rect 21269 32419 21327 32425
rect 21269 32385 21281 32419
rect 21315 32416 21327 32419
rect 21450 32416 21456 32428
rect 21315 32388 21456 32416
rect 21315 32385 21327 32388
rect 21269 32379 21327 32385
rect 21450 32376 21456 32388
rect 21508 32376 21514 32428
rect 21913 32419 21971 32425
rect 21913 32385 21925 32419
rect 21959 32416 21971 32419
rect 22094 32416 22100 32428
rect 21959 32388 22100 32416
rect 21959 32385 21971 32388
rect 21913 32379 21971 32385
rect 22094 32376 22100 32388
rect 22152 32416 22158 32428
rect 22278 32416 22284 32428
rect 22152 32388 22284 32416
rect 22152 32376 22158 32388
rect 22278 32376 22284 32388
rect 22336 32416 22342 32428
rect 22572 32425 22600 32456
rect 23201 32453 23213 32487
rect 23247 32484 23259 32487
rect 23566 32484 23572 32496
rect 23247 32456 23572 32484
rect 23247 32453 23259 32456
rect 23201 32447 23259 32453
rect 23566 32444 23572 32456
rect 23624 32484 23630 32496
rect 24596 32484 24624 32515
rect 25958 32512 25964 32524
rect 26016 32512 26022 32564
rect 27798 32512 27804 32564
rect 27856 32552 27862 32564
rect 27856 32524 28488 32552
rect 27856 32512 27862 32524
rect 23624 32456 24624 32484
rect 24673 32487 24731 32493
rect 23624 32444 23630 32456
rect 24673 32453 24685 32487
rect 24719 32484 24731 32487
rect 24946 32484 24952 32496
rect 24719 32456 24952 32484
rect 24719 32453 24731 32456
rect 24673 32447 24731 32453
rect 24946 32444 24952 32456
rect 25004 32484 25010 32496
rect 27522 32484 27528 32496
rect 25004 32456 26004 32484
rect 25004 32444 25010 32456
rect 22373 32419 22431 32425
rect 22373 32416 22385 32419
rect 22336 32388 22385 32416
rect 22336 32376 22342 32388
rect 22373 32385 22385 32388
rect 22419 32385 22431 32419
rect 22373 32379 22431 32385
rect 22557 32419 22615 32425
rect 22557 32385 22569 32419
rect 22603 32385 22615 32419
rect 23382 32416 23388 32428
rect 23343 32388 23388 32416
rect 22557 32379 22615 32385
rect 23382 32376 23388 32388
rect 23440 32376 23446 32428
rect 23477 32419 23535 32425
rect 23477 32385 23489 32419
rect 23523 32385 23535 32419
rect 23477 32379 23535 32385
rect 24581 32419 24639 32425
rect 24581 32385 24593 32419
rect 24627 32416 24639 32419
rect 24857 32419 24915 32425
rect 24627 32388 24808 32416
rect 24627 32385 24639 32388
rect 24581 32379 24639 32385
rect 18288 32320 19288 32348
rect 18288 32308 18294 32320
rect 22462 32308 22468 32360
rect 22520 32348 22526 32360
rect 23290 32348 23296 32360
rect 22520 32320 23296 32348
rect 22520 32308 22526 32320
rect 23290 32308 23296 32320
rect 23348 32348 23354 32360
rect 23492 32348 23520 32379
rect 23348 32320 23520 32348
rect 23348 32308 23354 32320
rect 12802 32280 12808 32292
rect 12763 32252 12808 32280
rect 12802 32240 12808 32252
rect 12860 32240 12866 32292
rect 13081 32283 13139 32289
rect 13081 32249 13093 32283
rect 13127 32280 13139 32283
rect 16666 32280 16672 32292
rect 13127 32252 16672 32280
rect 13127 32249 13139 32252
rect 13081 32243 13139 32249
rect 16666 32240 16672 32252
rect 16724 32240 16730 32292
rect 17954 32240 17960 32292
rect 18012 32280 18018 32292
rect 18877 32283 18935 32289
rect 18877 32280 18889 32283
rect 18012 32252 18889 32280
rect 18012 32240 18018 32252
rect 18877 32249 18889 32252
rect 18923 32249 18935 32283
rect 18877 32243 18935 32249
rect 20438 32240 20444 32292
rect 20496 32280 20502 32292
rect 20496 32252 21128 32280
rect 20496 32240 20502 32252
rect 1946 32212 1952 32224
rect 1907 32184 1952 32212
rect 1946 32172 1952 32184
rect 2004 32172 2010 32224
rect 8938 32172 8944 32224
rect 8996 32212 9002 32224
rect 10873 32215 10931 32221
rect 10873 32212 10885 32215
rect 8996 32184 10885 32212
rect 8996 32172 9002 32184
rect 10873 32181 10885 32184
rect 10919 32212 10931 32215
rect 11974 32212 11980 32224
rect 10919 32184 11980 32212
rect 10919 32181 10931 32184
rect 10873 32175 10931 32181
rect 11974 32172 11980 32184
rect 12032 32172 12038 32224
rect 13538 32212 13544 32224
rect 13499 32184 13544 32212
rect 13538 32172 13544 32184
rect 13596 32172 13602 32224
rect 14826 32172 14832 32224
rect 14884 32212 14890 32224
rect 15194 32212 15200 32224
rect 14884 32184 15200 32212
rect 14884 32172 14890 32184
rect 15194 32172 15200 32184
rect 15252 32172 15258 32224
rect 17034 32172 17040 32224
rect 17092 32212 17098 32224
rect 17497 32215 17555 32221
rect 17497 32212 17509 32215
rect 17092 32184 17509 32212
rect 17092 32172 17098 32184
rect 17497 32181 17509 32184
rect 17543 32181 17555 32215
rect 17497 32175 17555 32181
rect 17586 32172 17592 32224
rect 17644 32212 17650 32224
rect 18233 32215 18291 32221
rect 18233 32212 18245 32215
rect 17644 32184 18245 32212
rect 17644 32172 17650 32184
rect 18233 32181 18245 32184
rect 18279 32181 18291 32215
rect 18233 32175 18291 32181
rect 19981 32215 20039 32221
rect 19981 32181 19993 32215
rect 20027 32212 20039 32215
rect 20714 32212 20720 32224
rect 20027 32184 20720 32212
rect 20027 32181 20039 32184
rect 19981 32175 20039 32181
rect 20714 32172 20720 32184
rect 20772 32172 20778 32224
rect 20806 32172 20812 32224
rect 20864 32212 20870 32224
rect 21100 32221 21128 32252
rect 22278 32240 22284 32292
rect 22336 32280 22342 32292
rect 23474 32280 23480 32292
rect 22336 32252 23480 32280
rect 22336 32240 22342 32252
rect 23474 32240 23480 32252
rect 23532 32240 23538 32292
rect 23661 32283 23719 32289
rect 23661 32249 23673 32283
rect 23707 32280 23719 32283
rect 24670 32280 24676 32292
rect 23707 32252 24676 32280
rect 23707 32249 23719 32252
rect 23661 32243 23719 32249
rect 24670 32240 24676 32252
rect 24728 32240 24734 32292
rect 24780 32280 24808 32388
rect 24857 32385 24869 32419
rect 24903 32385 24915 32419
rect 25498 32416 25504 32428
rect 25459 32388 25504 32416
rect 24857 32379 24915 32385
rect 24872 32348 24900 32379
rect 25498 32376 25504 32388
rect 25556 32376 25562 32428
rect 25976 32425 26004 32456
rect 26988 32456 27528 32484
rect 25961 32419 26019 32425
rect 25961 32385 25973 32419
rect 26007 32385 26019 32419
rect 25961 32379 26019 32385
rect 26145 32419 26203 32425
rect 26145 32385 26157 32419
rect 26191 32385 26203 32419
rect 26145 32379 26203 32385
rect 25409 32351 25467 32357
rect 25409 32348 25421 32351
rect 24872 32320 25421 32348
rect 25409 32317 25421 32320
rect 25455 32348 25467 32351
rect 26160 32348 26188 32379
rect 26786 32376 26792 32428
rect 26844 32416 26850 32428
rect 26988 32425 27016 32456
rect 27522 32444 27528 32456
rect 27580 32444 27586 32496
rect 27982 32444 27988 32496
rect 28040 32444 28046 32496
rect 28460 32484 28488 32524
rect 28534 32512 28540 32564
rect 28592 32552 28598 32564
rect 28905 32555 28963 32561
rect 28905 32552 28917 32555
rect 28592 32524 28917 32552
rect 28592 32512 28598 32524
rect 28905 32521 28917 32524
rect 28951 32521 28963 32555
rect 29546 32552 29552 32564
rect 29507 32524 29552 32552
rect 28905 32515 28963 32521
rect 29546 32512 29552 32524
rect 29604 32512 29610 32564
rect 31478 32552 31484 32564
rect 31439 32524 31484 32552
rect 31478 32512 31484 32524
rect 31536 32512 31542 32564
rect 32493 32555 32551 32561
rect 32493 32521 32505 32555
rect 32539 32552 32551 32555
rect 32766 32552 32772 32564
rect 32539 32524 32772 32552
rect 32539 32521 32551 32524
rect 32493 32515 32551 32521
rect 32766 32512 32772 32524
rect 32824 32512 32830 32564
rect 32950 32512 32956 32564
rect 33008 32552 33014 32564
rect 33597 32555 33655 32561
rect 33597 32552 33609 32555
rect 33008 32524 33609 32552
rect 33008 32512 33014 32524
rect 33597 32521 33609 32524
rect 33643 32521 33655 32555
rect 33962 32552 33968 32564
rect 33923 32524 33968 32552
rect 33597 32515 33655 32521
rect 33962 32512 33968 32524
rect 34020 32512 34026 32564
rect 34977 32555 35035 32561
rect 34977 32521 34989 32555
rect 35023 32552 35035 32555
rect 35342 32552 35348 32564
rect 35023 32524 35348 32552
rect 35023 32521 35035 32524
rect 34977 32515 35035 32521
rect 35342 32512 35348 32524
rect 35400 32512 35406 32564
rect 35894 32512 35900 32564
rect 35952 32552 35958 32564
rect 36449 32555 36507 32561
rect 36449 32552 36461 32555
rect 35952 32524 36461 32552
rect 35952 32512 35958 32524
rect 36449 32521 36461 32524
rect 36495 32521 36507 32555
rect 36449 32515 36507 32521
rect 37642 32512 37648 32564
rect 37700 32552 37706 32564
rect 38105 32555 38163 32561
rect 38105 32552 38117 32555
rect 37700 32524 38117 32552
rect 37700 32512 37706 32524
rect 38105 32521 38117 32524
rect 38151 32521 38163 32555
rect 38105 32515 38163 32521
rect 39850 32512 39856 32564
rect 39908 32552 39914 32564
rect 40037 32555 40095 32561
rect 40037 32552 40049 32555
rect 39908 32524 40049 32552
rect 39908 32512 39914 32524
rect 40037 32521 40049 32524
rect 40083 32521 40095 32555
rect 40037 32515 40095 32521
rect 29825 32487 29883 32493
rect 29825 32484 29837 32487
rect 28460 32456 29837 32484
rect 29825 32453 29837 32456
rect 29871 32453 29883 32487
rect 30742 32484 30748 32496
rect 29825 32447 29883 32453
rect 30116 32456 30748 32484
rect 26973 32419 27031 32425
rect 26973 32416 26985 32419
rect 26844 32388 26985 32416
rect 26844 32376 26850 32388
rect 26973 32385 26985 32388
rect 27019 32385 27031 32419
rect 27154 32416 27160 32428
rect 27115 32388 27160 32416
rect 26973 32379 27031 32385
rect 27154 32376 27160 32388
rect 27212 32376 27218 32428
rect 27614 32376 27620 32428
rect 27672 32416 27678 32428
rect 27893 32419 27951 32425
rect 27893 32416 27905 32419
rect 27672 32388 27905 32416
rect 27672 32376 27678 32388
rect 27893 32385 27905 32388
rect 27939 32385 27951 32419
rect 28000 32416 28028 32444
rect 28077 32419 28135 32425
rect 28077 32416 28089 32419
rect 28000 32388 28089 32416
rect 27893 32379 27951 32385
rect 28077 32385 28089 32388
rect 28123 32385 28135 32419
rect 28077 32379 28135 32385
rect 28629 32419 28687 32425
rect 28629 32385 28641 32419
rect 28675 32385 28687 32419
rect 28810 32416 28816 32428
rect 28771 32388 28816 32416
rect 28629 32379 28687 32385
rect 27798 32348 27804 32360
rect 25455 32320 26188 32348
rect 27759 32320 27804 32348
rect 25455 32317 25467 32320
rect 25409 32311 25467 32317
rect 27798 32308 27804 32320
rect 27856 32308 27862 32360
rect 27985 32351 28043 32357
rect 27985 32317 27997 32351
rect 28031 32348 28043 32351
rect 28258 32348 28264 32360
rect 28031 32320 28264 32348
rect 28031 32317 28043 32320
rect 27985 32311 28043 32317
rect 28258 32308 28264 32320
rect 28316 32308 28322 32360
rect 28644 32348 28672 32379
rect 28810 32376 28816 32388
rect 28868 32376 28874 32428
rect 29730 32416 29736 32428
rect 29691 32388 29736 32416
rect 29730 32376 29736 32388
rect 29788 32376 29794 32428
rect 29914 32416 29920 32428
rect 29875 32388 29920 32416
rect 29914 32376 29920 32388
rect 29972 32376 29978 32428
rect 30116 32425 30144 32456
rect 30742 32444 30748 32456
rect 30800 32444 30806 32496
rect 30834 32444 30840 32496
rect 30892 32484 30898 32496
rect 30929 32487 30987 32493
rect 30929 32484 30941 32487
rect 30892 32456 30941 32484
rect 30892 32444 30898 32456
rect 30929 32453 30941 32456
rect 30975 32484 30987 32487
rect 31570 32484 31576 32496
rect 30975 32456 31576 32484
rect 30975 32453 30987 32456
rect 30929 32447 30987 32453
rect 31570 32444 31576 32456
rect 31628 32444 31634 32496
rect 32122 32444 32128 32496
rect 32180 32484 32186 32496
rect 32652 32487 32710 32493
rect 32652 32484 32664 32487
rect 32180 32456 32664 32484
rect 32180 32444 32186 32456
rect 32652 32453 32664 32456
rect 32698 32484 32710 32487
rect 33410 32484 33416 32496
rect 32698 32456 33416 32484
rect 32698 32453 32710 32456
rect 32652 32447 32710 32453
rect 33410 32444 33416 32456
rect 33468 32444 33474 32496
rect 33612 32456 34100 32484
rect 30101 32419 30159 32425
rect 30101 32385 30113 32419
rect 30147 32385 30159 32419
rect 30101 32379 30159 32385
rect 30193 32419 30251 32425
rect 30193 32385 30205 32419
rect 30239 32385 30251 32419
rect 30650 32416 30656 32428
rect 30611 32388 30656 32416
rect 30193 32379 30251 32385
rect 29362 32348 29368 32360
rect 28644 32320 29368 32348
rect 29362 32308 29368 32320
rect 29420 32308 29426 32360
rect 29638 32308 29644 32360
rect 29696 32348 29702 32360
rect 30208 32348 30236 32379
rect 30650 32376 30656 32388
rect 30708 32376 30714 32428
rect 32769 32419 32827 32425
rect 32769 32385 32781 32419
rect 32815 32416 32827 32419
rect 33612 32416 33640 32456
rect 34072 32428 34100 32456
rect 34698 32444 34704 32496
rect 34756 32484 34762 32496
rect 34756 32456 36400 32484
rect 34756 32444 34762 32456
rect 33778 32416 33784 32428
rect 32815 32388 33640 32416
rect 33739 32388 33784 32416
rect 32815 32385 32827 32388
rect 32769 32379 32827 32385
rect 33778 32376 33784 32388
rect 33836 32376 33842 32428
rect 34054 32416 34060 32428
rect 34015 32388 34060 32416
rect 34054 32376 34060 32388
rect 34112 32376 34118 32428
rect 34790 32416 34796 32428
rect 34751 32388 34796 32416
rect 34790 32376 34796 32388
rect 34848 32376 34854 32428
rect 35069 32419 35127 32425
rect 35069 32385 35081 32419
rect 35115 32416 35127 32419
rect 35434 32416 35440 32428
rect 35115 32388 35440 32416
rect 35115 32385 35127 32388
rect 35069 32379 35127 32385
rect 35434 32376 35440 32388
rect 35492 32376 35498 32428
rect 35710 32416 35716 32428
rect 35671 32388 35716 32416
rect 35710 32376 35716 32388
rect 35768 32376 35774 32428
rect 36372 32425 36400 32456
rect 38654 32444 38660 32496
rect 38712 32484 38718 32496
rect 39485 32487 39543 32493
rect 39485 32484 39497 32487
rect 38712 32456 39497 32484
rect 38712 32444 38718 32456
rect 39485 32453 39497 32456
rect 39531 32484 39543 32487
rect 39666 32484 39672 32496
rect 39531 32456 39672 32484
rect 39531 32453 39543 32456
rect 39485 32447 39543 32453
rect 39666 32444 39672 32456
rect 39724 32444 39730 32496
rect 36357 32419 36415 32425
rect 36357 32385 36369 32419
rect 36403 32385 36415 32419
rect 36357 32379 36415 32385
rect 36541 32419 36599 32425
rect 36541 32385 36553 32419
rect 36587 32385 36599 32419
rect 37458 32416 37464 32428
rect 37419 32388 37464 32416
rect 36541 32379 36599 32385
rect 29696 32320 30236 32348
rect 29696 32308 29702 32320
rect 32398 32308 32404 32360
rect 32456 32348 32462 32360
rect 32674 32348 32680 32360
rect 32456 32320 32680 32348
rect 32456 32308 32462 32320
rect 32674 32308 32680 32320
rect 32732 32348 32738 32360
rect 32861 32351 32919 32357
rect 32861 32348 32873 32351
rect 32732 32320 32873 32348
rect 32732 32308 32738 32320
rect 32861 32317 32873 32320
rect 32907 32317 32919 32351
rect 32861 32311 32919 32317
rect 33137 32351 33195 32357
rect 33137 32317 33149 32351
rect 33183 32348 33195 32351
rect 33318 32348 33324 32360
rect 33183 32320 33324 32348
rect 33183 32317 33195 32320
rect 33137 32311 33195 32317
rect 33318 32308 33324 32320
rect 33376 32308 33382 32360
rect 33796 32348 33824 32376
rect 34609 32351 34667 32357
rect 34609 32348 34621 32351
rect 33796 32320 34621 32348
rect 34609 32317 34621 32320
rect 34655 32317 34667 32351
rect 34609 32311 34667 32317
rect 34974 32308 34980 32360
rect 35032 32348 35038 32360
rect 35894 32348 35900 32360
rect 35032 32320 35900 32348
rect 35032 32308 35038 32320
rect 35894 32308 35900 32320
rect 35952 32308 35958 32360
rect 25222 32280 25228 32292
rect 24780 32252 25228 32280
rect 25222 32240 25228 32252
rect 25280 32280 25286 32292
rect 25590 32280 25596 32292
rect 25280 32252 25596 32280
rect 25280 32240 25286 32252
rect 25590 32240 25596 32252
rect 25648 32240 25654 32292
rect 27065 32283 27123 32289
rect 27065 32249 27077 32283
rect 27111 32280 27123 32283
rect 28350 32280 28356 32292
rect 27111 32252 28356 32280
rect 27111 32249 27123 32252
rect 27065 32243 27123 32249
rect 28350 32240 28356 32252
rect 28408 32240 28414 32292
rect 28626 32240 28632 32292
rect 28684 32280 28690 32292
rect 30926 32280 30932 32292
rect 28684 32252 30788 32280
rect 30887 32252 30932 32280
rect 28684 32240 28690 32252
rect 20901 32215 20959 32221
rect 20901 32212 20913 32215
rect 20864 32184 20913 32212
rect 20864 32172 20870 32184
rect 20901 32181 20913 32184
rect 20947 32181 20959 32215
rect 20901 32175 20959 32181
rect 21085 32215 21143 32221
rect 21085 32181 21097 32215
rect 21131 32181 21143 32215
rect 21085 32175 21143 32181
rect 22186 32172 22192 32224
rect 22244 32212 22250 32224
rect 23201 32215 23259 32221
rect 23201 32212 23213 32215
rect 22244 32184 23213 32212
rect 22244 32172 22250 32184
rect 23201 32181 23213 32184
rect 23247 32181 23259 32215
rect 23201 32175 23259 32181
rect 27617 32215 27675 32221
rect 27617 32181 27629 32215
rect 27663 32212 27675 32215
rect 27890 32212 27896 32224
rect 27663 32184 27896 32212
rect 27663 32181 27675 32184
rect 27617 32175 27675 32181
rect 27890 32172 27896 32184
rect 27948 32172 27954 32224
rect 28994 32172 29000 32224
rect 29052 32212 29058 32224
rect 29089 32215 29147 32221
rect 29089 32212 29101 32215
rect 29052 32184 29101 32212
rect 29052 32172 29058 32184
rect 29089 32181 29101 32184
rect 29135 32181 29147 32215
rect 29089 32175 29147 32181
rect 29730 32172 29736 32224
rect 29788 32212 29794 32224
rect 30006 32212 30012 32224
rect 29788 32184 30012 32212
rect 29788 32172 29794 32184
rect 30006 32172 30012 32184
rect 30064 32172 30070 32224
rect 30760 32212 30788 32252
rect 30926 32240 30932 32252
rect 30984 32240 30990 32292
rect 35802 32280 35808 32292
rect 35544 32252 35808 32280
rect 30834 32212 30840 32224
rect 30760 32184 30840 32212
rect 30834 32172 30840 32184
rect 30892 32172 30898 32224
rect 33962 32172 33968 32224
rect 34020 32212 34026 32224
rect 34514 32212 34520 32224
rect 34020 32184 34520 32212
rect 34020 32172 34026 32184
rect 34514 32172 34520 32184
rect 34572 32212 34578 32224
rect 35544 32221 35572 32252
rect 35802 32240 35808 32252
rect 35860 32280 35866 32292
rect 36556 32280 36584 32379
rect 37458 32376 37464 32388
rect 37516 32376 37522 32428
rect 37645 32419 37703 32425
rect 37645 32385 37657 32419
rect 37691 32416 37703 32419
rect 37734 32416 37740 32428
rect 37691 32388 37740 32416
rect 37691 32385 37703 32388
rect 37645 32379 37703 32385
rect 37734 32376 37740 32388
rect 37792 32376 37798 32428
rect 38102 32376 38108 32428
rect 38160 32416 38166 32428
rect 38289 32419 38347 32425
rect 38289 32416 38301 32419
rect 38160 32388 38301 32416
rect 38160 32376 38166 32388
rect 38289 32385 38301 32388
rect 38335 32416 38347 32419
rect 38746 32416 38752 32428
rect 38335 32388 38752 32416
rect 38335 32385 38347 32388
rect 38289 32379 38347 32385
rect 38746 32376 38752 32388
rect 38804 32416 38810 32428
rect 40589 32419 40647 32425
rect 40589 32416 40601 32419
rect 38804 32388 40601 32416
rect 38804 32376 38810 32388
rect 40589 32385 40601 32388
rect 40635 32385 40647 32419
rect 40589 32379 40647 32385
rect 43254 32376 43260 32428
rect 43312 32416 43318 32428
rect 47670 32416 47676 32428
rect 43312 32388 47676 32416
rect 43312 32376 43318 32388
rect 47670 32376 47676 32388
rect 47728 32416 47734 32428
rect 47857 32419 47915 32425
rect 47857 32416 47869 32419
rect 47728 32388 47869 32416
rect 47728 32376 47734 32388
rect 47857 32385 47869 32388
rect 47903 32385 47915 32419
rect 47857 32379 47915 32385
rect 38378 32308 38384 32360
rect 38436 32348 38442 32360
rect 38473 32351 38531 32357
rect 38473 32348 38485 32351
rect 38436 32320 38485 32348
rect 38436 32308 38442 32320
rect 38473 32317 38485 32320
rect 38519 32317 38531 32351
rect 38473 32311 38531 32317
rect 39574 32308 39580 32360
rect 39632 32348 39638 32360
rect 40954 32348 40960 32360
rect 39632 32320 40960 32348
rect 39632 32308 39638 32320
rect 40954 32308 40960 32320
rect 41012 32348 41018 32360
rect 41693 32351 41751 32357
rect 41693 32348 41705 32351
rect 41012 32320 41705 32348
rect 41012 32308 41018 32320
rect 41693 32317 41705 32320
rect 41739 32317 41751 32351
rect 41693 32311 41751 32317
rect 35860 32252 36584 32280
rect 35860 32240 35866 32252
rect 38562 32240 38568 32292
rect 38620 32280 38626 32292
rect 38933 32283 38991 32289
rect 38933 32280 38945 32283
rect 38620 32252 38945 32280
rect 38620 32240 38626 32252
rect 38933 32249 38945 32252
rect 38979 32249 38991 32283
rect 38933 32243 38991 32249
rect 35529 32215 35587 32221
rect 35529 32212 35541 32215
rect 34572 32184 35541 32212
rect 34572 32172 34578 32184
rect 35529 32181 35541 32184
rect 35575 32181 35587 32215
rect 35529 32175 35587 32181
rect 36538 32172 36544 32224
rect 36596 32212 36602 32224
rect 37277 32215 37335 32221
rect 37277 32212 37289 32215
rect 36596 32184 37289 32212
rect 36596 32172 36602 32184
rect 37277 32181 37289 32184
rect 37323 32181 37335 32215
rect 37277 32175 37335 32181
rect 40402 32172 40408 32224
rect 40460 32212 40466 32224
rect 41141 32215 41199 32221
rect 41141 32212 41153 32215
rect 40460 32184 41153 32212
rect 40460 32172 40466 32184
rect 41141 32181 41153 32184
rect 41187 32212 41199 32215
rect 41966 32212 41972 32224
rect 41187 32184 41972 32212
rect 41187 32181 41199 32184
rect 41141 32175 41199 32181
rect 41966 32172 41972 32184
rect 42024 32172 42030 32224
rect 48038 32212 48044 32224
rect 47999 32184 48044 32212
rect 48038 32172 48044 32184
rect 48096 32172 48102 32224
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 1578 32008 1584 32020
rect 1539 31980 1584 32008
rect 1578 31968 1584 31980
rect 1636 31968 1642 32020
rect 10686 32008 10692 32020
rect 10647 31980 10692 32008
rect 10686 31968 10692 31980
rect 10744 31968 10750 32020
rect 11333 32011 11391 32017
rect 11333 31977 11345 32011
rect 11379 32008 11391 32011
rect 11790 32008 11796 32020
rect 11379 31980 11796 32008
rect 11379 31977 11391 31980
rect 11333 31971 11391 31977
rect 11790 31968 11796 31980
rect 11848 31968 11854 32020
rect 12621 32011 12679 32017
rect 12621 31977 12633 32011
rect 12667 32008 12679 32011
rect 12802 32008 12808 32020
rect 12667 31980 12808 32008
rect 12667 31977 12679 31980
rect 12621 31971 12679 31977
rect 12802 31968 12808 31980
rect 12860 31968 12866 32020
rect 14277 32011 14335 32017
rect 14277 31977 14289 32011
rect 14323 32008 14335 32011
rect 15013 32011 15071 32017
rect 15013 32008 15025 32011
rect 14323 31980 15025 32008
rect 14323 31977 14335 31980
rect 14277 31971 14335 31977
rect 15013 31977 15025 31980
rect 15059 32008 15071 32011
rect 15059 31980 15608 32008
rect 15059 31977 15071 31980
rect 15013 31971 15071 31977
rect 1946 31900 1952 31952
rect 2004 31940 2010 31952
rect 15194 31940 15200 31952
rect 2004 31912 15200 31940
rect 2004 31900 2010 31912
rect 15194 31900 15200 31912
rect 15252 31900 15258 31952
rect 13722 31832 13728 31884
rect 13780 31872 13786 31884
rect 15580 31872 15608 31980
rect 15654 31968 15660 32020
rect 15712 32008 15718 32020
rect 15933 32011 15991 32017
rect 15933 32008 15945 32011
rect 15712 31980 15945 32008
rect 15712 31968 15718 31980
rect 15933 31977 15945 31980
rect 15979 31977 15991 32011
rect 16574 32008 16580 32020
rect 16535 31980 16580 32008
rect 15933 31971 15991 31977
rect 16574 31968 16580 31980
rect 16632 31968 16638 32020
rect 19245 32011 19303 32017
rect 19245 31977 19257 32011
rect 19291 32008 19303 32011
rect 19334 32008 19340 32020
rect 19291 31980 19340 32008
rect 19291 31977 19303 31980
rect 19245 31971 19303 31977
rect 19334 31968 19340 31980
rect 19392 31968 19398 32020
rect 20441 32011 20499 32017
rect 20441 31977 20453 32011
rect 20487 32008 20499 32011
rect 22833 32011 22891 32017
rect 20487 31980 22784 32008
rect 20487 31977 20499 31980
rect 20441 31971 20499 31977
rect 17129 31943 17187 31949
rect 17129 31909 17141 31943
rect 17175 31909 17187 31943
rect 17129 31903 17187 31909
rect 17144 31872 17172 31903
rect 18874 31900 18880 31952
rect 18932 31940 18938 31952
rect 20806 31940 20812 31952
rect 18932 31912 19564 31940
rect 20767 31912 20812 31940
rect 18932 31900 18938 31912
rect 13780 31844 14412 31872
rect 15580 31844 15792 31872
rect 17144 31844 19288 31872
rect 13780 31832 13786 31844
rect 10229 31807 10287 31813
rect 10229 31773 10241 31807
rect 10275 31804 10287 31807
rect 12342 31804 12348 31816
rect 10275 31776 12348 31804
rect 10275 31773 10287 31776
rect 10229 31767 10287 31773
rect 12342 31764 12348 31776
rect 12400 31764 12406 31816
rect 12437 31807 12495 31813
rect 12437 31773 12449 31807
rect 12483 31804 12495 31807
rect 12526 31804 12532 31816
rect 12483 31776 12532 31804
rect 12483 31773 12495 31776
rect 12437 31767 12495 31773
rect 12526 31764 12532 31776
rect 12584 31764 12590 31816
rect 12621 31807 12679 31813
rect 12621 31773 12633 31807
rect 12667 31804 12679 31807
rect 13357 31807 13415 31813
rect 13357 31804 13369 31807
rect 12667 31776 13369 31804
rect 12667 31773 12679 31776
rect 12621 31767 12679 31773
rect 13357 31773 13369 31776
rect 13403 31804 13415 31807
rect 13538 31804 13544 31816
rect 13403 31776 13544 31804
rect 13403 31773 13415 31776
rect 13357 31767 13415 31773
rect 13538 31764 13544 31776
rect 13596 31764 13602 31816
rect 13630 31764 13636 31816
rect 13688 31764 13694 31816
rect 13814 31764 13820 31816
rect 13872 31804 13878 31816
rect 14093 31807 14151 31813
rect 14093 31804 14105 31807
rect 13872 31776 14105 31804
rect 13872 31764 13878 31776
rect 14093 31773 14105 31776
rect 14139 31773 14151 31807
rect 14093 31767 14151 31773
rect 14182 31764 14188 31816
rect 14240 31804 14246 31816
rect 14384 31813 14412 31844
rect 14369 31807 14427 31813
rect 14240 31776 14285 31804
rect 14240 31764 14246 31776
rect 14369 31773 14381 31807
rect 14415 31773 14427 31807
rect 14369 31767 14427 31773
rect 14826 31764 14832 31816
rect 14884 31764 14890 31816
rect 15764 31813 15792 31844
rect 15657 31807 15715 31813
rect 15657 31804 15669 31807
rect 15028 31776 15669 31804
rect 13173 31739 13231 31745
rect 13173 31705 13185 31739
rect 13219 31736 13231 31739
rect 13648 31736 13676 31764
rect 13219 31708 13676 31736
rect 13219 31705 13231 31708
rect 13173 31699 13231 31705
rect 13541 31671 13599 31677
rect 13541 31637 13553 31671
rect 13587 31668 13599 31671
rect 13722 31668 13728 31680
rect 13587 31640 13728 31668
rect 13587 31637 13599 31640
rect 13541 31631 13599 31637
rect 13722 31628 13728 31640
rect 13780 31628 13786 31680
rect 14844 31677 14872 31764
rect 15028 31748 15056 31776
rect 15657 31773 15669 31776
rect 15703 31773 15715 31807
rect 15657 31767 15715 31773
rect 15749 31807 15807 31813
rect 15749 31773 15761 31807
rect 15795 31773 15807 31807
rect 17126 31804 17132 31816
rect 17087 31776 17132 31804
rect 15749 31767 15807 31773
rect 17126 31764 17132 31776
rect 17184 31764 17190 31816
rect 17402 31804 17408 31816
rect 17363 31776 17408 31804
rect 17402 31764 17408 31776
rect 17460 31804 17466 31816
rect 17862 31804 17868 31816
rect 17460 31776 17868 31804
rect 17460 31764 17466 31776
rect 17862 31764 17868 31776
rect 17920 31764 17926 31816
rect 18233 31807 18291 31813
rect 18233 31804 18245 31807
rect 17972 31776 18245 31804
rect 15010 31745 15016 31748
rect 14997 31739 15016 31745
rect 14997 31705 15009 31739
rect 15068 31736 15074 31748
rect 15197 31739 15255 31745
rect 15068 31708 15145 31736
rect 14997 31699 15016 31705
rect 15010 31696 15016 31699
rect 15068 31696 15074 31708
rect 15197 31705 15209 31739
rect 15243 31736 15255 31739
rect 15378 31736 15384 31748
rect 15243 31708 15384 31736
rect 15243 31705 15255 31708
rect 15197 31699 15255 31705
rect 15378 31696 15384 31708
rect 15436 31736 15442 31748
rect 15933 31739 15991 31745
rect 15933 31736 15945 31739
rect 15436 31708 15945 31736
rect 15436 31696 15442 31708
rect 15933 31705 15945 31708
rect 15979 31705 15991 31739
rect 15933 31699 15991 31705
rect 17494 31696 17500 31748
rect 17552 31736 17558 31748
rect 17972 31736 18000 31776
rect 18233 31773 18245 31776
rect 18279 31773 18291 31807
rect 18233 31767 18291 31773
rect 18322 31764 18328 31816
rect 18380 31804 18386 31816
rect 18509 31807 18567 31813
rect 18380 31776 18425 31804
rect 18380 31764 18386 31776
rect 18509 31773 18521 31807
rect 18555 31804 18567 31807
rect 18782 31804 18788 31816
rect 18555 31776 18788 31804
rect 18555 31773 18567 31776
rect 18509 31767 18567 31773
rect 18782 31764 18788 31776
rect 18840 31764 18846 31816
rect 19260 31813 19288 31844
rect 19245 31807 19303 31813
rect 19245 31773 19257 31807
rect 19291 31773 19303 31807
rect 19426 31804 19432 31816
rect 19387 31776 19432 31804
rect 19245 31767 19303 31773
rect 19426 31764 19432 31776
rect 19484 31764 19490 31816
rect 19536 31804 19564 31912
rect 20806 31900 20812 31912
rect 20864 31900 20870 31952
rect 22005 31943 22063 31949
rect 22005 31909 22017 31943
rect 22051 31940 22063 31943
rect 22278 31940 22284 31952
rect 22051 31912 22284 31940
rect 22051 31909 22063 31912
rect 22005 31903 22063 31909
rect 22278 31900 22284 31912
rect 22336 31900 22342 31952
rect 22646 31940 22652 31952
rect 22480 31912 22652 31940
rect 20714 31872 20720 31884
rect 20675 31844 20720 31872
rect 20714 31832 20720 31844
rect 20772 31832 20778 31884
rect 22370 31872 22376 31884
rect 20916 31844 22376 31872
rect 20916 31813 20944 31844
rect 22370 31832 22376 31844
rect 22428 31832 22434 31884
rect 22480 31881 22508 31912
rect 22646 31900 22652 31912
rect 22704 31900 22710 31952
rect 22756 31940 22784 31980
rect 22833 31977 22845 32011
rect 22879 32008 22891 32011
rect 23385 32011 23443 32017
rect 23385 32008 23397 32011
rect 22879 31980 23397 32008
rect 22879 31977 22891 31980
rect 22833 31971 22891 31977
rect 23385 31977 23397 31980
rect 23431 31977 23443 32011
rect 23385 31971 23443 31977
rect 24489 32011 24547 32017
rect 24489 31977 24501 32011
rect 24535 32008 24547 32011
rect 25498 32008 25504 32020
rect 24535 31980 25504 32008
rect 24535 31977 24547 31980
rect 24489 31971 24547 31977
rect 25498 31968 25504 31980
rect 25556 31968 25562 32020
rect 25590 31968 25596 32020
rect 25648 32008 25654 32020
rect 27893 32011 27951 32017
rect 25648 31980 25693 32008
rect 25648 31968 25654 31980
rect 27893 31977 27905 32011
rect 27939 32008 27951 32011
rect 28074 32008 28080 32020
rect 27939 31980 28080 32008
rect 27939 31977 27951 31980
rect 27893 31971 27951 31977
rect 28074 31968 28080 31980
rect 28132 31968 28138 32020
rect 28350 31968 28356 32020
rect 28408 32008 28414 32020
rect 28994 32008 29000 32020
rect 28408 31980 28856 32008
rect 28955 31980 29000 32008
rect 28408 31968 28414 31980
rect 25133 31943 25191 31949
rect 22756 31912 23244 31940
rect 22465 31875 22523 31881
rect 22465 31841 22477 31875
rect 22511 31841 22523 31875
rect 23106 31872 23112 31884
rect 22465 31835 22523 31841
rect 22664 31844 23112 31872
rect 20625 31807 20683 31813
rect 20625 31804 20637 31807
rect 19536 31776 20637 31804
rect 20625 31773 20637 31776
rect 20671 31773 20683 31807
rect 20625 31767 20683 31773
rect 20901 31807 20959 31813
rect 20901 31773 20913 31807
rect 20947 31773 20959 31807
rect 21082 31804 21088 31816
rect 21043 31776 21088 31804
rect 20901 31767 20959 31773
rect 21082 31764 21088 31776
rect 21140 31764 21146 31816
rect 21637 31807 21695 31813
rect 21637 31773 21649 31807
rect 21683 31804 21695 31807
rect 21726 31804 21732 31816
rect 21683 31776 21732 31804
rect 21683 31773 21695 31776
rect 21637 31767 21695 31773
rect 21726 31764 21732 31776
rect 21784 31764 21790 31816
rect 22664 31813 22692 31844
rect 23106 31832 23112 31844
rect 23164 31832 23170 31884
rect 22649 31807 22707 31813
rect 22649 31773 22661 31807
rect 22695 31773 22707 31807
rect 22649 31767 22707 31773
rect 17552 31708 18000 31736
rect 21821 31739 21879 31745
rect 17552 31696 17558 31708
rect 21821 31705 21833 31739
rect 21867 31736 21879 31739
rect 21910 31736 21916 31748
rect 21867 31708 21916 31736
rect 21867 31705 21879 31708
rect 21821 31699 21879 31705
rect 21910 31696 21916 31708
rect 21968 31696 21974 31748
rect 23216 31736 23244 31912
rect 25133 31909 25145 31943
rect 25179 31940 25191 31943
rect 26694 31940 26700 31952
rect 25179 31912 26700 31940
rect 25179 31909 25191 31912
rect 25133 31903 25191 31909
rect 26694 31900 26700 31912
rect 26752 31900 26758 31952
rect 27798 31900 27804 31952
rect 27856 31940 27862 31952
rect 28828 31940 28856 31980
rect 28994 31968 29000 31980
rect 29052 31968 29058 32020
rect 29914 31968 29920 32020
rect 29972 31968 29978 32020
rect 30101 32011 30159 32017
rect 30101 31977 30113 32011
rect 30147 32008 30159 32011
rect 30650 32008 30656 32020
rect 30147 31980 30656 32008
rect 30147 31977 30159 31980
rect 30101 31971 30159 31977
rect 30650 31968 30656 31980
rect 30708 31968 30714 32020
rect 30834 31968 30840 32020
rect 30892 32008 30898 32020
rect 31849 32011 31907 32017
rect 31849 32008 31861 32011
rect 30892 31980 31861 32008
rect 30892 31968 30898 31980
rect 31849 31977 31861 31980
rect 31895 31977 31907 32011
rect 31849 31971 31907 31977
rect 32582 31968 32588 32020
rect 32640 32008 32646 32020
rect 32769 32011 32827 32017
rect 32769 32008 32781 32011
rect 32640 31980 32781 32008
rect 32640 31968 32646 31980
rect 32769 31977 32781 31980
rect 32815 31977 32827 32011
rect 32769 31971 32827 31977
rect 34054 31968 34060 32020
rect 34112 32008 34118 32020
rect 34149 32011 34207 32017
rect 34149 32008 34161 32011
rect 34112 31980 34161 32008
rect 34112 31968 34118 31980
rect 34149 31977 34161 31980
rect 34195 31977 34207 32011
rect 34790 32008 34796 32020
rect 34751 31980 34796 32008
rect 34149 31971 34207 31977
rect 34790 31968 34796 31980
rect 34848 31968 34854 32020
rect 38378 31968 38384 32020
rect 38436 32008 38442 32020
rect 39853 32011 39911 32017
rect 39853 32008 39865 32011
rect 38436 31980 39865 32008
rect 38436 31968 38442 31980
rect 39853 31977 39865 31980
rect 39899 32008 39911 32011
rect 40402 32008 40408 32020
rect 39899 31980 40408 32008
rect 39899 31977 39911 31980
rect 39853 31971 39911 31977
rect 40402 31968 40408 31980
rect 40460 31968 40466 32020
rect 40678 31968 40684 32020
rect 40736 32008 40742 32020
rect 40957 32011 41015 32017
rect 40957 32008 40969 32011
rect 40736 31980 40969 32008
rect 40736 31968 40742 31980
rect 40957 31977 40969 31980
rect 41003 31977 41015 32011
rect 47670 32008 47676 32020
rect 47631 31980 47676 32008
rect 40957 31971 41015 31977
rect 47670 31968 47676 31980
rect 47728 31968 47734 32020
rect 29932 31940 29960 31968
rect 30742 31940 30748 31952
rect 27856 31912 28764 31940
rect 28828 31912 29960 31940
rect 30668 31912 30748 31940
rect 27856 31900 27862 31912
rect 23566 31872 23572 31884
rect 23527 31844 23572 31872
rect 23566 31832 23572 31844
rect 23624 31832 23630 31884
rect 24397 31875 24455 31881
rect 24397 31841 24409 31875
rect 24443 31872 24455 31875
rect 25682 31872 25688 31884
rect 24443 31844 25688 31872
rect 24443 31841 24455 31844
rect 24397 31835 24455 31841
rect 25682 31832 25688 31844
rect 25740 31872 25746 31884
rect 25961 31875 26019 31881
rect 25961 31872 25973 31875
rect 25740 31844 25973 31872
rect 25740 31832 25746 31844
rect 25961 31841 25973 31844
rect 26007 31841 26019 31875
rect 25961 31835 26019 31841
rect 27157 31875 27215 31881
rect 27157 31841 27169 31875
rect 27203 31872 27215 31875
rect 28258 31872 28264 31884
rect 27203 31844 28264 31872
rect 27203 31841 27215 31844
rect 27157 31835 27215 31841
rect 28258 31832 28264 31844
rect 28316 31832 28322 31884
rect 28350 31832 28356 31884
rect 28408 31872 28414 31884
rect 28736 31881 28764 31912
rect 28629 31875 28687 31881
rect 28629 31872 28641 31875
rect 28408 31844 28641 31872
rect 28408 31832 28414 31844
rect 28629 31841 28641 31844
rect 28675 31841 28687 31875
rect 28629 31835 28687 31841
rect 28721 31875 28779 31881
rect 28721 31841 28733 31875
rect 28767 31872 28779 31875
rect 29638 31872 29644 31884
rect 28767 31844 29500 31872
rect 29599 31844 29644 31872
rect 28767 31841 28779 31844
rect 28721 31835 28779 31841
rect 23293 31807 23351 31813
rect 23293 31773 23305 31807
rect 23339 31804 23351 31807
rect 23474 31804 23480 31816
rect 23339 31776 23480 31804
rect 23339 31773 23351 31776
rect 23293 31767 23351 31773
rect 23474 31764 23480 31776
rect 23532 31764 23538 31816
rect 24857 31807 24915 31813
rect 24857 31773 24869 31807
rect 24903 31804 24915 31807
rect 24946 31804 24952 31816
rect 24903 31776 24952 31804
rect 24903 31773 24915 31776
rect 24857 31767 24915 31773
rect 24946 31764 24952 31776
rect 25004 31764 25010 31816
rect 25774 31804 25780 31816
rect 25735 31776 25780 31804
rect 25774 31764 25780 31776
rect 25832 31764 25838 31816
rect 26602 31764 26608 31816
rect 26660 31804 26666 31816
rect 26973 31807 27031 31813
rect 26973 31804 26985 31807
rect 26660 31776 26985 31804
rect 26660 31764 26666 31776
rect 26973 31773 26985 31776
rect 27019 31804 27031 31807
rect 27062 31804 27068 31816
rect 27019 31776 27068 31804
rect 27019 31773 27031 31776
rect 26973 31767 27031 31773
rect 27062 31764 27068 31776
rect 27120 31804 27126 31816
rect 27614 31804 27620 31816
rect 27120 31776 27476 31804
rect 27575 31776 27620 31804
rect 27120 31764 27126 31776
rect 24302 31736 24308 31748
rect 23216 31708 24308 31736
rect 24302 31696 24308 31708
rect 24360 31696 24366 31748
rect 24670 31736 24676 31748
rect 24631 31708 24676 31736
rect 24670 31696 24676 31708
rect 24728 31696 24734 31748
rect 26786 31736 26792 31748
rect 26747 31708 26792 31736
rect 26786 31696 26792 31708
rect 26844 31696 26850 31748
rect 27448 31736 27476 31776
rect 27614 31764 27620 31776
rect 27672 31764 27678 31816
rect 27890 31804 27896 31816
rect 27851 31776 27896 31804
rect 27890 31764 27896 31776
rect 27948 31764 27954 31816
rect 28000 31776 28488 31804
rect 28000 31736 28028 31776
rect 27448 31708 28028 31736
rect 28460 31736 28488 31776
rect 28534 31764 28540 31816
rect 28592 31804 28598 31816
rect 28813 31807 28871 31813
rect 28592 31776 28637 31804
rect 28592 31764 28598 31776
rect 28813 31773 28825 31807
rect 28859 31804 28871 31807
rect 29362 31804 29368 31816
rect 28859 31776 29368 31804
rect 28859 31773 28871 31776
rect 28813 31767 28871 31773
rect 29362 31764 29368 31776
rect 29420 31764 29426 31816
rect 29472 31804 29500 31844
rect 29638 31832 29644 31844
rect 29696 31832 29702 31884
rect 29748 31881 29776 31912
rect 29733 31875 29791 31881
rect 29733 31841 29745 31875
rect 29779 31841 29791 31875
rect 29733 31835 29791 31841
rect 29917 31875 29975 31881
rect 29917 31841 29929 31875
rect 29963 31872 29975 31875
rect 30006 31872 30012 31884
rect 29963 31844 30012 31872
rect 29963 31841 29975 31844
rect 29917 31835 29975 31841
rect 30006 31832 30012 31844
rect 30064 31832 30070 31884
rect 30668 31881 30696 31912
rect 30742 31900 30748 31912
rect 30800 31900 30806 31952
rect 35434 31940 35440 31952
rect 35176 31912 35440 31940
rect 30653 31875 30711 31881
rect 30653 31841 30665 31875
rect 30699 31841 30711 31875
rect 32214 31872 32220 31884
rect 32175 31844 32220 31872
rect 30653 31835 30711 31841
rect 32214 31832 32220 31844
rect 32272 31832 32278 31884
rect 33873 31875 33931 31881
rect 32324 31844 32996 31872
rect 29825 31807 29883 31813
rect 29472 31776 29684 31804
rect 28994 31736 29000 31748
rect 28460 31708 29000 31736
rect 28994 31696 29000 31708
rect 29052 31696 29058 31748
rect 29656 31736 29684 31776
rect 29825 31773 29837 31807
rect 29871 31804 29883 31807
rect 29871 31776 29905 31804
rect 29871 31773 29883 31776
rect 29825 31767 29883 31773
rect 29840 31736 29868 31767
rect 30466 31764 30472 31816
rect 30524 31804 30530 31816
rect 30561 31807 30619 31813
rect 30561 31804 30573 31807
rect 30524 31776 30573 31804
rect 30524 31764 30530 31776
rect 30561 31773 30573 31776
rect 30607 31773 30619 31807
rect 30742 31804 30748 31816
rect 30703 31776 30748 31804
rect 30561 31767 30619 31773
rect 30742 31764 30748 31776
rect 30800 31764 30806 31816
rect 32122 31804 32128 31816
rect 32083 31776 32128 31804
rect 32122 31764 32128 31776
rect 32180 31764 32186 31816
rect 32324 31804 32352 31844
rect 32968 31813 32996 31844
rect 33873 31841 33885 31875
rect 33919 31872 33931 31875
rect 33962 31872 33968 31884
rect 33919 31844 33968 31872
rect 33919 31841 33931 31844
rect 33873 31835 33931 31841
rect 33962 31832 33968 31844
rect 34020 31832 34026 31884
rect 34057 31875 34115 31881
rect 34057 31841 34069 31875
rect 34103 31872 34115 31875
rect 34698 31872 34704 31884
rect 34103 31844 34704 31872
rect 34103 31841 34115 31844
rect 34057 31835 34115 31841
rect 34698 31832 34704 31844
rect 34756 31832 34762 31884
rect 32232 31776 32352 31804
rect 32953 31807 33011 31813
rect 32232 31748 32260 31776
rect 32953 31773 32965 31807
rect 32999 31773 33011 31807
rect 32953 31767 33011 31773
rect 33045 31807 33103 31813
rect 33045 31773 33057 31807
rect 33091 31773 33103 31807
rect 33045 31767 33103 31773
rect 34149 31807 34207 31813
rect 34149 31773 34161 31807
rect 34195 31804 34207 31807
rect 34514 31804 34520 31816
rect 34195 31776 34520 31804
rect 34195 31773 34207 31776
rect 34149 31767 34207 31773
rect 29656 31708 29868 31736
rect 30190 31696 30196 31748
rect 30248 31736 30254 31748
rect 30248 31708 32168 31736
rect 30248 31696 30254 31708
rect 14829 31671 14887 31677
rect 14829 31637 14841 31671
rect 14875 31637 14887 31671
rect 14829 31631 14887 31637
rect 17313 31671 17371 31677
rect 17313 31637 17325 31671
rect 17359 31668 17371 31671
rect 17402 31668 17408 31680
rect 17359 31640 17408 31668
rect 17359 31637 17371 31640
rect 17313 31631 17371 31637
rect 17402 31628 17408 31640
rect 17460 31668 17466 31680
rect 17586 31668 17592 31680
rect 17460 31640 17592 31668
rect 17460 31628 17466 31640
rect 17586 31628 17592 31640
rect 17644 31628 17650 31680
rect 17865 31671 17923 31677
rect 17865 31637 17877 31671
rect 17911 31668 17923 31671
rect 17954 31668 17960 31680
rect 17911 31640 17960 31668
rect 17911 31637 17923 31640
rect 17865 31631 17923 31637
rect 17954 31628 17960 31640
rect 18012 31628 18018 31680
rect 19981 31671 20039 31677
rect 19981 31637 19993 31671
rect 20027 31668 20039 31671
rect 22094 31668 22100 31680
rect 20027 31640 22100 31668
rect 20027 31637 20039 31640
rect 19981 31631 20039 31637
rect 22094 31628 22100 31640
rect 22152 31628 22158 31680
rect 23845 31671 23903 31677
rect 23845 31637 23857 31671
rect 23891 31668 23903 31671
rect 24765 31671 24823 31677
rect 24765 31668 24777 31671
rect 23891 31640 24777 31668
rect 23891 31637 23903 31640
rect 23845 31631 23903 31637
rect 24765 31637 24777 31640
rect 24811 31637 24823 31671
rect 27706 31668 27712 31680
rect 27667 31640 27712 31668
rect 24765 31631 24823 31637
rect 27706 31628 27712 31640
rect 27764 31628 27770 31680
rect 30650 31628 30656 31680
rect 30708 31668 30714 31680
rect 31294 31668 31300 31680
rect 30708 31640 31300 31668
rect 30708 31628 30714 31640
rect 31294 31628 31300 31640
rect 31352 31628 31358 31680
rect 32140 31668 32168 31708
rect 32214 31696 32220 31748
rect 32272 31696 32278 31748
rect 32950 31668 32956 31680
rect 32140 31640 32956 31668
rect 32950 31628 32956 31640
rect 33008 31668 33014 31680
rect 33060 31668 33088 31767
rect 34514 31764 34520 31776
rect 34572 31764 34578 31816
rect 35176 31813 35204 31912
rect 35434 31900 35440 31912
rect 35492 31900 35498 31952
rect 35894 31900 35900 31952
rect 35952 31940 35958 31952
rect 35952 31912 38654 31940
rect 35952 31900 35958 31912
rect 38626 31884 38654 31912
rect 35710 31872 35716 31884
rect 35289 31844 35716 31872
rect 35289 31813 35317 31844
rect 35710 31832 35716 31844
rect 35768 31832 35774 31884
rect 36538 31872 36544 31884
rect 36499 31844 36544 31872
rect 36538 31832 36544 31844
rect 36596 31832 36602 31884
rect 37826 31872 37832 31884
rect 37200 31844 37832 31872
rect 35049 31807 35107 31813
rect 35049 31773 35061 31807
rect 35095 31804 35107 31807
rect 35142 31807 35204 31813
rect 35095 31773 35112 31804
rect 35049 31767 35112 31773
rect 35142 31773 35154 31807
rect 35188 31776 35204 31807
rect 35253 31807 35317 31813
rect 35188 31773 35200 31776
rect 35142 31767 35200 31773
rect 35253 31773 35265 31807
rect 35299 31776 35317 31807
rect 35437 31807 35495 31813
rect 35299 31773 35311 31776
rect 35253 31767 35311 31773
rect 35437 31773 35449 31807
rect 35483 31804 35495 31807
rect 35894 31804 35900 31816
rect 35483 31776 35900 31804
rect 35483 31773 35495 31776
rect 35437 31767 35495 31773
rect 35084 31736 35112 31767
rect 35894 31764 35900 31776
rect 35952 31764 35958 31816
rect 36722 31804 36728 31816
rect 36683 31776 36728 31804
rect 36722 31764 36728 31776
rect 36780 31764 36786 31816
rect 37200 31813 37228 31844
rect 37826 31832 37832 31844
rect 37884 31832 37890 31884
rect 38197 31875 38255 31881
rect 38197 31841 38209 31875
rect 38243 31872 38255 31875
rect 38470 31872 38476 31884
rect 38243 31844 38476 31872
rect 38243 31841 38255 31844
rect 38197 31835 38255 31841
rect 38470 31832 38476 31844
rect 38528 31832 38534 31884
rect 38626 31872 38660 31884
rect 38567 31844 38660 31872
rect 38654 31832 38660 31844
rect 38712 31832 38718 31884
rect 37185 31807 37243 31813
rect 37185 31773 37197 31807
rect 37231 31773 37243 31807
rect 37458 31804 37464 31816
rect 37419 31776 37464 31804
rect 37185 31767 37243 31773
rect 37458 31764 37464 31776
rect 37516 31764 37522 31816
rect 38838 31804 38844 31816
rect 38626 31776 38844 31804
rect 35342 31736 35348 31748
rect 35084 31708 35348 31736
rect 35342 31696 35348 31708
rect 35400 31696 35406 31748
rect 36265 31739 36323 31745
rect 36265 31705 36277 31739
rect 36311 31705 36323 31739
rect 36740 31736 36768 31764
rect 37642 31736 37648 31748
rect 36740 31708 37648 31736
rect 36265 31699 36323 31705
rect 33008 31640 33088 31668
rect 33008 31628 33014 31640
rect 33318 31628 33324 31680
rect 33376 31668 33382 31680
rect 36280 31668 36308 31699
rect 37642 31696 37648 31708
rect 37700 31736 37706 31748
rect 38626 31736 38654 31776
rect 38838 31764 38844 31776
rect 38896 31804 38902 31816
rect 39209 31807 39267 31813
rect 39209 31804 39221 31807
rect 38896 31776 39221 31804
rect 38896 31764 38902 31776
rect 39209 31773 39221 31776
rect 39255 31773 39267 31807
rect 39209 31767 39267 31773
rect 37700 31708 38654 31736
rect 37700 31696 37706 31708
rect 33376 31640 36308 31668
rect 33376 31628 33382 31640
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 10965 31467 11023 31473
rect 10965 31433 10977 31467
rect 11011 31464 11023 31467
rect 13541 31467 13599 31473
rect 11011 31436 12572 31464
rect 11011 31433 11023 31436
rect 10965 31427 11023 31433
rect 12342 31396 12348 31408
rect 12303 31368 12348 31396
rect 12342 31356 12348 31368
rect 12400 31356 12406 31408
rect 12544 31340 12572 31436
rect 13541 31433 13553 31467
rect 13587 31464 13599 31467
rect 13814 31464 13820 31476
rect 13587 31436 13820 31464
rect 13587 31433 13599 31436
rect 13541 31427 13599 31433
rect 13814 31424 13820 31436
rect 13872 31424 13878 31476
rect 13909 31467 13967 31473
rect 13909 31433 13921 31467
rect 13955 31464 13967 31467
rect 15010 31464 15016 31476
rect 13955 31436 15016 31464
rect 13955 31433 13967 31436
rect 13909 31427 13967 31433
rect 15010 31424 15016 31436
rect 15068 31424 15074 31476
rect 15194 31424 15200 31476
rect 15252 31464 15258 31476
rect 16482 31464 16488 31476
rect 15252 31436 16488 31464
rect 15252 31424 15258 31436
rect 16482 31424 16488 31436
rect 16540 31464 16546 31476
rect 16853 31467 16911 31473
rect 16853 31464 16865 31467
rect 16540 31436 16865 31464
rect 16540 31424 16546 31436
rect 16853 31433 16865 31436
rect 16899 31433 16911 31467
rect 17862 31464 17868 31476
rect 17823 31436 17868 31464
rect 16853 31427 16911 31433
rect 17862 31424 17868 31436
rect 17920 31424 17926 31476
rect 19797 31467 19855 31473
rect 17972 31436 19380 31464
rect 15838 31396 15844 31408
rect 12728 31368 15056 31396
rect 11885 31331 11943 31337
rect 11885 31297 11897 31331
rect 11931 31328 11943 31331
rect 11931 31300 12434 31328
rect 11931 31297 11943 31300
rect 11885 31291 11943 31297
rect 12406 31260 12434 31300
rect 12526 31288 12532 31340
rect 12584 31328 12590 31340
rect 12584 31300 12629 31328
rect 12584 31288 12590 31300
rect 12728 31260 12756 31368
rect 15028 31340 15056 31368
rect 15120 31368 15844 31396
rect 13446 31328 13452 31340
rect 13359 31300 13452 31328
rect 13446 31288 13452 31300
rect 13504 31288 13510 31340
rect 13722 31328 13728 31340
rect 13683 31300 13728 31328
rect 13722 31288 13728 31300
rect 13780 31288 13786 31340
rect 14826 31328 14832 31340
rect 14787 31300 14832 31328
rect 14826 31288 14832 31300
rect 14884 31288 14890 31340
rect 15010 31328 15016 31340
rect 14971 31300 15016 31328
rect 15010 31288 15016 31300
rect 15068 31288 15074 31340
rect 15120 31337 15148 31368
rect 15838 31356 15844 31368
rect 15896 31396 15902 31408
rect 17972 31396 18000 31436
rect 19242 31396 19248 31408
rect 15896 31368 18000 31396
rect 18800 31368 19248 31396
rect 15896 31356 15902 31368
rect 15105 31331 15163 31337
rect 15105 31297 15117 31331
rect 15151 31297 15163 31331
rect 15105 31291 15163 31297
rect 15749 31331 15807 31337
rect 15749 31297 15761 31331
rect 15795 31297 15807 31331
rect 15749 31291 15807 31297
rect 12406 31232 12756 31260
rect 13464 31260 13492 31288
rect 14182 31260 14188 31272
rect 13464 31232 14188 31260
rect 14182 31220 14188 31232
rect 14240 31260 14246 31272
rect 15194 31260 15200 31272
rect 14240 31232 15200 31260
rect 14240 31220 14246 31232
rect 15194 31220 15200 31232
rect 15252 31260 15258 31272
rect 15565 31263 15623 31269
rect 15565 31260 15577 31263
rect 15252 31232 15577 31260
rect 15252 31220 15258 31232
rect 15565 31229 15577 31232
rect 15611 31229 15623 31263
rect 15565 31223 15623 31229
rect 15105 31195 15163 31201
rect 15105 31161 15117 31195
rect 15151 31192 15163 31195
rect 15764 31192 15792 31291
rect 17310 31288 17316 31340
rect 17368 31328 17374 31340
rect 17405 31331 17463 31337
rect 17405 31328 17417 31331
rect 17368 31300 17417 31328
rect 17368 31288 17374 31300
rect 17405 31297 17417 31300
rect 17451 31297 17463 31331
rect 17405 31291 17463 31297
rect 17494 31288 17500 31340
rect 17552 31328 17558 31340
rect 17681 31331 17739 31337
rect 17552 31300 17597 31328
rect 17552 31288 17558 31300
rect 17681 31297 17693 31331
rect 17727 31328 17739 31331
rect 18046 31328 18052 31340
rect 17727 31300 18052 31328
rect 17727 31297 17739 31300
rect 17681 31291 17739 31297
rect 18046 31288 18052 31300
rect 18104 31288 18110 31340
rect 18800 31337 18828 31368
rect 19242 31356 19248 31368
rect 19300 31356 19306 31408
rect 19352 31396 19380 31436
rect 19797 31433 19809 31467
rect 19843 31464 19855 31467
rect 19978 31464 19984 31476
rect 19843 31436 19984 31464
rect 19843 31433 19855 31436
rect 19797 31427 19855 31433
rect 19978 31424 19984 31436
rect 20036 31424 20042 31476
rect 21082 31464 21088 31476
rect 21043 31436 21088 31464
rect 21082 31424 21088 31436
rect 21140 31424 21146 31476
rect 23290 31424 23296 31476
rect 23348 31464 23354 31476
rect 23385 31467 23443 31473
rect 23385 31464 23397 31467
rect 23348 31436 23397 31464
rect 23348 31424 23354 31436
rect 23385 31433 23397 31436
rect 23431 31433 23443 31467
rect 24210 31464 24216 31476
rect 24171 31436 24216 31464
rect 23385 31427 23443 31433
rect 24210 31424 24216 31436
rect 24268 31424 24274 31476
rect 24854 31424 24860 31476
rect 24912 31424 24918 31476
rect 24946 31424 24952 31476
rect 25004 31464 25010 31476
rect 25501 31467 25559 31473
rect 25501 31464 25513 31467
rect 25004 31436 25513 31464
rect 25004 31424 25010 31436
rect 25501 31433 25513 31436
rect 25547 31433 25559 31467
rect 25501 31427 25559 31433
rect 26234 31424 26240 31476
rect 26292 31464 26298 31476
rect 27246 31464 27252 31476
rect 26292 31436 27252 31464
rect 26292 31424 26298 31436
rect 27246 31424 27252 31436
rect 27304 31424 27310 31476
rect 27522 31424 27528 31476
rect 27580 31424 27586 31476
rect 27614 31424 27620 31476
rect 27672 31473 27678 31476
rect 27672 31464 27681 31473
rect 27672 31436 27717 31464
rect 27672 31427 27681 31436
rect 27672 31424 27678 31427
rect 27982 31424 27988 31476
rect 28040 31464 28046 31476
rect 28353 31467 28411 31473
rect 28353 31464 28365 31467
rect 28040 31436 28365 31464
rect 28040 31424 28046 31436
rect 28353 31433 28365 31436
rect 28399 31433 28411 31467
rect 28994 31464 29000 31476
rect 28955 31436 29000 31464
rect 28353 31427 28411 31433
rect 28994 31424 29000 31436
rect 29052 31424 29058 31476
rect 29454 31464 29460 31476
rect 29415 31436 29460 31464
rect 29454 31424 29460 31436
rect 29512 31424 29518 31476
rect 30466 31424 30472 31476
rect 30524 31464 30530 31476
rect 31021 31467 31079 31473
rect 31021 31464 31033 31467
rect 30524 31436 31033 31464
rect 30524 31424 30530 31436
rect 31021 31433 31033 31436
rect 31067 31433 31079 31467
rect 31021 31427 31079 31433
rect 32309 31467 32367 31473
rect 32309 31433 32321 31467
rect 32355 31464 32367 31467
rect 32858 31464 32864 31476
rect 32355 31436 32864 31464
rect 32355 31433 32367 31436
rect 32309 31427 32367 31433
rect 32858 31424 32864 31436
rect 32916 31424 32922 31476
rect 34514 31424 34520 31476
rect 34572 31464 34578 31476
rect 35526 31464 35532 31476
rect 34572 31436 35532 31464
rect 34572 31424 34578 31436
rect 35526 31424 35532 31436
rect 35584 31424 35590 31476
rect 37642 31464 37648 31476
rect 37603 31436 37648 31464
rect 37642 31424 37648 31436
rect 37700 31424 37706 31476
rect 38838 31464 38844 31476
rect 38799 31436 38844 31464
rect 38838 31424 38844 31436
rect 38896 31424 38902 31476
rect 39942 31424 39948 31476
rect 40000 31464 40006 31476
rect 40497 31467 40555 31473
rect 40497 31464 40509 31467
rect 40000 31436 40509 31464
rect 40000 31424 40006 31436
rect 40497 31433 40509 31436
rect 40543 31433 40555 31467
rect 40497 31427 40555 31433
rect 20625 31399 20683 31405
rect 19352 31368 20024 31396
rect 18785 31331 18843 31337
rect 18785 31297 18797 31331
rect 18831 31297 18843 31331
rect 18966 31328 18972 31340
rect 18927 31300 18972 31328
rect 18785 31291 18843 31297
rect 18966 31288 18972 31300
rect 19024 31328 19030 31340
rect 19705 31331 19763 31337
rect 19705 31328 19717 31331
rect 19024 31300 19717 31328
rect 19024 31288 19030 31300
rect 19705 31297 19717 31300
rect 19751 31297 19763 31331
rect 19886 31328 19892 31340
rect 19847 31300 19892 31328
rect 19705 31291 19763 31297
rect 19886 31288 19892 31300
rect 19944 31288 19950 31340
rect 19996 31328 20024 31368
rect 20625 31365 20637 31399
rect 20671 31396 20683 31399
rect 21450 31396 21456 31408
rect 20671 31368 21456 31396
rect 20671 31365 20683 31368
rect 20625 31359 20683 31365
rect 21450 31356 21456 31368
rect 21508 31356 21514 31408
rect 22094 31356 22100 31408
rect 22152 31396 22158 31408
rect 22465 31399 22523 31405
rect 22465 31396 22477 31399
rect 22152 31368 22477 31396
rect 22152 31356 22158 31368
rect 22465 31365 22477 31368
rect 22511 31365 22523 31399
rect 22465 31359 22523 31365
rect 22554 31356 22560 31408
rect 22612 31396 22618 31408
rect 22833 31399 22891 31405
rect 22612 31368 22784 31396
rect 22612 31356 22618 31368
rect 20901 31331 20959 31337
rect 19996 31300 20852 31328
rect 19245 31263 19303 31269
rect 19245 31229 19257 31263
rect 19291 31260 19303 31263
rect 19904 31260 19932 31288
rect 19291 31232 19932 31260
rect 20717 31263 20775 31269
rect 19291 31229 19303 31232
rect 19245 31223 19303 31229
rect 20717 31229 20729 31263
rect 20763 31229 20775 31263
rect 20824 31260 20852 31300
rect 20901 31297 20913 31331
rect 20947 31328 20959 31331
rect 20990 31328 20996 31340
rect 20947 31300 20996 31328
rect 20947 31297 20959 31300
rect 20901 31291 20959 31297
rect 20990 31288 20996 31300
rect 21048 31288 21054 31340
rect 22002 31288 22008 31340
rect 22060 31328 22066 31340
rect 22278 31328 22284 31340
rect 22060 31300 22284 31328
rect 22060 31288 22066 31300
rect 22278 31288 22284 31300
rect 22336 31328 22342 31340
rect 22649 31331 22707 31337
rect 22649 31328 22661 31331
rect 22336 31300 22661 31328
rect 22336 31288 22342 31300
rect 22649 31297 22661 31300
rect 22695 31297 22707 31331
rect 22756 31328 22784 31368
rect 22833 31365 22845 31399
rect 22879 31396 22891 31399
rect 22879 31368 23520 31396
rect 22879 31365 22891 31368
rect 22833 31359 22891 31365
rect 23492 31337 23520 31368
rect 23293 31331 23351 31337
rect 23293 31328 23305 31331
rect 22756 31300 23305 31328
rect 22649 31291 22707 31297
rect 23293 31297 23305 31300
rect 23339 31297 23351 31331
rect 23293 31291 23351 31297
rect 23477 31331 23535 31337
rect 23477 31297 23489 31331
rect 23523 31297 23535 31331
rect 24228 31328 24256 31424
rect 24673 31399 24731 31405
rect 24673 31365 24685 31399
rect 24719 31396 24731 31399
rect 24872 31396 24900 31424
rect 24719 31368 24900 31396
rect 25041 31399 25099 31405
rect 24719 31365 24731 31368
rect 24673 31359 24731 31365
rect 25041 31365 25053 31399
rect 25087 31396 25099 31399
rect 25774 31396 25780 31408
rect 25087 31368 25780 31396
rect 25087 31365 25099 31368
rect 25041 31359 25099 31365
rect 25774 31356 25780 31368
rect 25832 31356 25838 31408
rect 26050 31356 26056 31408
rect 26108 31396 26114 31408
rect 27540 31396 27568 31424
rect 27709 31399 27767 31405
rect 27709 31396 27721 31399
rect 26108 31368 27476 31396
rect 27540 31368 27721 31396
rect 26108 31356 26114 31368
rect 24857 31331 24915 31337
rect 24857 31328 24869 31331
rect 24228 31300 24869 31328
rect 23477 31291 23535 31297
rect 24857 31297 24869 31300
rect 24903 31297 24915 31331
rect 24857 31291 24915 31297
rect 25501 31331 25559 31337
rect 25501 31297 25513 31331
rect 25547 31297 25559 31331
rect 25501 31291 25559 31297
rect 25685 31331 25743 31337
rect 25685 31297 25697 31331
rect 25731 31328 25743 31331
rect 26145 31331 26203 31337
rect 26145 31328 26157 31331
rect 25731 31300 26157 31328
rect 25731 31297 25743 31300
rect 25685 31291 25743 31297
rect 26145 31297 26157 31300
rect 26191 31328 26203 31331
rect 26234 31328 26240 31340
rect 26191 31300 26240 31328
rect 26191 31297 26203 31300
rect 26145 31291 26203 31297
rect 25516 31260 25544 31291
rect 26234 31288 26240 31300
rect 26292 31288 26298 31340
rect 26329 31331 26387 31337
rect 26329 31297 26341 31331
rect 26375 31328 26387 31331
rect 27062 31328 27068 31340
rect 26375 31300 27068 31328
rect 26375 31297 26387 31300
rect 26329 31291 26387 31297
rect 26344 31260 26372 31291
rect 27062 31288 27068 31300
rect 27120 31288 27126 31340
rect 27448 31328 27476 31368
rect 27709 31365 27721 31368
rect 27755 31365 27767 31399
rect 29086 31396 29092 31408
rect 27709 31359 27767 31365
rect 28092 31368 29092 31396
rect 27525 31331 27583 31337
rect 27525 31328 27537 31331
rect 27448 31300 27537 31328
rect 27525 31297 27537 31300
rect 27571 31297 27583 31331
rect 27525 31291 27583 31297
rect 27801 31331 27859 31337
rect 27801 31297 27813 31331
rect 27847 31328 27859 31331
rect 27890 31328 27896 31340
rect 27847 31300 27896 31328
rect 27847 31297 27859 31300
rect 27801 31291 27859 31297
rect 20824 31232 22094 31260
rect 25516 31232 26372 31260
rect 27540 31260 27568 31291
rect 27890 31288 27896 31300
rect 27948 31288 27954 31340
rect 28092 31260 28120 31368
rect 29086 31356 29092 31368
rect 29144 31356 29150 31408
rect 31478 31396 31484 31408
rect 29472 31368 31484 31396
rect 29472 31340 29500 31368
rect 28258 31328 28264 31340
rect 28219 31300 28264 31328
rect 28258 31288 28264 31300
rect 28316 31288 28322 31340
rect 28350 31288 28356 31340
rect 28408 31328 28414 31340
rect 28445 31331 28503 31337
rect 28445 31328 28457 31331
rect 28408 31300 28457 31328
rect 28408 31288 28414 31300
rect 28445 31297 28457 31300
rect 28491 31297 28503 31331
rect 28445 31291 28503 31297
rect 29454 31288 29460 31340
rect 29512 31288 29518 31340
rect 29917 31331 29975 31337
rect 29917 31297 29929 31331
rect 29963 31328 29975 31331
rect 30006 31328 30012 31340
rect 29963 31300 30012 31328
rect 29963 31297 29975 31300
rect 29917 31291 29975 31297
rect 30006 31288 30012 31300
rect 30064 31288 30070 31340
rect 30392 31337 30420 31368
rect 31478 31356 31484 31368
rect 31536 31356 31542 31408
rect 32585 31399 32643 31405
rect 32585 31365 32597 31399
rect 32631 31396 32643 31399
rect 33778 31396 33784 31408
rect 32631 31368 33784 31396
rect 32631 31365 32643 31368
rect 32585 31359 32643 31365
rect 33778 31356 33784 31368
rect 33836 31356 33842 31408
rect 35342 31396 35348 31408
rect 35176 31368 35348 31396
rect 30377 31331 30435 31337
rect 30377 31297 30389 31331
rect 30423 31297 30435 31331
rect 30377 31291 30435 31297
rect 30561 31331 30619 31337
rect 30561 31297 30573 31331
rect 30607 31328 30619 31331
rect 30650 31328 30656 31340
rect 30607 31300 30656 31328
rect 30607 31297 30619 31300
rect 30561 31291 30619 31297
rect 30650 31288 30656 31300
rect 30708 31288 30714 31340
rect 31018 31328 31024 31340
rect 30979 31300 31024 31328
rect 31018 31288 31024 31300
rect 31076 31288 31082 31340
rect 31205 31331 31263 31337
rect 31205 31297 31217 31331
rect 31251 31328 31263 31331
rect 31386 31328 31392 31340
rect 31251 31300 31392 31328
rect 31251 31297 31263 31300
rect 31205 31291 31263 31297
rect 31386 31288 31392 31300
rect 31444 31288 31450 31340
rect 32122 31288 32128 31340
rect 32180 31328 32186 31340
rect 32493 31331 32551 31337
rect 32493 31328 32505 31331
rect 32180 31300 32505 31328
rect 32180 31288 32186 31300
rect 32493 31297 32505 31300
rect 32539 31297 32551 31331
rect 32674 31328 32680 31340
rect 32635 31300 32680 31328
rect 32493 31291 32551 31297
rect 27540 31232 28120 31260
rect 20717 31223 20775 31229
rect 15151 31164 15792 31192
rect 18969 31195 19027 31201
rect 15151 31161 15163 31164
rect 15105 31155 15163 31161
rect 18969 31161 18981 31195
rect 19015 31192 19027 31195
rect 20070 31192 20076 31204
rect 19015 31164 20076 31192
rect 19015 31161 19027 31164
rect 18969 31155 19027 31161
rect 20070 31152 20076 31164
rect 20128 31192 20134 31204
rect 20732 31192 20760 31223
rect 20128 31164 20760 31192
rect 22066 31192 22094 31232
rect 28166 31220 28172 31272
rect 28224 31260 28230 31272
rect 28534 31260 28540 31272
rect 28224 31232 28540 31260
rect 28224 31220 28230 31232
rect 28534 31220 28540 31232
rect 28592 31260 28598 31272
rect 31478 31260 31484 31272
rect 28592 31232 31484 31260
rect 28592 31220 28598 31232
rect 31478 31220 31484 31232
rect 31536 31220 31542 31272
rect 32508 31260 32536 31291
rect 32674 31288 32680 31300
rect 32732 31288 32738 31340
rect 32766 31288 32772 31340
rect 32824 31337 32830 31340
rect 32824 31331 32853 31337
rect 32841 31297 32853 31331
rect 33134 31328 33140 31340
rect 32824 31291 32853 31297
rect 32892 31300 33140 31328
rect 32824 31288 32830 31291
rect 32892 31260 32920 31300
rect 33134 31288 33140 31300
rect 33192 31288 33198 31340
rect 33410 31328 33416 31340
rect 33371 31300 33416 31328
rect 33410 31288 33416 31300
rect 33468 31288 33474 31340
rect 35176 31337 35204 31368
rect 35342 31356 35348 31368
rect 35400 31396 35406 31408
rect 38562 31396 38568 31408
rect 35400 31368 38568 31396
rect 35400 31356 35406 31368
rect 38562 31356 38568 31368
rect 38620 31356 38626 31408
rect 34057 31331 34115 31337
rect 34057 31297 34069 31331
rect 34103 31297 34115 31331
rect 34057 31291 34115 31297
rect 35161 31331 35219 31337
rect 35161 31297 35173 31331
rect 35207 31297 35219 31331
rect 35161 31291 35219 31297
rect 37461 31331 37519 31337
rect 37461 31297 37473 31331
rect 37507 31328 37519 31331
rect 37642 31328 37648 31340
rect 37507 31300 37648 31328
rect 37507 31297 37519 31300
rect 37461 31291 37519 31297
rect 32508 31232 32920 31260
rect 32953 31263 33011 31269
rect 32953 31229 32965 31263
rect 32999 31260 33011 31263
rect 33505 31263 33563 31269
rect 33505 31260 33517 31263
rect 32999 31232 33517 31260
rect 32999 31229 33011 31232
rect 32953 31223 33011 31229
rect 33505 31229 33517 31232
rect 33551 31229 33563 31263
rect 33505 31223 33563 31229
rect 33318 31192 33324 31204
rect 22066 31164 33324 31192
rect 20128 31152 20134 31164
rect 33318 31152 33324 31164
rect 33376 31152 33382 31204
rect 12713 31127 12771 31133
rect 12713 31093 12725 31127
rect 12759 31124 12771 31127
rect 12986 31124 12992 31136
rect 12759 31096 12992 31124
rect 12759 31093 12771 31096
rect 12713 31087 12771 31093
rect 12986 31084 12992 31096
rect 13044 31084 13050 31136
rect 15933 31127 15991 31133
rect 15933 31093 15945 31127
rect 15979 31124 15991 31127
rect 16390 31124 16396 31136
rect 15979 31096 16396 31124
rect 15979 31093 15991 31096
rect 15933 31087 15991 31093
rect 16390 31084 16396 31096
rect 16448 31084 16454 31136
rect 16482 31084 16488 31136
rect 16540 31124 16546 31136
rect 19794 31124 19800 31136
rect 16540 31096 19800 31124
rect 16540 31084 16546 31096
rect 19794 31084 19800 31096
rect 19852 31084 19858 31136
rect 19978 31084 19984 31136
rect 20036 31124 20042 31136
rect 20438 31124 20444 31136
rect 20036 31096 20444 31124
rect 20036 31084 20042 31096
rect 20438 31084 20444 31096
rect 20496 31124 20502 31136
rect 20625 31127 20683 31133
rect 20625 31124 20637 31127
rect 20496 31096 20637 31124
rect 20496 31084 20502 31096
rect 20625 31093 20637 31096
rect 20671 31093 20683 31127
rect 22002 31124 22008 31136
rect 21963 31096 22008 31124
rect 20625 31087 20683 31093
rect 22002 31084 22008 31096
rect 22060 31084 22066 31136
rect 25498 31084 25504 31136
rect 25556 31124 25562 31136
rect 26145 31127 26203 31133
rect 26145 31124 26157 31127
rect 25556 31096 26157 31124
rect 25556 31084 25562 31096
rect 26145 31093 26157 31096
rect 26191 31093 26203 31127
rect 27062 31124 27068 31136
rect 27023 31096 27068 31124
rect 26145 31087 26203 31093
rect 27062 31084 27068 31096
rect 27120 31084 27126 31136
rect 29638 31124 29644 31136
rect 29599 31096 29644 31124
rect 29638 31084 29644 31096
rect 29696 31124 29702 31136
rect 30377 31127 30435 31133
rect 30377 31124 30389 31127
rect 29696 31096 30389 31124
rect 29696 31084 29702 31096
rect 30377 31093 30389 31096
rect 30423 31093 30435 31127
rect 30377 31087 30435 31093
rect 31478 31084 31484 31136
rect 31536 31124 31542 31136
rect 34072 31124 34100 31291
rect 37642 31288 37648 31300
rect 37700 31288 37706 31340
rect 37737 31331 37795 31337
rect 37737 31297 37749 31331
rect 37783 31328 37795 31331
rect 37826 31328 37832 31340
rect 37783 31300 37832 31328
rect 37783 31297 37795 31300
rect 37737 31291 37795 31297
rect 37826 31288 37832 31300
rect 37884 31288 37890 31340
rect 34146 31220 34152 31272
rect 34204 31260 34210 31272
rect 34241 31263 34299 31269
rect 34241 31260 34253 31263
rect 34204 31232 34253 31260
rect 34204 31220 34210 31232
rect 34241 31229 34253 31232
rect 34287 31229 34299 31263
rect 34241 31223 34299 31229
rect 35253 31263 35311 31269
rect 35253 31229 35265 31263
rect 35299 31260 35311 31263
rect 35434 31260 35440 31272
rect 35299 31232 35440 31260
rect 35299 31229 35311 31232
rect 35253 31223 35311 31229
rect 35434 31220 35440 31232
rect 35492 31220 35498 31272
rect 36078 31124 36084 31136
rect 31536 31096 34100 31124
rect 36039 31096 36084 31124
rect 31536 31084 31542 31096
rect 36078 31084 36084 31096
rect 36136 31084 36142 31136
rect 36446 31084 36452 31136
rect 36504 31124 36510 31136
rect 36541 31127 36599 31133
rect 36541 31124 36553 31127
rect 36504 31096 36553 31124
rect 36504 31084 36510 31096
rect 36541 31093 36553 31096
rect 36587 31093 36599 31127
rect 37274 31124 37280 31136
rect 37235 31096 37280 31124
rect 36541 31087 36599 31093
rect 37274 31084 37280 31096
rect 37332 31084 37338 31136
rect 38289 31127 38347 31133
rect 38289 31093 38301 31127
rect 38335 31124 38347 31127
rect 38654 31124 38660 31136
rect 38335 31096 38660 31124
rect 38335 31093 38347 31096
rect 38289 31087 38347 31093
rect 38654 31084 38660 31096
rect 38712 31084 38718 31136
rect 38746 31084 38752 31136
rect 38804 31124 38810 31136
rect 39301 31127 39359 31133
rect 39301 31124 39313 31127
rect 38804 31096 39313 31124
rect 38804 31084 38810 31096
rect 39301 31093 39313 31096
rect 39347 31124 39359 31127
rect 39853 31127 39911 31133
rect 39853 31124 39865 31127
rect 39347 31096 39865 31124
rect 39347 31093 39359 31096
rect 39301 31087 39359 31093
rect 39853 31093 39865 31096
rect 39899 31093 39911 31127
rect 39853 31087 39911 31093
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 13722 30880 13728 30932
rect 13780 30920 13786 30932
rect 14093 30923 14151 30929
rect 14093 30920 14105 30923
rect 13780 30892 14105 30920
rect 13780 30880 13786 30892
rect 14093 30889 14105 30892
rect 14139 30889 14151 30923
rect 15194 30920 15200 30932
rect 15155 30892 15200 30920
rect 14093 30883 14151 30889
rect 15194 30880 15200 30892
rect 15252 30880 15258 30932
rect 16577 30923 16635 30929
rect 16577 30889 16589 30923
rect 16623 30920 16635 30923
rect 16850 30920 16856 30932
rect 16623 30892 16856 30920
rect 16623 30889 16635 30892
rect 16577 30883 16635 30889
rect 16850 30880 16856 30892
rect 16908 30880 16914 30932
rect 17402 30920 17408 30932
rect 17363 30892 17408 30920
rect 17402 30880 17408 30892
rect 17460 30880 17466 30932
rect 18690 30920 18696 30932
rect 18651 30892 18696 30920
rect 18690 30880 18696 30892
rect 18748 30880 18754 30932
rect 19978 30920 19984 30932
rect 19939 30892 19984 30920
rect 19978 30880 19984 30892
rect 20036 30880 20042 30932
rect 20070 30880 20076 30932
rect 20128 30920 20134 30932
rect 20625 30923 20683 30929
rect 20625 30920 20637 30923
rect 20128 30892 20637 30920
rect 20128 30880 20134 30892
rect 20625 30889 20637 30892
rect 20671 30889 20683 30923
rect 20625 30883 20683 30889
rect 20809 30923 20867 30929
rect 20809 30889 20821 30923
rect 20855 30920 20867 30923
rect 20990 30920 20996 30932
rect 20855 30892 20996 30920
rect 20855 30889 20867 30892
rect 20809 30883 20867 30889
rect 20990 30880 20996 30892
rect 21048 30880 21054 30932
rect 21361 30923 21419 30929
rect 21361 30889 21373 30923
rect 21407 30920 21419 30923
rect 21450 30920 21456 30932
rect 21407 30892 21456 30920
rect 21407 30889 21419 30892
rect 21361 30883 21419 30889
rect 21450 30880 21456 30892
rect 21508 30880 21514 30932
rect 22370 30920 22376 30932
rect 22331 30892 22376 30920
rect 22370 30880 22376 30892
rect 22428 30880 22434 30932
rect 27525 30923 27583 30929
rect 27525 30889 27537 30923
rect 27571 30920 27583 30923
rect 27706 30920 27712 30932
rect 27571 30892 27712 30920
rect 27571 30889 27583 30892
rect 27525 30883 27583 30889
rect 27706 30880 27712 30892
rect 27764 30880 27770 30932
rect 29641 30923 29699 30929
rect 29641 30889 29653 30923
rect 29687 30920 29699 30923
rect 30006 30920 30012 30932
rect 29687 30892 30012 30920
rect 29687 30889 29699 30892
rect 29641 30883 29699 30889
rect 30006 30880 30012 30892
rect 30064 30880 30070 30932
rect 30742 30920 30748 30932
rect 30703 30892 30748 30920
rect 30742 30880 30748 30892
rect 30800 30880 30806 30932
rect 33134 30880 33140 30932
rect 33192 30920 33198 30932
rect 33505 30923 33563 30929
rect 33505 30920 33517 30923
rect 33192 30892 33517 30920
rect 33192 30880 33198 30892
rect 33505 30889 33517 30892
rect 33551 30889 33563 30923
rect 37090 30920 37096 30932
rect 37051 30892 37096 30920
rect 33505 30883 33563 30889
rect 37090 30880 37096 30892
rect 37148 30880 37154 30932
rect 38010 30880 38016 30932
rect 38068 30920 38074 30932
rect 38197 30923 38255 30929
rect 38197 30920 38209 30923
rect 38068 30892 38209 30920
rect 38068 30880 38074 30892
rect 38197 30889 38209 30892
rect 38243 30889 38255 30923
rect 38746 30920 38752 30932
rect 38707 30892 38752 30920
rect 38197 30883 38255 30889
rect 38746 30880 38752 30892
rect 38804 30880 38810 30932
rect 14461 30855 14519 30861
rect 14461 30821 14473 30855
rect 14507 30852 14519 30855
rect 15562 30852 15568 30864
rect 14507 30824 15568 30852
rect 14507 30821 14519 30824
rect 14461 30815 14519 30821
rect 15562 30812 15568 30824
rect 15620 30812 15626 30864
rect 16485 30855 16543 30861
rect 16485 30821 16497 30855
rect 16531 30852 16543 30855
rect 17310 30852 17316 30864
rect 16531 30824 17316 30852
rect 16531 30821 16543 30824
rect 16485 30815 16543 30821
rect 17310 30812 17316 30824
rect 17368 30812 17374 30864
rect 19794 30812 19800 30864
rect 19852 30852 19858 30864
rect 20438 30852 20444 30864
rect 19852 30824 20444 30852
rect 19852 30812 19858 30824
rect 20438 30812 20444 30824
rect 20496 30812 20502 30864
rect 20530 30812 20536 30864
rect 20588 30852 20594 30864
rect 20588 30824 22324 30852
rect 20588 30812 20594 30824
rect 11885 30787 11943 30793
rect 11885 30753 11897 30787
rect 11931 30784 11943 30787
rect 13081 30787 13139 30793
rect 11931 30756 12572 30784
rect 11931 30753 11943 30756
rect 11885 30747 11943 30753
rect 12544 30728 12572 30756
rect 13081 30753 13093 30787
rect 13127 30784 13139 30787
rect 14185 30787 14243 30793
rect 14185 30784 14197 30787
rect 13127 30756 14197 30784
rect 13127 30753 13139 30756
rect 13081 30747 13139 30753
rect 14185 30753 14197 30756
rect 14231 30784 14243 30787
rect 14826 30784 14832 30796
rect 14231 30756 14832 30784
rect 14231 30753 14243 30756
rect 14185 30747 14243 30753
rect 14826 30744 14832 30756
rect 14884 30784 14890 30796
rect 17494 30784 17500 30796
rect 14884 30756 15424 30784
rect 14884 30744 14890 30756
rect 11333 30719 11391 30725
rect 11333 30685 11345 30719
rect 11379 30716 11391 30719
rect 12342 30716 12348 30728
rect 11379 30688 12348 30716
rect 11379 30685 11391 30688
rect 11333 30679 11391 30685
rect 12342 30676 12348 30688
rect 12400 30676 12406 30728
rect 12526 30716 12532 30728
rect 12487 30688 12532 30716
rect 12526 30676 12532 30688
rect 12584 30676 12590 30728
rect 12986 30716 12992 30728
rect 12947 30688 12992 30716
rect 12986 30676 12992 30688
rect 13044 30676 13050 30728
rect 13173 30719 13231 30725
rect 13173 30685 13185 30719
rect 13219 30685 13231 30719
rect 13173 30679 13231 30685
rect 12437 30651 12495 30657
rect 12437 30617 12449 30651
rect 12483 30648 12495 30651
rect 13188 30648 13216 30679
rect 13262 30676 13268 30728
rect 13320 30716 13326 30728
rect 15396 30725 15424 30756
rect 17420 30756 17500 30784
rect 14093 30719 14151 30725
rect 14093 30716 14105 30719
rect 13320 30688 14105 30716
rect 13320 30676 13326 30688
rect 14093 30685 14105 30688
rect 14139 30685 14151 30719
rect 14093 30679 14151 30685
rect 15381 30719 15439 30725
rect 15381 30685 15393 30719
rect 15427 30685 15439 30719
rect 15657 30719 15715 30725
rect 15657 30716 15669 30719
rect 15381 30679 15439 30685
rect 15488 30688 15669 30716
rect 13814 30648 13820 30660
rect 12483 30620 13820 30648
rect 12483 30617 12495 30620
rect 12437 30611 12495 30617
rect 13814 30608 13820 30620
rect 13872 30608 13878 30660
rect 15286 30608 15292 30660
rect 15344 30648 15350 30660
rect 15488 30648 15516 30688
rect 15657 30685 15669 30688
rect 15703 30685 15715 30719
rect 15657 30679 15715 30685
rect 16850 30676 16856 30728
rect 16908 30716 16914 30728
rect 17420 30725 17448 30756
rect 17494 30744 17500 30756
rect 17552 30744 17558 30796
rect 21174 30744 21180 30796
rect 21232 30784 21238 30796
rect 22296 30793 22324 30824
rect 27246 30812 27252 30864
rect 27304 30852 27310 30864
rect 28353 30855 28411 30861
rect 28353 30852 28365 30855
rect 27304 30824 28365 30852
rect 27304 30812 27310 30824
rect 28353 30821 28365 30824
rect 28399 30821 28411 30855
rect 28353 30815 28411 30821
rect 21729 30787 21787 30793
rect 21729 30784 21741 30787
rect 21232 30756 21741 30784
rect 21232 30744 21238 30756
rect 21729 30753 21741 30756
rect 21775 30753 21787 30787
rect 21729 30747 21787 30753
rect 22281 30787 22339 30793
rect 22281 30753 22293 30787
rect 22327 30753 22339 30787
rect 22281 30747 22339 30753
rect 17405 30719 17463 30725
rect 17405 30716 17417 30719
rect 16908 30688 17417 30716
rect 16908 30676 16914 30688
rect 17405 30685 17417 30688
rect 17451 30685 17463 30719
rect 17405 30679 17463 30685
rect 17681 30719 17739 30725
rect 17681 30685 17693 30719
rect 17727 30716 17739 30719
rect 18046 30716 18052 30728
rect 17727 30688 18052 30716
rect 17727 30685 17739 30688
rect 17681 30679 17739 30685
rect 18046 30676 18052 30688
rect 18104 30676 18110 30728
rect 19426 30676 19432 30728
rect 19484 30716 19490 30728
rect 19705 30719 19763 30725
rect 19705 30716 19717 30719
rect 19484 30688 19717 30716
rect 19484 30676 19490 30688
rect 19705 30685 19717 30688
rect 19751 30716 19763 30719
rect 19751 30688 20576 30716
rect 19751 30685 19763 30688
rect 19705 30679 19763 30685
rect 15344 30620 15516 30648
rect 15565 30651 15623 30657
rect 15344 30608 15350 30620
rect 15565 30617 15577 30651
rect 15611 30648 15623 30651
rect 15838 30648 15844 30660
rect 15611 30620 15844 30648
rect 15611 30617 15623 30620
rect 15565 30611 15623 30617
rect 15838 30608 15844 30620
rect 15896 30608 15902 30660
rect 16022 30608 16028 30660
rect 16080 30648 16086 30660
rect 16117 30651 16175 30657
rect 16117 30648 16129 30651
rect 16080 30620 16129 30648
rect 16080 30608 16086 30620
rect 16117 30617 16129 30620
rect 16163 30617 16175 30651
rect 16117 30611 16175 30617
rect 17310 30608 17316 30660
rect 17368 30648 17374 30660
rect 17497 30651 17555 30657
rect 17497 30648 17509 30651
rect 17368 30620 17509 30648
rect 17368 30608 17374 30620
rect 17497 30617 17509 30620
rect 17543 30617 17555 30651
rect 17497 30611 17555 30617
rect 19981 30651 20039 30657
rect 19981 30617 19993 30651
rect 20027 30648 20039 30651
rect 20346 30648 20352 30660
rect 20027 30620 20352 30648
rect 20027 30617 20039 30620
rect 19981 30611 20039 30617
rect 20346 30608 20352 30620
rect 20404 30648 20410 30660
rect 20441 30651 20499 30657
rect 20441 30648 20453 30651
rect 20404 30620 20453 30648
rect 20404 30608 20410 30620
rect 20441 30617 20453 30620
rect 20487 30617 20499 30651
rect 20548 30648 20576 30688
rect 21266 30676 21272 30728
rect 21324 30716 21330 30728
rect 21637 30719 21695 30725
rect 21637 30716 21649 30719
rect 21324 30688 21649 30716
rect 21324 30676 21330 30688
rect 21637 30685 21649 30688
rect 21683 30685 21695 30719
rect 21744 30716 21772 30747
rect 24302 30744 24308 30796
rect 24360 30784 24366 30796
rect 32033 30787 32091 30793
rect 24360 30756 24624 30784
rect 24360 30744 24366 30756
rect 22465 30719 22523 30725
rect 22465 30716 22477 30719
rect 21744 30688 22477 30716
rect 21637 30679 21695 30685
rect 22465 30685 22477 30688
rect 22511 30685 22523 30719
rect 22465 30679 22523 30685
rect 22557 30719 22615 30725
rect 22557 30685 22569 30719
rect 22603 30685 22615 30719
rect 22557 30679 22615 30685
rect 20622 30648 20628 30660
rect 20680 30657 20686 30660
rect 20680 30651 20699 30657
rect 20548 30620 20628 30648
rect 20441 30611 20499 30617
rect 19797 30583 19855 30589
rect 19797 30549 19809 30583
rect 19843 30580 19855 30583
rect 20070 30580 20076 30592
rect 19843 30552 20076 30580
rect 19843 30549 19855 30552
rect 19797 30543 19855 30549
rect 20070 30540 20076 30552
rect 20128 30540 20134 30592
rect 20456 30580 20484 30611
rect 20622 30608 20628 30620
rect 20687 30648 20699 30651
rect 21652 30648 21680 30679
rect 22094 30648 22100 30660
rect 20687 30620 20773 30648
rect 21652 30620 22100 30648
rect 20687 30617 20699 30620
rect 20680 30611 20699 30617
rect 20680 30608 20686 30611
rect 22094 30608 22100 30620
rect 22152 30648 22158 30660
rect 22572 30648 22600 30679
rect 24118 30676 24124 30728
rect 24176 30716 24182 30728
rect 24397 30719 24455 30725
rect 24397 30716 24409 30719
rect 24176 30688 24409 30716
rect 24176 30676 24182 30688
rect 24397 30685 24409 30688
rect 24443 30716 24455 30719
rect 24486 30716 24492 30728
rect 24443 30688 24492 30716
rect 24443 30685 24455 30688
rect 24397 30679 24455 30685
rect 24486 30676 24492 30688
rect 24544 30676 24550 30728
rect 24596 30725 24624 30756
rect 32033 30753 32045 30787
rect 32079 30784 32091 30787
rect 32674 30784 32680 30796
rect 32079 30756 32680 30784
rect 32079 30753 32091 30756
rect 32033 30747 32091 30753
rect 32674 30744 32680 30756
rect 32732 30744 32738 30796
rect 33226 30744 33232 30796
rect 33284 30784 33290 30796
rect 36541 30787 36599 30793
rect 36541 30784 36553 30787
rect 33284 30756 36553 30784
rect 33284 30744 33290 30756
rect 36541 30753 36553 30756
rect 36587 30753 36599 30787
rect 36541 30747 36599 30753
rect 24581 30719 24639 30725
rect 24581 30685 24593 30719
rect 24627 30716 24639 30719
rect 25958 30716 25964 30728
rect 24627 30688 25964 30716
rect 24627 30685 24639 30688
rect 24581 30679 24639 30685
rect 25958 30676 25964 30688
rect 26016 30676 26022 30728
rect 26786 30716 26792 30728
rect 26747 30688 26792 30716
rect 26786 30676 26792 30688
rect 26844 30676 26850 30728
rect 29454 30676 29460 30728
rect 29512 30716 29518 30728
rect 29549 30719 29607 30725
rect 29549 30716 29561 30719
rect 29512 30688 29561 30716
rect 29512 30676 29518 30688
rect 29549 30685 29561 30688
rect 29595 30685 29607 30719
rect 29549 30679 29607 30685
rect 29733 30719 29791 30725
rect 29733 30685 29745 30719
rect 29779 30716 29791 30719
rect 30650 30716 30656 30728
rect 29779 30688 30656 30716
rect 29779 30685 29791 30688
rect 29733 30679 29791 30685
rect 22152 30620 22600 30648
rect 22152 30608 22158 30620
rect 27522 30608 27528 30660
rect 27580 30648 27586 30660
rect 27709 30651 27767 30657
rect 27709 30648 27721 30651
rect 27580 30620 27721 30648
rect 27580 30608 27586 30620
rect 27709 30617 27721 30620
rect 27755 30617 27767 30651
rect 27890 30648 27896 30660
rect 27851 30620 27896 30648
rect 27709 30611 27767 30617
rect 27890 30608 27896 30620
rect 27948 30608 27954 30660
rect 29270 30608 29276 30660
rect 29328 30648 29334 30660
rect 29748 30648 29776 30679
rect 30650 30676 30656 30688
rect 30708 30676 30714 30728
rect 31113 30719 31171 30725
rect 31113 30685 31125 30719
rect 31159 30716 31171 30719
rect 31386 30716 31392 30728
rect 31159 30688 31392 30716
rect 31159 30685 31171 30688
rect 31113 30679 31171 30685
rect 31386 30676 31392 30688
rect 31444 30716 31450 30728
rect 31444 30688 31754 30716
rect 31444 30676 31450 30688
rect 29328 30620 29776 30648
rect 30929 30651 30987 30657
rect 29328 30608 29334 30620
rect 30929 30617 30941 30651
rect 30975 30648 30987 30651
rect 31018 30648 31024 30660
rect 30975 30620 31024 30648
rect 30975 30617 30987 30620
rect 30929 30611 30987 30617
rect 20990 30580 20996 30592
rect 20456 30552 20996 30580
rect 20990 30540 20996 30552
rect 21048 30540 21054 30592
rect 21726 30540 21732 30592
rect 21784 30580 21790 30592
rect 23109 30583 23167 30589
rect 23109 30580 23121 30583
rect 21784 30552 23121 30580
rect 21784 30540 21790 30552
rect 23109 30549 23121 30552
rect 23155 30580 23167 30583
rect 23750 30580 23756 30592
rect 23155 30552 23756 30580
rect 23155 30549 23167 30552
rect 23109 30543 23167 30549
rect 23750 30540 23756 30552
rect 23808 30540 23814 30592
rect 24026 30540 24032 30592
rect 24084 30580 24090 30592
rect 24489 30583 24547 30589
rect 24489 30580 24501 30583
rect 24084 30552 24501 30580
rect 24084 30540 24090 30552
rect 24489 30549 24501 30552
rect 24535 30580 24547 30583
rect 24762 30580 24768 30592
rect 24535 30552 24768 30580
rect 24535 30549 24547 30552
rect 24489 30543 24547 30549
rect 24762 30540 24768 30552
rect 24820 30540 24826 30592
rect 24854 30540 24860 30592
rect 24912 30580 24918 30592
rect 25133 30583 25191 30589
rect 25133 30580 25145 30583
rect 24912 30552 25145 30580
rect 24912 30540 24918 30552
rect 25133 30549 25145 30552
rect 25179 30549 25191 30583
rect 25133 30543 25191 30549
rect 26053 30583 26111 30589
rect 26053 30549 26065 30583
rect 26099 30580 26111 30583
rect 26234 30580 26240 30592
rect 26099 30552 26240 30580
rect 26099 30549 26111 30552
rect 26053 30543 26111 30549
rect 26234 30540 26240 30552
rect 26292 30580 26298 30592
rect 26510 30580 26516 30592
rect 26292 30552 26516 30580
rect 26292 30540 26298 30552
rect 26510 30540 26516 30552
rect 26568 30540 26574 30592
rect 26881 30583 26939 30589
rect 26881 30549 26893 30583
rect 26927 30580 26939 30583
rect 26970 30580 26976 30592
rect 26927 30552 26976 30580
rect 26927 30549 26939 30552
rect 26881 30543 26939 30549
rect 26970 30540 26976 30552
rect 27028 30540 27034 30592
rect 28994 30580 29000 30592
rect 28955 30552 29000 30580
rect 28994 30540 29000 30552
rect 29052 30580 29058 30592
rect 29178 30580 29184 30592
rect 29052 30552 29184 30580
rect 29052 30540 29058 30552
rect 29178 30540 29184 30552
rect 29236 30540 29242 30592
rect 29546 30540 29552 30592
rect 29604 30580 29610 30592
rect 30098 30580 30104 30592
rect 29604 30552 30104 30580
rect 29604 30540 29610 30552
rect 30098 30540 30104 30552
rect 30156 30580 30162 30592
rect 30193 30583 30251 30589
rect 30193 30580 30205 30583
rect 30156 30552 30205 30580
rect 30156 30540 30162 30552
rect 30193 30549 30205 30552
rect 30239 30549 30251 30583
rect 30944 30580 30972 30611
rect 31018 30608 31024 30620
rect 31076 30608 31082 30660
rect 31726 30648 31754 30688
rect 32214 30676 32220 30728
rect 32272 30716 32278 30728
rect 32272 30688 32338 30716
rect 32272 30676 32278 30688
rect 32950 30676 32956 30728
rect 33008 30716 33014 30728
rect 33502 30716 33508 30728
rect 33008 30688 33053 30716
rect 33463 30688 33508 30716
rect 33008 30676 33014 30688
rect 33502 30676 33508 30688
rect 33560 30676 33566 30728
rect 33689 30719 33747 30725
rect 33689 30685 33701 30719
rect 33735 30685 33747 30719
rect 36446 30716 36452 30728
rect 33689 30679 33747 30685
rect 35176 30688 36452 30716
rect 32030 30648 32036 30660
rect 31726 30620 32036 30648
rect 32030 30608 32036 30620
rect 32088 30608 32094 30660
rect 32490 30608 32496 30660
rect 32548 30648 32554 30660
rect 33704 30648 33732 30679
rect 32548 30620 33732 30648
rect 32548 30608 32554 30620
rect 34698 30608 34704 30660
rect 34756 30648 34762 30660
rect 35176 30657 35204 30688
rect 36446 30676 36452 30688
rect 36504 30716 36510 30728
rect 37645 30719 37703 30725
rect 37645 30716 37657 30719
rect 36504 30688 37657 30716
rect 36504 30676 36510 30688
rect 37645 30685 37657 30688
rect 37691 30685 37703 30719
rect 37645 30679 37703 30685
rect 35161 30651 35219 30657
rect 35161 30648 35173 30651
rect 34756 30620 35173 30648
rect 34756 30608 34762 30620
rect 35161 30617 35173 30620
rect 35207 30617 35219 30651
rect 35161 30611 35219 30617
rect 35345 30651 35403 30657
rect 35345 30617 35357 30651
rect 35391 30648 35403 30651
rect 37090 30648 37096 30660
rect 35391 30620 37096 30648
rect 35391 30617 35403 30620
rect 35345 30611 35403 30617
rect 33226 30580 33232 30592
rect 30944 30552 33232 30580
rect 30193 30543 30251 30549
rect 33226 30540 33232 30552
rect 33284 30540 33290 30592
rect 34054 30540 34060 30592
rect 34112 30580 34118 30592
rect 35360 30580 35388 30611
rect 37090 30608 37096 30620
rect 37148 30608 37154 30660
rect 34112 30552 35388 30580
rect 35529 30583 35587 30589
rect 34112 30540 34118 30552
rect 35529 30549 35541 30583
rect 35575 30580 35587 30583
rect 35894 30580 35900 30592
rect 35575 30552 35900 30580
rect 35575 30549 35587 30552
rect 35529 30543 35587 30549
rect 35894 30540 35900 30552
rect 35952 30540 35958 30592
rect 35986 30540 35992 30592
rect 36044 30580 36050 30592
rect 36044 30552 36089 30580
rect 36044 30540 36050 30552
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 12069 30379 12127 30385
rect 12069 30345 12081 30379
rect 12115 30376 12127 30379
rect 12342 30376 12348 30388
rect 12115 30348 12348 30376
rect 12115 30345 12127 30348
rect 12069 30339 12127 30345
rect 12342 30336 12348 30348
rect 12400 30336 12406 30388
rect 12526 30376 12532 30388
rect 12487 30348 12532 30376
rect 12526 30336 12532 30348
rect 12584 30336 12590 30388
rect 13725 30379 13783 30385
rect 13725 30345 13737 30379
rect 13771 30376 13783 30379
rect 15378 30376 15384 30388
rect 13771 30348 15384 30376
rect 13771 30345 13783 30348
rect 13725 30339 13783 30345
rect 15378 30336 15384 30348
rect 15436 30376 15442 30388
rect 15838 30376 15844 30388
rect 15436 30348 15844 30376
rect 15436 30336 15442 30348
rect 15838 30336 15844 30348
rect 15896 30336 15902 30388
rect 17129 30379 17187 30385
rect 17129 30345 17141 30379
rect 17175 30376 17187 30379
rect 17310 30376 17316 30388
rect 17175 30348 17316 30376
rect 17175 30345 17187 30348
rect 17129 30339 17187 30345
rect 17310 30336 17316 30348
rect 17368 30336 17374 30388
rect 18046 30376 18052 30388
rect 17604 30348 18052 30376
rect 17604 30317 17632 30348
rect 18046 30336 18052 30348
rect 18104 30336 18110 30388
rect 19426 30336 19432 30388
rect 19484 30376 19490 30388
rect 19613 30379 19671 30385
rect 19613 30376 19625 30379
rect 19484 30348 19625 30376
rect 19484 30336 19490 30348
rect 19613 30345 19625 30348
rect 19659 30345 19671 30379
rect 19613 30339 19671 30345
rect 20530 30336 20536 30388
rect 20588 30376 20594 30388
rect 20625 30379 20683 30385
rect 20625 30376 20637 30379
rect 20588 30348 20637 30376
rect 20588 30336 20594 30348
rect 20625 30345 20637 30348
rect 20671 30345 20683 30379
rect 22278 30376 22284 30388
rect 20625 30339 20683 30345
rect 21008 30348 21312 30376
rect 22239 30348 22284 30376
rect 2041 30311 2099 30317
rect 2041 30277 2053 30311
rect 2087 30308 2099 30311
rect 17589 30311 17647 30317
rect 2087 30280 16896 30308
rect 2087 30277 2099 30280
rect 2041 30271 2099 30277
rect 1578 30200 1584 30252
rect 1636 30240 1642 30252
rect 1857 30243 1915 30249
rect 1857 30240 1869 30243
rect 1636 30212 1869 30240
rect 1636 30200 1642 30212
rect 1857 30209 1869 30212
rect 1903 30209 1915 30243
rect 13170 30240 13176 30252
rect 13131 30212 13176 30240
rect 1857 30203 1915 30209
rect 13170 30200 13176 30212
rect 13228 30200 13234 30252
rect 14277 30243 14335 30249
rect 14277 30209 14289 30243
rect 14323 30240 14335 30243
rect 15286 30240 15292 30252
rect 14323 30212 15292 30240
rect 14323 30209 14335 30212
rect 14277 30203 14335 30209
rect 15286 30200 15292 30212
rect 15344 30200 15350 30252
rect 15562 30240 15568 30252
rect 15523 30212 15568 30240
rect 15562 30200 15568 30212
rect 15620 30200 15626 30252
rect 16298 30200 16304 30252
rect 16356 30240 16362 30252
rect 16666 30240 16672 30252
rect 16356 30212 16672 30240
rect 16356 30200 16362 30212
rect 16666 30200 16672 30212
rect 16724 30200 16730 30252
rect 16761 30243 16819 30249
rect 16761 30209 16773 30243
rect 16807 30209 16819 30243
rect 16761 30203 16819 30209
rect 15749 30175 15807 30181
rect 15749 30141 15761 30175
rect 15795 30172 15807 30175
rect 16574 30172 16580 30184
rect 15795 30144 16580 30172
rect 15795 30141 15807 30144
rect 15749 30135 15807 30141
rect 16574 30132 16580 30144
rect 16632 30172 16638 30184
rect 16776 30172 16804 30203
rect 16632 30144 16804 30172
rect 16868 30172 16896 30280
rect 17589 30277 17601 30311
rect 17635 30277 17647 30311
rect 21008 30308 21036 30348
rect 21174 30317 21180 30320
rect 17589 30271 17647 30277
rect 17880 30280 21036 30308
rect 21131 30311 21180 30317
rect 16942 30200 16948 30252
rect 17000 30240 17006 30252
rect 17773 30243 17831 30249
rect 17773 30240 17785 30243
rect 17000 30212 17785 30240
rect 17000 30200 17006 30212
rect 17773 30209 17785 30212
rect 17819 30209 17831 30243
rect 17773 30203 17831 30209
rect 17880 30172 17908 30280
rect 21131 30277 21143 30311
rect 21177 30277 21180 30311
rect 21131 30271 21180 30277
rect 21174 30268 21180 30271
rect 21232 30268 21238 30320
rect 21284 30308 21312 30348
rect 22278 30336 22284 30348
rect 22336 30336 22342 30388
rect 24762 30336 24768 30388
rect 24820 30376 24826 30388
rect 24949 30379 25007 30385
rect 24949 30376 24961 30379
rect 24820 30348 24961 30376
rect 24820 30336 24826 30348
rect 24949 30345 24961 30348
rect 24995 30345 25007 30379
rect 24949 30339 25007 30345
rect 27356 30348 27936 30376
rect 27356 30308 27384 30348
rect 21284 30280 27384 30308
rect 27430 30268 27436 30320
rect 27488 30308 27494 30320
rect 27801 30311 27859 30317
rect 27801 30308 27813 30311
rect 27488 30280 27813 30308
rect 27488 30268 27494 30280
rect 27801 30277 27813 30280
rect 27847 30277 27859 30311
rect 27908 30308 27936 30348
rect 29086 30336 29092 30388
rect 29144 30376 29150 30388
rect 32309 30379 32367 30385
rect 29144 30348 31340 30376
rect 29144 30336 29150 30348
rect 27908 30280 28672 30308
rect 27801 30271 27859 30277
rect 18877 30243 18935 30249
rect 18877 30209 18889 30243
rect 18923 30209 18935 30243
rect 18877 30203 18935 30209
rect 19061 30243 19119 30249
rect 19061 30209 19073 30243
rect 19107 30240 19119 30243
rect 19242 30240 19248 30252
rect 19107 30212 19248 30240
rect 19107 30209 19119 30212
rect 19061 30203 19119 30209
rect 16868 30144 17908 30172
rect 16632 30132 16638 30144
rect 18892 30104 18920 30203
rect 19242 30200 19248 30212
rect 19300 30200 19306 30252
rect 19518 30240 19524 30252
rect 19479 30212 19524 30240
rect 19518 30200 19524 30212
rect 19576 30200 19582 30252
rect 19705 30243 19763 30249
rect 19705 30209 19717 30243
rect 19751 30209 19763 30243
rect 19705 30203 19763 30209
rect 19797 30243 19855 30249
rect 19797 30209 19809 30243
rect 19843 30209 19855 30243
rect 19797 30203 19855 30209
rect 19334 30132 19340 30184
rect 19392 30172 19398 30184
rect 19720 30172 19748 30203
rect 19392 30144 19748 30172
rect 19392 30132 19398 30144
rect 17788 30076 18920 30104
rect 17788 30048 17816 30076
rect 14829 30039 14887 30045
rect 14829 30005 14841 30039
rect 14875 30036 14887 30039
rect 17770 30036 17776 30048
rect 14875 30008 17776 30036
rect 14875 30005 14887 30008
rect 14829 29999 14887 30005
rect 17770 29996 17776 30008
rect 17828 29996 17834 30048
rect 17954 30036 17960 30048
rect 17915 30008 17960 30036
rect 17954 29996 17960 30008
rect 18012 29996 18018 30048
rect 18892 30036 18920 30076
rect 18969 30107 19027 30113
rect 18969 30073 18981 30107
rect 19015 30104 19027 30107
rect 19426 30104 19432 30116
rect 19015 30076 19432 30104
rect 19015 30073 19027 30076
rect 18969 30067 19027 30073
rect 19426 30064 19432 30076
rect 19484 30104 19490 30116
rect 19812 30104 19840 30203
rect 20622 30200 20628 30252
rect 20680 30240 20686 30252
rect 20809 30243 20867 30249
rect 20809 30240 20821 30243
rect 20680 30212 20821 30240
rect 20680 30200 20686 30212
rect 20809 30209 20821 30212
rect 20855 30209 20867 30243
rect 20809 30203 20867 30209
rect 20901 30243 20959 30249
rect 20901 30209 20913 30243
rect 20947 30209 20959 30243
rect 20901 30203 20959 30209
rect 20070 30132 20076 30184
rect 20128 30172 20134 30184
rect 20916 30172 20944 30203
rect 20990 30200 20996 30252
rect 21048 30240 21054 30252
rect 21048 30212 21093 30240
rect 21048 30200 21054 30212
rect 21266 30200 21272 30252
rect 21324 30240 21330 30252
rect 23014 30240 23020 30252
rect 21324 30212 21369 30240
rect 22975 30212 23020 30240
rect 21324 30200 21330 30212
rect 23014 30200 23020 30212
rect 23072 30200 23078 30252
rect 24026 30240 24032 30252
rect 23987 30212 24032 30240
rect 24026 30200 24032 30212
rect 24084 30200 24090 30252
rect 24857 30243 24915 30249
rect 24857 30240 24869 30243
rect 24228 30212 24869 30240
rect 23934 30172 23940 30184
rect 20128 30144 20944 30172
rect 23895 30144 23940 30172
rect 20128 30132 20134 30144
rect 23934 30132 23940 30144
rect 23992 30172 23998 30184
rect 24228 30172 24256 30212
rect 24857 30209 24869 30212
rect 24903 30209 24915 30243
rect 25130 30240 25136 30252
rect 25091 30212 25136 30240
rect 24857 30203 24915 30209
rect 24394 30172 24400 30184
rect 23992 30144 24256 30172
rect 24355 30144 24400 30172
rect 23992 30132 23998 30144
rect 24394 30132 24400 30144
rect 24452 30132 24458 30184
rect 24872 30172 24900 30203
rect 25130 30200 25136 30212
rect 25188 30200 25194 30252
rect 25774 30240 25780 30252
rect 25735 30212 25780 30240
rect 25774 30200 25780 30212
rect 25832 30200 25838 30252
rect 25961 30243 26019 30249
rect 25961 30209 25973 30243
rect 26007 30209 26019 30243
rect 25961 30203 26019 30209
rect 25976 30172 26004 30203
rect 26878 30200 26884 30252
rect 26936 30240 26942 30252
rect 27525 30243 27583 30249
rect 27525 30240 27537 30243
rect 26936 30212 27537 30240
rect 26936 30200 26942 30212
rect 27525 30209 27537 30212
rect 27571 30209 27583 30243
rect 28261 30243 28319 30249
rect 28261 30240 28273 30243
rect 27525 30203 27583 30209
rect 27632 30212 28273 30240
rect 24872 30144 26004 30172
rect 19484 30076 19840 30104
rect 25869 30107 25927 30113
rect 19484 30064 19490 30076
rect 25869 30073 25881 30107
rect 25915 30104 25927 30107
rect 26786 30104 26792 30116
rect 25915 30076 26792 30104
rect 25915 30073 25927 30076
rect 25869 30067 25927 30073
rect 26786 30064 26792 30076
rect 26844 30064 26850 30116
rect 27632 30048 27660 30212
rect 28261 30209 28273 30212
rect 28307 30209 28319 30243
rect 28261 30203 28319 30209
rect 28350 30200 28356 30252
rect 28408 30240 28414 30252
rect 28534 30240 28540 30252
rect 28408 30212 28453 30240
rect 28495 30212 28540 30240
rect 28408 30200 28414 30212
rect 28534 30200 28540 30212
rect 28592 30200 28598 30252
rect 27801 30175 27859 30181
rect 27801 30141 27813 30175
rect 27847 30141 27859 30175
rect 27801 30135 27859 30141
rect 27816 30104 27844 30135
rect 28537 30107 28595 30113
rect 28537 30104 28549 30107
rect 27816 30076 28549 30104
rect 28537 30073 28549 30076
rect 28583 30073 28595 30107
rect 28644 30104 28672 30280
rect 28810 30268 28816 30320
rect 28868 30308 28874 30320
rect 31312 30308 31340 30348
rect 32309 30345 32321 30379
rect 32355 30376 32367 30379
rect 32677 30379 32735 30385
rect 32355 30348 32628 30376
rect 32355 30345 32367 30348
rect 32309 30339 32367 30345
rect 31573 30311 31631 30317
rect 28868 30280 31248 30308
rect 31312 30280 31524 30308
rect 28868 30268 28874 30280
rect 29086 30240 29092 30252
rect 29047 30212 29092 30240
rect 29086 30200 29092 30212
rect 29144 30200 29150 30252
rect 29638 30200 29644 30252
rect 29696 30240 29702 30252
rect 29825 30243 29883 30249
rect 29825 30240 29837 30243
rect 29696 30212 29837 30240
rect 29696 30200 29702 30212
rect 29825 30209 29837 30212
rect 29871 30209 29883 30243
rect 29825 30203 29883 30209
rect 29914 30200 29920 30252
rect 29972 30240 29978 30252
rect 30285 30243 30343 30249
rect 30285 30240 30297 30243
rect 29972 30212 30297 30240
rect 29972 30200 29978 30212
rect 30285 30209 30297 30212
rect 30331 30209 30343 30243
rect 30285 30203 30343 30209
rect 30469 30243 30527 30249
rect 30469 30209 30481 30243
rect 30515 30209 30527 30243
rect 30469 30203 30527 30209
rect 29546 30172 29552 30184
rect 29507 30144 29552 30172
rect 29546 30132 29552 30144
rect 29604 30132 29610 30184
rect 30190 30132 30196 30184
rect 30248 30172 30254 30184
rect 30484 30172 30512 30203
rect 31220 30181 31248 30280
rect 31386 30240 31392 30252
rect 31347 30212 31392 30240
rect 31386 30200 31392 30212
rect 31444 30200 31450 30252
rect 31496 30240 31524 30280
rect 31573 30277 31585 30311
rect 31619 30308 31631 30311
rect 32600 30308 32628 30348
rect 32677 30345 32689 30379
rect 32723 30376 32735 30379
rect 32766 30376 32772 30388
rect 32723 30348 32772 30376
rect 32723 30345 32735 30348
rect 32677 30339 32735 30345
rect 32766 30336 32772 30348
rect 32824 30336 32830 30388
rect 35253 30379 35311 30385
rect 35253 30345 35265 30379
rect 35299 30376 35311 30379
rect 35710 30376 35716 30388
rect 35299 30348 35716 30376
rect 35299 30345 35311 30348
rect 35253 30339 35311 30345
rect 35710 30336 35716 30348
rect 35768 30336 35774 30388
rect 37090 30336 37096 30388
rect 37148 30376 37154 30388
rect 37277 30379 37335 30385
rect 37277 30376 37289 30379
rect 37148 30348 37289 30376
rect 37148 30336 37154 30348
rect 37277 30345 37289 30348
rect 37323 30345 37335 30379
rect 37277 30339 37335 30345
rect 38654 30336 38660 30388
rect 38712 30376 38718 30388
rect 39390 30376 39396 30388
rect 38712 30348 39396 30376
rect 38712 30336 38718 30348
rect 39390 30336 39396 30348
rect 39448 30336 39454 30388
rect 32950 30308 32956 30320
rect 31619 30280 32536 30308
rect 32600 30280 32956 30308
rect 31619 30277 31631 30280
rect 31573 30271 31631 30277
rect 32508 30252 32536 30280
rect 32950 30268 32956 30280
rect 33008 30268 33014 30320
rect 33505 30311 33563 30317
rect 33505 30277 33517 30311
rect 33551 30308 33563 30311
rect 33551 30280 34928 30308
rect 33551 30277 33563 30280
rect 33505 30271 33563 30277
rect 32214 30240 32220 30252
rect 31496 30212 31754 30240
rect 32175 30212 32220 30240
rect 30248 30144 30512 30172
rect 31205 30175 31263 30181
rect 30248 30132 30254 30144
rect 31205 30141 31217 30175
rect 31251 30172 31263 30175
rect 31478 30172 31484 30184
rect 31251 30144 31484 30172
rect 31251 30141 31263 30144
rect 31205 30135 31263 30141
rect 31478 30132 31484 30144
rect 31536 30132 31542 30184
rect 31726 30172 31754 30212
rect 32214 30200 32220 30212
rect 32272 30200 32278 30252
rect 32490 30240 32496 30252
rect 32451 30212 32496 30240
rect 32490 30200 32496 30212
rect 32548 30200 32554 30252
rect 33134 30200 33140 30252
rect 33192 30240 33198 30252
rect 33413 30243 33471 30249
rect 33413 30240 33425 30243
rect 33192 30212 33425 30240
rect 33192 30200 33198 30212
rect 33413 30209 33425 30212
rect 33459 30209 33471 30243
rect 33594 30240 33600 30252
rect 33555 30212 33600 30240
rect 33413 30203 33471 30209
rect 33594 30200 33600 30212
rect 33652 30200 33658 30252
rect 34054 30200 34060 30252
rect 34112 30240 34118 30252
rect 34241 30243 34299 30249
rect 34112 30212 34157 30240
rect 34112 30200 34118 30212
rect 34241 30209 34253 30243
rect 34287 30240 34299 30243
rect 34698 30240 34704 30252
rect 34287 30212 34704 30240
rect 34287 30209 34299 30212
rect 34241 30203 34299 30209
rect 34146 30172 34152 30184
rect 31726 30144 34152 30172
rect 34146 30132 34152 30144
rect 34204 30132 34210 30184
rect 34256 30104 34284 30203
rect 34698 30200 34704 30212
rect 34756 30200 34762 30252
rect 34900 30249 34928 30280
rect 34885 30243 34943 30249
rect 34885 30209 34897 30243
rect 34931 30240 34943 30243
rect 35250 30240 35256 30252
rect 34931 30212 35256 30240
rect 34931 30209 34943 30212
rect 34885 30203 34943 30209
rect 35250 30200 35256 30212
rect 35308 30200 35314 30252
rect 36357 30243 36415 30249
rect 36357 30209 36369 30243
rect 36403 30240 36415 30243
rect 36538 30240 36544 30252
rect 36403 30212 36544 30240
rect 36403 30209 36415 30212
rect 36357 30203 36415 30209
rect 36538 30200 36544 30212
rect 36596 30200 36602 30252
rect 37274 30240 37280 30252
rect 36648 30212 37280 30240
rect 34790 30172 34796 30184
rect 34751 30144 34796 30172
rect 34790 30132 34796 30144
rect 34848 30132 34854 30184
rect 36449 30175 36507 30181
rect 36449 30141 36461 30175
rect 36495 30172 36507 30175
rect 36648 30172 36676 30212
rect 37274 30200 37280 30212
rect 37332 30200 37338 30252
rect 36495 30144 36676 30172
rect 36725 30175 36783 30181
rect 36495 30141 36507 30144
rect 36449 30135 36507 30141
rect 36725 30141 36737 30175
rect 36771 30172 36783 30175
rect 39482 30172 39488 30184
rect 36771 30144 39488 30172
rect 36771 30141 36783 30144
rect 36725 30135 36783 30141
rect 39482 30132 39488 30144
rect 39540 30132 39546 30184
rect 28644 30076 34284 30104
rect 28537 30067 28595 30073
rect 20622 30036 20628 30048
rect 18892 30008 20628 30036
rect 20622 29996 20628 30008
rect 20680 29996 20686 30048
rect 25222 29996 25228 30048
rect 25280 30036 25286 30048
rect 25317 30039 25375 30045
rect 25317 30036 25329 30039
rect 25280 30008 25329 30036
rect 25280 29996 25286 30008
rect 25317 30005 25329 30008
rect 25363 30005 25375 30039
rect 25317 29999 25375 30005
rect 26234 29996 26240 30048
rect 26292 30036 26298 30048
rect 26973 30039 27031 30045
rect 26973 30036 26985 30039
rect 26292 30008 26985 30036
rect 26292 29996 26298 30008
rect 26973 30005 26985 30008
rect 27019 30036 27031 30039
rect 27062 30036 27068 30048
rect 27019 30008 27068 30036
rect 27019 30005 27031 30008
rect 26973 29999 27031 30005
rect 27062 29996 27068 30008
rect 27120 29996 27126 30048
rect 27614 30036 27620 30048
rect 27575 30008 27620 30036
rect 27614 29996 27620 30008
rect 27672 29996 27678 30048
rect 27798 29996 27804 30048
rect 27856 30036 27862 30048
rect 28810 30036 28816 30048
rect 27856 30008 28816 30036
rect 27856 29996 27862 30008
rect 28810 29996 28816 30008
rect 28868 29996 28874 30048
rect 29546 29996 29552 30048
rect 29604 30036 29610 30048
rect 29641 30039 29699 30045
rect 29641 30036 29653 30039
rect 29604 30008 29653 30036
rect 29604 29996 29610 30008
rect 29641 30005 29653 30008
rect 29687 30005 29699 30039
rect 29641 29999 29699 30005
rect 29733 30039 29791 30045
rect 29733 30005 29745 30039
rect 29779 30036 29791 30039
rect 29822 30036 29828 30048
rect 29779 30008 29828 30036
rect 29779 30005 29791 30008
rect 29733 29999 29791 30005
rect 29822 29996 29828 30008
rect 29880 30036 29886 30048
rect 30285 30039 30343 30045
rect 30285 30036 30297 30039
rect 29880 30008 30297 30036
rect 29880 29996 29886 30008
rect 30285 30005 30297 30008
rect 30331 30005 30343 30039
rect 30285 29999 30343 30005
rect 31478 29996 31484 30048
rect 31536 30036 31542 30048
rect 33318 30036 33324 30048
rect 31536 30008 33324 30036
rect 31536 29996 31542 30008
rect 33318 29996 33324 30008
rect 33376 29996 33382 30048
rect 33686 29996 33692 30048
rect 33744 30036 33750 30048
rect 34149 30039 34207 30045
rect 34149 30036 34161 30039
rect 33744 30008 34161 30036
rect 33744 29996 33750 30008
rect 34149 30005 34161 30008
rect 34195 30005 34207 30039
rect 34149 29999 34207 30005
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 1578 29832 1584 29844
rect 1539 29804 1584 29832
rect 1578 29792 1584 29804
rect 1636 29792 1642 29844
rect 15013 29835 15071 29841
rect 15013 29801 15025 29835
rect 15059 29832 15071 29835
rect 15378 29832 15384 29844
rect 15059 29804 15384 29832
rect 15059 29801 15071 29804
rect 15013 29795 15071 29801
rect 15378 29792 15384 29804
rect 15436 29792 15442 29844
rect 16022 29832 16028 29844
rect 15983 29804 16028 29832
rect 16022 29792 16028 29804
rect 16080 29792 16086 29844
rect 16209 29835 16267 29841
rect 16209 29801 16221 29835
rect 16255 29801 16267 29835
rect 16942 29832 16948 29844
rect 16903 29804 16948 29832
rect 16209 29795 16267 29801
rect 14461 29767 14519 29773
rect 14461 29733 14473 29767
rect 14507 29764 14519 29767
rect 15286 29764 15292 29776
rect 14507 29736 15292 29764
rect 14507 29733 14519 29736
rect 14461 29727 14519 29733
rect 15286 29724 15292 29736
rect 15344 29724 15350 29776
rect 16224 29764 16252 29795
rect 16942 29792 16948 29804
rect 17000 29792 17006 29844
rect 17770 29832 17776 29844
rect 17731 29804 17776 29832
rect 17770 29792 17776 29804
rect 17828 29792 17834 29844
rect 18509 29835 18567 29841
rect 18509 29801 18521 29835
rect 18555 29801 18567 29835
rect 18509 29795 18567 29801
rect 18693 29835 18751 29841
rect 18693 29801 18705 29835
rect 18739 29832 18751 29835
rect 18966 29832 18972 29844
rect 18739 29804 18972 29832
rect 18739 29801 18751 29804
rect 18693 29795 18751 29801
rect 16298 29764 16304 29776
rect 16224 29736 16304 29764
rect 16298 29724 16304 29736
rect 16356 29724 16362 29776
rect 16960 29764 16988 29792
rect 16408 29736 16988 29764
rect 18524 29764 18552 29795
rect 18966 29792 18972 29804
rect 19024 29792 19030 29844
rect 19797 29835 19855 29841
rect 19797 29801 19809 29835
rect 19843 29832 19855 29835
rect 20070 29832 20076 29844
rect 19843 29804 20076 29832
rect 19843 29801 19855 29804
rect 19797 29795 19855 29801
rect 20070 29792 20076 29804
rect 20128 29792 20134 29844
rect 21174 29832 21180 29844
rect 21135 29804 21180 29832
rect 21174 29792 21180 29804
rect 21232 29792 21238 29844
rect 22830 29832 22836 29844
rect 22791 29804 22836 29832
rect 22830 29792 22836 29804
rect 22888 29792 22894 29844
rect 23017 29835 23075 29841
rect 23017 29801 23029 29835
rect 23063 29832 23075 29835
rect 25130 29832 25136 29844
rect 23063 29804 25136 29832
rect 23063 29801 23075 29804
rect 23017 29795 23075 29801
rect 25130 29792 25136 29804
rect 25188 29792 25194 29844
rect 25240 29804 26004 29832
rect 19334 29764 19340 29776
rect 18524 29736 19340 29764
rect 16408 29628 16436 29736
rect 19334 29724 19340 29736
rect 19392 29724 19398 29776
rect 25240 29764 25268 29804
rect 20456 29736 25268 29764
rect 25501 29767 25559 29773
rect 16482 29656 16488 29708
rect 16540 29696 16546 29708
rect 20456 29696 20484 29736
rect 25501 29733 25513 29767
rect 25547 29764 25559 29767
rect 25866 29764 25872 29776
rect 25547 29736 25872 29764
rect 25547 29733 25559 29736
rect 25501 29727 25559 29733
rect 25866 29724 25872 29736
rect 25924 29724 25930 29776
rect 25976 29764 26004 29804
rect 26786 29792 26792 29844
rect 26844 29832 26850 29844
rect 26881 29835 26939 29841
rect 26881 29832 26893 29835
rect 26844 29804 26893 29832
rect 26844 29792 26850 29804
rect 26881 29801 26893 29804
rect 26927 29801 26939 29835
rect 26881 29795 26939 29801
rect 27709 29835 27767 29841
rect 27709 29801 27721 29835
rect 27755 29832 27767 29835
rect 27890 29832 27896 29844
rect 27755 29804 27896 29832
rect 27755 29801 27767 29804
rect 27709 29795 27767 29801
rect 27890 29792 27896 29804
rect 27948 29792 27954 29844
rect 28902 29832 28908 29844
rect 28863 29804 28908 29832
rect 28902 29792 28908 29804
rect 28960 29792 28966 29844
rect 29549 29835 29607 29841
rect 29549 29801 29561 29835
rect 29595 29832 29607 29835
rect 29730 29832 29736 29844
rect 29595 29804 29736 29832
rect 29595 29801 29607 29804
rect 29549 29795 29607 29801
rect 29730 29792 29736 29804
rect 29788 29792 29794 29844
rect 30466 29832 30472 29844
rect 30427 29804 30472 29832
rect 30466 29792 30472 29804
rect 30524 29792 30530 29844
rect 30558 29792 30564 29844
rect 30616 29832 30622 29844
rect 30653 29835 30711 29841
rect 30653 29832 30665 29835
rect 30616 29804 30665 29832
rect 30616 29792 30622 29804
rect 30653 29801 30665 29804
rect 30699 29801 30711 29835
rect 30653 29795 30711 29801
rect 31297 29835 31355 29841
rect 31297 29801 31309 29835
rect 31343 29832 31355 29835
rect 33502 29832 33508 29844
rect 31343 29804 33508 29832
rect 31343 29801 31355 29804
rect 31297 29795 31355 29801
rect 33502 29792 33508 29804
rect 33560 29792 33566 29844
rect 34149 29835 34207 29841
rect 34149 29801 34161 29835
rect 34195 29832 34207 29835
rect 34238 29832 34244 29844
rect 34195 29804 34244 29832
rect 34195 29801 34207 29804
rect 34149 29795 34207 29801
rect 34238 29792 34244 29804
rect 34296 29792 34302 29844
rect 34793 29835 34851 29841
rect 34793 29801 34805 29835
rect 34839 29832 34851 29835
rect 35986 29832 35992 29844
rect 34839 29804 35992 29832
rect 34839 29801 34851 29804
rect 34793 29795 34851 29801
rect 31386 29764 31392 29776
rect 25976 29736 31392 29764
rect 16540 29668 20484 29696
rect 16540 29656 16546 29668
rect 20530 29656 20536 29708
rect 20588 29696 20594 29708
rect 22278 29696 22284 29708
rect 20588 29668 22284 29696
rect 20588 29656 20594 29668
rect 16850 29628 16856 29640
rect 16208 29603 16436 29628
rect 16163 29600 16436 29603
rect 16811 29600 16856 29628
rect 16163 29597 16236 29600
rect 16163 29563 16175 29597
rect 16209 29566 16236 29597
rect 16850 29588 16856 29600
rect 16908 29588 16914 29640
rect 17034 29628 17040 29640
rect 16995 29600 17040 29628
rect 17034 29588 17040 29600
rect 17092 29588 17098 29640
rect 18598 29588 18604 29640
rect 18656 29588 18662 29640
rect 19334 29628 19340 29640
rect 19295 29600 19340 29628
rect 19334 29588 19340 29600
rect 19392 29588 19398 29640
rect 19518 29588 19524 29640
rect 19576 29628 19582 29640
rect 19613 29631 19671 29637
rect 19613 29628 19625 29631
rect 19576 29600 19625 29628
rect 19576 29588 19582 29600
rect 19613 29597 19625 29600
rect 19659 29628 19671 29631
rect 20070 29628 20076 29640
rect 19659 29600 20076 29628
rect 19659 29597 19671 29600
rect 19613 29591 19671 29597
rect 20070 29588 20076 29600
rect 20128 29588 20134 29640
rect 20162 29588 20168 29640
rect 20220 29628 20226 29640
rect 20441 29631 20499 29637
rect 20441 29628 20453 29631
rect 20220 29600 20453 29628
rect 20220 29588 20226 29600
rect 20441 29597 20453 29600
rect 20487 29597 20499 29631
rect 20622 29628 20628 29640
rect 20583 29600 20628 29628
rect 20441 29591 20499 29597
rect 20622 29588 20628 29600
rect 20680 29588 20686 29640
rect 20990 29588 20996 29640
rect 21048 29628 21054 29640
rect 21836 29637 21864 29668
rect 22278 29656 22284 29668
rect 22336 29696 22342 29708
rect 22738 29696 22744 29708
rect 22336 29668 22744 29696
rect 22336 29656 22342 29668
rect 22738 29656 22744 29668
rect 22796 29656 22802 29708
rect 22830 29656 22836 29708
rect 22888 29696 22894 29708
rect 23290 29696 23296 29708
rect 22888 29668 23296 29696
rect 22888 29656 22894 29668
rect 23290 29656 23296 29668
rect 23348 29696 23354 29708
rect 25222 29696 25228 29708
rect 23348 29668 23612 29696
rect 25183 29668 25228 29696
rect 23348 29656 23354 29668
rect 21177 29631 21235 29637
rect 21177 29628 21189 29631
rect 21048 29600 21189 29628
rect 21048 29588 21054 29600
rect 21177 29597 21189 29600
rect 21223 29597 21235 29631
rect 21177 29591 21235 29597
rect 21361 29631 21419 29637
rect 21361 29597 21373 29631
rect 21407 29597 21419 29631
rect 21361 29591 21419 29597
rect 21821 29631 21879 29637
rect 21821 29597 21833 29631
rect 21867 29597 21879 29631
rect 22002 29628 22008 29640
rect 21963 29600 22008 29628
rect 21821 29591 21879 29597
rect 16209 29563 16221 29566
rect 16163 29557 16221 29563
rect 16393 29563 16451 29569
rect 16393 29529 16405 29563
rect 16439 29560 16451 29563
rect 16574 29560 16580 29572
rect 16439 29532 16580 29560
rect 16439 29529 16451 29532
rect 16393 29523 16451 29529
rect 16574 29520 16580 29532
rect 16632 29560 16638 29572
rect 17678 29560 17684 29572
rect 16632 29532 17684 29560
rect 16632 29520 16638 29532
rect 17678 29520 17684 29532
rect 17736 29520 17742 29572
rect 18325 29563 18383 29569
rect 18325 29529 18337 29563
rect 18371 29560 18383 29563
rect 18616 29560 18644 29588
rect 19150 29560 19156 29572
rect 18371 29532 19156 29560
rect 18371 29529 18383 29532
rect 18325 29523 18383 29529
rect 19150 29520 19156 29532
rect 19208 29520 19214 29572
rect 21376 29560 21404 29591
rect 22002 29588 22008 29600
rect 22060 29588 22066 29640
rect 23584 29637 23612 29668
rect 25222 29656 25228 29668
rect 25280 29656 25286 29708
rect 26418 29656 26424 29708
rect 26476 29696 26482 29708
rect 26973 29699 27031 29705
rect 26973 29696 26985 29699
rect 26476 29668 26985 29696
rect 26476 29656 26482 29668
rect 26973 29665 26985 29668
rect 27019 29696 27031 29699
rect 27522 29696 27528 29708
rect 27019 29668 27528 29696
rect 27019 29665 27031 29668
rect 26973 29659 27031 29665
rect 27522 29656 27528 29668
rect 27580 29656 27586 29708
rect 27614 29656 27620 29708
rect 27672 29696 27678 29708
rect 27672 29668 28212 29696
rect 27672 29656 27678 29668
rect 23477 29631 23535 29637
rect 23477 29628 23489 29631
rect 22572 29600 23489 29628
rect 22370 29560 22376 29572
rect 21376 29532 22376 29560
rect 22370 29520 22376 29532
rect 22428 29520 22434 29572
rect 22572 29504 22600 29600
rect 23477 29597 23489 29600
rect 23523 29597 23535 29631
rect 23477 29591 23535 29597
rect 23569 29631 23627 29637
rect 23569 29597 23581 29631
rect 23615 29597 23627 29631
rect 23750 29628 23756 29640
rect 23711 29600 23756 29628
rect 23569 29591 23627 29597
rect 23750 29588 23756 29600
rect 23808 29588 23814 29640
rect 25038 29588 25044 29640
rect 25096 29628 25102 29640
rect 25133 29631 25191 29637
rect 25133 29628 25145 29631
rect 25096 29600 25145 29628
rect 25096 29588 25102 29600
rect 25133 29597 25145 29600
rect 25179 29628 25191 29631
rect 25774 29628 25780 29640
rect 25179 29600 25780 29628
rect 25179 29597 25191 29600
rect 25133 29591 25191 29597
rect 25774 29588 25780 29600
rect 25832 29588 25838 29640
rect 25958 29588 25964 29640
rect 26016 29628 26022 29640
rect 26513 29631 26571 29637
rect 26513 29628 26525 29631
rect 26016 29600 26525 29628
rect 26016 29588 26022 29600
rect 26513 29597 26525 29600
rect 26559 29597 26571 29631
rect 26513 29591 26571 29597
rect 26789 29631 26847 29637
rect 26789 29597 26801 29631
rect 26835 29628 26847 29631
rect 26878 29628 26884 29640
rect 26835 29600 26884 29628
rect 26835 29597 26847 29600
rect 26789 29591 26847 29597
rect 26878 29588 26884 29600
rect 26936 29588 26942 29640
rect 27154 29588 27160 29640
rect 27212 29628 27218 29640
rect 28184 29637 28212 29668
rect 27893 29631 27951 29637
rect 27893 29628 27905 29631
rect 27212 29600 27905 29628
rect 27212 29588 27218 29600
rect 27893 29597 27905 29600
rect 27939 29597 27951 29631
rect 27893 29591 27951 29597
rect 28169 29631 28227 29637
rect 28169 29597 28181 29631
rect 28215 29597 28227 29631
rect 28169 29591 28227 29597
rect 28350 29588 28356 29640
rect 28408 29628 28414 29640
rect 28997 29631 29055 29637
rect 28408 29600 28501 29628
rect 28408 29588 28414 29600
rect 28997 29597 29009 29631
rect 29043 29628 29055 29631
rect 29362 29628 29368 29640
rect 29043 29600 29368 29628
rect 29043 29597 29055 29600
rect 28997 29591 29055 29597
rect 29362 29588 29368 29600
rect 29420 29588 29426 29640
rect 29546 29628 29552 29640
rect 29507 29600 29552 29628
rect 29546 29588 29552 29600
rect 29604 29588 29610 29640
rect 29822 29628 29828 29640
rect 29783 29600 29828 29628
rect 29822 29588 29828 29600
rect 29880 29588 29886 29640
rect 31312 29637 31340 29736
rect 31386 29724 31392 29736
rect 31444 29724 31450 29776
rect 31726 29736 33272 29764
rect 31297 29631 31355 29637
rect 31297 29597 31309 29631
rect 31343 29597 31355 29631
rect 31478 29628 31484 29640
rect 31439 29600 31484 29628
rect 31297 29591 31355 29597
rect 31478 29588 31484 29600
rect 31536 29588 31542 29640
rect 22649 29563 22707 29569
rect 22649 29529 22661 29563
rect 22695 29560 22707 29563
rect 23768 29560 23796 29588
rect 22695 29532 23796 29560
rect 22695 29529 22707 29532
rect 22649 29523 22707 29529
rect 24486 29520 24492 29572
rect 24544 29560 24550 29572
rect 26896 29560 26924 29588
rect 28368 29560 28396 29588
rect 24544 29532 26648 29560
rect 26896 29532 28396 29560
rect 30285 29563 30343 29569
rect 24544 29520 24550 29532
rect 15470 29492 15476 29504
rect 15431 29464 15476 29492
rect 15470 29452 15476 29464
rect 15528 29452 15534 29504
rect 18414 29452 18420 29504
rect 18472 29492 18478 29504
rect 18525 29495 18583 29501
rect 18525 29492 18537 29495
rect 18472 29464 18537 29492
rect 18472 29452 18478 29464
rect 18525 29461 18537 29464
rect 18571 29461 18583 29495
rect 19426 29492 19432 29504
rect 19387 29464 19432 29492
rect 18525 29455 18583 29461
rect 19426 29452 19432 29464
rect 19484 29452 19490 29504
rect 20254 29492 20260 29504
rect 20215 29464 20260 29492
rect 20254 29452 20260 29464
rect 20312 29452 20318 29504
rect 21910 29492 21916 29504
rect 21871 29464 21916 29492
rect 21910 29452 21916 29464
rect 21968 29452 21974 29504
rect 22554 29452 22560 29504
rect 22612 29492 22618 29504
rect 23658 29501 23664 29504
rect 22849 29495 22907 29501
rect 22849 29492 22861 29495
rect 22612 29464 22861 29492
rect 22612 29452 22618 29464
rect 22849 29461 22861 29464
rect 22895 29461 22907 29495
rect 22849 29455 22907 29461
rect 23654 29455 23664 29501
rect 23716 29492 23722 29504
rect 24397 29495 24455 29501
rect 23716 29464 23754 29492
rect 23658 29452 23664 29455
rect 23716 29452 23722 29464
rect 24397 29461 24409 29495
rect 24443 29492 24455 29495
rect 24854 29492 24860 29504
rect 24443 29464 24860 29492
rect 24443 29461 24455 29464
rect 24397 29455 24455 29461
rect 24854 29452 24860 29464
rect 24912 29452 24918 29504
rect 25682 29452 25688 29504
rect 25740 29492 25746 29504
rect 26620 29501 26648 29532
rect 30285 29529 30297 29563
rect 30331 29560 30343 29563
rect 31726 29560 31754 29736
rect 33134 29696 33140 29708
rect 33095 29668 33140 29696
rect 33134 29656 33140 29668
rect 33192 29656 33198 29708
rect 33244 29696 33272 29736
rect 33318 29724 33324 29776
rect 33376 29764 33382 29776
rect 34808 29764 34836 29795
rect 35986 29792 35992 29804
rect 36044 29792 36050 29844
rect 36081 29835 36139 29841
rect 36081 29801 36093 29835
rect 36127 29832 36139 29835
rect 37458 29832 37464 29844
rect 36127 29804 37464 29832
rect 36127 29801 36139 29804
rect 36081 29795 36139 29801
rect 37458 29792 37464 29804
rect 37516 29792 37522 29844
rect 35342 29764 35348 29776
rect 33376 29736 34836 29764
rect 35303 29736 35348 29764
rect 33376 29724 33382 29736
rect 35342 29724 35348 29736
rect 35400 29724 35406 29776
rect 34238 29696 34244 29708
rect 33244 29668 34244 29696
rect 34238 29656 34244 29668
rect 34296 29656 34302 29708
rect 35894 29696 35900 29708
rect 35855 29668 35900 29696
rect 35894 29656 35900 29668
rect 35952 29696 35958 29708
rect 48130 29696 48136 29708
rect 35952 29668 36768 29696
rect 48091 29668 48136 29696
rect 35952 29656 35958 29668
rect 32490 29628 32496 29640
rect 32451 29600 32496 29628
rect 32490 29588 32496 29600
rect 32548 29588 32554 29640
rect 32674 29628 32680 29640
rect 32635 29600 32680 29628
rect 32674 29588 32680 29600
rect 32732 29588 32738 29640
rect 33594 29628 33600 29640
rect 33507 29600 33600 29628
rect 33594 29588 33600 29600
rect 33652 29588 33658 29640
rect 33686 29588 33692 29640
rect 33744 29628 33750 29640
rect 35802 29628 35808 29640
rect 33744 29600 35808 29628
rect 33744 29588 33750 29600
rect 35802 29588 35808 29600
rect 35860 29588 35866 29640
rect 36740 29637 36768 29668
rect 48130 29656 48136 29668
rect 48188 29656 48194 29708
rect 36725 29631 36783 29637
rect 36725 29597 36737 29631
rect 36771 29597 36783 29631
rect 36725 29591 36783 29597
rect 36817 29631 36875 29637
rect 36817 29597 36829 29631
rect 36863 29597 36875 29631
rect 36817 29591 36875 29597
rect 30331 29532 31754 29560
rect 32585 29563 32643 29569
rect 30331 29529 30343 29532
rect 30285 29523 30343 29529
rect 32585 29529 32597 29563
rect 32631 29560 32643 29563
rect 33612 29560 33640 29588
rect 32631 29532 33640 29560
rect 32631 29529 32643 29532
rect 32585 29523 32643 29529
rect 34606 29520 34612 29572
rect 34664 29560 34670 29572
rect 35345 29563 35403 29569
rect 35345 29560 35357 29563
rect 34664 29532 35357 29560
rect 34664 29520 34670 29532
rect 35345 29529 35357 29532
rect 35391 29529 35403 29563
rect 35820 29560 35848 29588
rect 36832 29560 36860 29591
rect 46382 29588 46388 29640
rect 46440 29628 46446 29640
rect 47857 29631 47915 29637
rect 47857 29628 47869 29631
rect 46440 29600 47869 29628
rect 46440 29588 46446 29600
rect 47857 29597 47869 29600
rect 47903 29597 47915 29631
rect 47857 29591 47915 29597
rect 35820 29532 36860 29560
rect 35345 29523 35403 29529
rect 25961 29495 26019 29501
rect 25961 29492 25973 29495
rect 25740 29464 25973 29492
rect 25740 29452 25746 29464
rect 25961 29461 25973 29464
rect 26007 29461 26019 29495
rect 25961 29455 26019 29461
rect 26605 29495 26663 29501
rect 26605 29461 26617 29495
rect 26651 29461 26663 29495
rect 26605 29455 26663 29461
rect 27249 29495 27307 29501
rect 27249 29461 27261 29495
rect 27295 29492 27307 29495
rect 28258 29492 28264 29504
rect 27295 29464 28264 29492
rect 27295 29461 27307 29464
rect 27249 29455 27307 29461
rect 28258 29452 28264 29464
rect 28316 29452 28322 29504
rect 29638 29452 29644 29504
rect 29696 29492 29702 29504
rect 29733 29495 29791 29501
rect 29733 29492 29745 29495
rect 29696 29464 29745 29492
rect 29696 29452 29702 29464
rect 29733 29461 29745 29464
rect 29779 29461 29791 29495
rect 29733 29455 29791 29461
rect 30495 29495 30553 29501
rect 30495 29461 30507 29495
rect 30541 29492 30553 29495
rect 30926 29492 30932 29504
rect 30541 29464 30932 29492
rect 30541 29461 30553 29464
rect 30495 29455 30553 29461
rect 30926 29452 30932 29464
rect 30984 29452 30990 29504
rect 32030 29492 32036 29504
rect 31991 29464 32036 29492
rect 32030 29452 32036 29464
rect 32088 29452 32094 29504
rect 33410 29492 33416 29504
rect 33371 29464 33416 29492
rect 33410 29452 33416 29464
rect 33468 29452 33474 29504
rect 33505 29495 33563 29501
rect 33505 29461 33517 29495
rect 33551 29492 33563 29495
rect 33686 29492 33692 29504
rect 33551 29464 33692 29492
rect 33551 29461 33563 29464
rect 33505 29455 33563 29461
rect 33686 29452 33692 29464
rect 33744 29452 33750 29504
rect 36538 29492 36544 29504
rect 36499 29464 36544 29492
rect 36538 29452 36544 29464
rect 36596 29452 36602 29504
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 16117 29291 16175 29297
rect 16117 29257 16129 29291
rect 16163 29288 16175 29291
rect 16850 29288 16856 29300
rect 16163 29260 16856 29288
rect 16163 29257 16175 29260
rect 16117 29251 16175 29257
rect 16850 29248 16856 29260
rect 16908 29248 16914 29300
rect 17034 29288 17040 29300
rect 16995 29260 17040 29288
rect 17034 29248 17040 29260
rect 17092 29248 17098 29300
rect 17678 29288 17684 29300
rect 17639 29260 17684 29288
rect 17678 29248 17684 29260
rect 17736 29248 17742 29300
rect 18874 29288 18880 29300
rect 18835 29260 18880 29288
rect 18874 29248 18880 29260
rect 18932 29248 18938 29300
rect 19245 29291 19303 29297
rect 19245 29257 19257 29291
rect 19291 29288 19303 29291
rect 19334 29288 19340 29300
rect 19291 29260 19340 29288
rect 19291 29257 19303 29260
rect 19245 29251 19303 29257
rect 19334 29248 19340 29260
rect 19392 29288 19398 29300
rect 19797 29291 19855 29297
rect 19797 29288 19809 29291
rect 19392 29260 19809 29288
rect 19392 29248 19398 29260
rect 19797 29257 19809 29260
rect 19843 29257 19855 29291
rect 20990 29288 20996 29300
rect 20951 29260 20996 29288
rect 19797 29251 19855 29257
rect 20990 29248 20996 29260
rect 21048 29248 21054 29300
rect 22554 29288 22560 29300
rect 22515 29260 22560 29288
rect 22554 29248 22560 29260
rect 22612 29248 22618 29300
rect 23290 29288 23296 29300
rect 23251 29260 23296 29288
rect 23290 29248 23296 29260
rect 23348 29248 23354 29300
rect 23845 29291 23903 29297
rect 23845 29257 23857 29291
rect 23891 29288 23903 29291
rect 23934 29288 23940 29300
rect 23891 29260 23940 29288
rect 23891 29257 23903 29260
rect 23845 29251 23903 29257
rect 23934 29248 23940 29260
rect 23992 29248 23998 29300
rect 24762 29248 24768 29300
rect 24820 29288 24826 29300
rect 27065 29291 27123 29297
rect 27065 29288 27077 29291
rect 24820 29260 27077 29288
rect 24820 29248 24826 29260
rect 27065 29257 27077 29260
rect 27111 29257 27123 29291
rect 27065 29251 27123 29257
rect 27157 29291 27215 29297
rect 27157 29257 27169 29291
rect 27203 29288 27215 29291
rect 27614 29288 27620 29300
rect 27203 29260 27620 29288
rect 27203 29257 27215 29260
rect 27157 29251 27215 29257
rect 27614 29248 27620 29260
rect 27672 29248 27678 29300
rect 28258 29288 28264 29300
rect 28219 29260 28264 29288
rect 28258 29248 28264 29260
rect 28316 29248 28322 29300
rect 28445 29291 28503 29297
rect 28445 29257 28457 29291
rect 28491 29288 28503 29291
rect 28718 29288 28724 29300
rect 28491 29260 28724 29288
rect 28491 29257 28503 29260
rect 28445 29251 28503 29257
rect 28718 29248 28724 29260
rect 28776 29248 28782 29300
rect 30466 29288 30472 29300
rect 30427 29260 30472 29288
rect 30466 29248 30472 29260
rect 30524 29248 30530 29300
rect 30926 29288 30932 29300
rect 30887 29260 30932 29288
rect 30926 29248 30932 29260
rect 30984 29248 30990 29300
rect 33134 29248 33140 29300
rect 33192 29288 33198 29300
rect 33229 29291 33287 29297
rect 33229 29288 33241 29291
rect 33192 29260 33241 29288
rect 33192 29248 33198 29260
rect 33229 29257 33241 29260
rect 33275 29257 33287 29291
rect 33229 29251 33287 29257
rect 34790 29248 34796 29300
rect 34848 29288 34854 29300
rect 35161 29291 35219 29297
rect 35161 29288 35173 29291
rect 34848 29260 35173 29288
rect 34848 29248 34854 29260
rect 35161 29257 35173 29260
rect 35207 29257 35219 29291
rect 35802 29288 35808 29300
rect 35763 29260 35808 29288
rect 35161 29251 35219 29257
rect 35802 29248 35808 29260
rect 35860 29248 35866 29300
rect 48130 29288 48136 29300
rect 48091 29260 48136 29288
rect 48130 29248 48136 29260
rect 48188 29248 48194 29300
rect 16669 29223 16727 29229
rect 16669 29220 16681 29223
rect 15948 29192 16681 29220
rect 15948 29161 15976 29192
rect 16669 29189 16681 29192
rect 16715 29189 16727 29223
rect 16669 29183 16727 29189
rect 18414 29180 18420 29232
rect 18472 29220 18478 29232
rect 20622 29220 20628 29232
rect 18472 29192 19748 29220
rect 20583 29192 20628 29220
rect 18472 29180 18478 29192
rect 15933 29155 15991 29161
rect 15933 29152 15945 29155
rect 15396 29124 15945 29152
rect 14826 29016 14832 29028
rect 14787 28988 14832 29016
rect 14826 28976 14832 28988
rect 14884 29016 14890 29028
rect 15396 29025 15424 29124
rect 15933 29121 15945 29124
rect 15979 29121 15991 29155
rect 16114 29152 16120 29164
rect 16075 29124 16120 29152
rect 15933 29115 15991 29121
rect 16114 29112 16120 29124
rect 16172 29152 16178 29164
rect 16853 29155 16911 29161
rect 16853 29152 16865 29155
rect 16172 29124 16865 29152
rect 16172 29112 16178 29124
rect 16853 29121 16865 29124
rect 16899 29152 16911 29155
rect 17218 29152 17224 29164
rect 16899 29124 17224 29152
rect 16899 29121 16911 29124
rect 16853 29115 16911 29121
rect 17218 29112 17224 29124
rect 17276 29112 17282 29164
rect 17586 29152 17592 29164
rect 17547 29124 17592 29152
rect 17586 29112 17592 29124
rect 17644 29112 17650 29164
rect 17954 29152 17960 29164
rect 17915 29124 17960 29152
rect 17954 29112 17960 29124
rect 18012 29112 18018 29164
rect 18782 29152 18788 29164
rect 18743 29124 18788 29152
rect 18782 29112 18788 29124
rect 18840 29112 18846 29164
rect 19058 29152 19064 29164
rect 18971 29124 19064 29152
rect 19058 29112 19064 29124
rect 19116 29112 19122 29164
rect 19150 29112 19156 29164
rect 19208 29152 19214 29164
rect 19518 29152 19524 29164
rect 19208 29124 19524 29152
rect 19208 29112 19214 29124
rect 19518 29112 19524 29124
rect 19576 29112 19582 29164
rect 19720 29161 19748 29192
rect 20622 29180 20628 29192
rect 20680 29180 20686 29232
rect 20841 29223 20899 29229
rect 20841 29189 20853 29223
rect 20887 29220 20899 29223
rect 21082 29220 21088 29232
rect 20887 29192 21088 29220
rect 20887 29189 20899 29192
rect 20841 29183 20899 29189
rect 21082 29180 21088 29192
rect 21140 29180 21146 29232
rect 29457 29223 29515 29229
rect 24504 29192 25636 29220
rect 24504 29164 24532 29192
rect 19705 29155 19763 29161
rect 19705 29121 19717 29155
rect 19751 29121 19763 29155
rect 19705 29115 19763 29121
rect 19794 29112 19800 29164
rect 19852 29152 19858 29164
rect 19981 29155 20039 29161
rect 19981 29152 19993 29155
rect 19852 29124 19993 29152
rect 19852 29112 19858 29124
rect 19981 29121 19993 29124
rect 20027 29121 20039 29155
rect 19981 29115 20039 29121
rect 22002 29112 22008 29164
rect 22060 29152 22066 29164
rect 22189 29155 22247 29161
rect 22189 29152 22201 29155
rect 22060 29124 22201 29152
rect 22060 29112 22066 29124
rect 22189 29121 22201 29124
rect 22235 29152 22247 29155
rect 23014 29152 23020 29164
rect 22235 29124 22508 29152
rect 22975 29124 23020 29152
rect 22235 29121 22247 29124
rect 22189 29115 22247 29121
rect 17865 29087 17923 29093
rect 17865 29053 17877 29087
rect 17911 29084 17923 29087
rect 18230 29084 18236 29096
rect 17911 29056 18236 29084
rect 17911 29053 17923 29056
rect 17865 29047 17923 29053
rect 18230 29044 18236 29056
rect 18288 29084 18294 29096
rect 19076 29084 19104 29112
rect 20070 29084 20076 29096
rect 18288 29056 19104 29084
rect 19168 29056 20076 29084
rect 18288 29044 18294 29056
rect 15381 29019 15439 29025
rect 15381 29016 15393 29019
rect 14884 28988 15393 29016
rect 14884 28976 14890 28988
rect 15381 28985 15393 28988
rect 15427 28985 15439 29019
rect 15381 28979 15439 28985
rect 15470 28976 15476 29028
rect 15528 29016 15534 29028
rect 16942 29016 16948 29028
rect 15528 28988 16948 29016
rect 15528 28976 15534 28988
rect 16942 28976 16948 28988
rect 17000 29016 17006 29028
rect 17770 29016 17776 29028
rect 17000 28988 17776 29016
rect 17000 28976 17006 28988
rect 17770 28976 17776 28988
rect 17828 28976 17834 29028
rect 18049 29019 18107 29025
rect 18049 28985 18061 29019
rect 18095 29016 18107 29019
rect 19168 29016 19196 29056
rect 20070 29044 20076 29056
rect 20128 29044 20134 29096
rect 22094 29044 22100 29096
rect 22152 29084 22158 29096
rect 22281 29087 22339 29093
rect 22281 29084 22293 29087
rect 22152 29056 22293 29084
rect 22152 29044 22158 29056
rect 22281 29053 22293 29056
rect 22327 29053 22339 29087
rect 22480 29084 22508 29124
rect 23014 29112 23020 29124
rect 23072 29112 23078 29164
rect 23658 29112 23664 29164
rect 23716 29152 23722 29164
rect 23753 29155 23811 29161
rect 23753 29152 23765 29155
rect 23716 29124 23765 29152
rect 23716 29112 23722 29124
rect 23753 29121 23765 29124
rect 23799 29121 23811 29155
rect 23753 29115 23811 29121
rect 23937 29155 23995 29161
rect 23937 29121 23949 29155
rect 23983 29121 23995 29155
rect 24486 29152 24492 29164
rect 24447 29124 24492 29152
rect 23937 29115 23995 29121
rect 23293 29087 23351 29093
rect 23293 29084 23305 29087
rect 22480 29056 23305 29084
rect 22281 29047 22339 29053
rect 23293 29053 23305 29056
rect 23339 29053 23351 29087
rect 23952 29084 23980 29115
rect 24486 29112 24492 29124
rect 24544 29112 24550 29164
rect 24581 29155 24639 29161
rect 24581 29121 24593 29155
rect 24627 29152 24639 29155
rect 24670 29152 24676 29164
rect 24627 29124 24676 29152
rect 24627 29121 24639 29124
rect 24581 29115 24639 29121
rect 24670 29112 24676 29124
rect 24728 29112 24734 29164
rect 24765 29155 24823 29161
rect 24765 29121 24777 29155
rect 24811 29152 24823 29155
rect 25130 29152 25136 29164
rect 24811 29124 25136 29152
rect 24811 29121 24823 29124
rect 24765 29115 24823 29121
rect 24780 29084 24808 29115
rect 25130 29112 25136 29124
rect 25188 29112 25194 29164
rect 25608 29161 25636 29192
rect 29457 29189 29469 29223
rect 29503 29220 29515 29223
rect 29730 29220 29736 29232
rect 29503 29192 29736 29220
rect 29503 29189 29515 29192
rect 29457 29183 29515 29189
rect 29730 29180 29736 29192
rect 29788 29180 29794 29232
rect 32490 29180 32496 29232
rect 32548 29220 32554 29232
rect 32861 29223 32919 29229
rect 32861 29220 32873 29223
rect 32548 29192 32873 29220
rect 32548 29180 32554 29192
rect 32861 29189 32873 29192
rect 32907 29220 32919 29223
rect 33962 29220 33968 29232
rect 32907 29192 33968 29220
rect 32907 29189 32919 29192
rect 32861 29183 32919 29189
rect 33962 29180 33968 29192
rect 34020 29220 34026 29232
rect 36265 29223 36323 29229
rect 36265 29220 36277 29223
rect 34020 29192 36277 29220
rect 34020 29180 34026 29192
rect 36265 29189 36277 29192
rect 36311 29189 36323 29223
rect 36265 29183 36323 29189
rect 25593 29155 25651 29161
rect 25593 29121 25605 29155
rect 25639 29121 25651 29155
rect 25593 29115 25651 29121
rect 25682 29112 25688 29164
rect 25740 29152 25746 29164
rect 26970 29152 26976 29164
rect 25740 29124 25785 29152
rect 26931 29124 26976 29152
rect 25740 29112 25746 29124
rect 26970 29112 26976 29124
rect 27028 29112 27034 29164
rect 27982 29112 27988 29164
rect 28040 29152 28046 29164
rect 28077 29155 28135 29161
rect 28077 29152 28089 29155
rect 28040 29124 28089 29152
rect 28040 29112 28046 29124
rect 28077 29121 28089 29124
rect 28123 29121 28135 29155
rect 28077 29115 28135 29121
rect 28166 29112 28172 29164
rect 28224 29152 28230 29164
rect 29362 29152 29368 29164
rect 28224 29124 28269 29152
rect 29323 29124 29368 29152
rect 28224 29112 28230 29124
rect 29362 29112 29368 29124
rect 29420 29112 29426 29164
rect 29641 29155 29699 29161
rect 29641 29121 29653 29155
rect 29687 29152 29699 29155
rect 29914 29152 29920 29164
rect 29687 29124 29920 29152
rect 29687 29121 29699 29124
rect 29641 29115 29699 29121
rect 29914 29112 29920 29124
rect 29972 29112 29978 29164
rect 30098 29152 30104 29164
rect 30059 29124 30104 29152
rect 30098 29112 30104 29124
rect 30156 29112 30162 29164
rect 30190 29112 30196 29164
rect 30248 29152 30254 29164
rect 31205 29155 31263 29161
rect 31205 29152 31217 29155
rect 30248 29124 31217 29152
rect 30248 29112 30254 29124
rect 31205 29121 31217 29124
rect 31251 29121 31263 29155
rect 31205 29115 31263 29121
rect 32674 29112 32680 29164
rect 32732 29152 32738 29164
rect 33045 29155 33103 29161
rect 33045 29152 33057 29155
rect 32732 29124 33057 29152
rect 32732 29112 32738 29124
rect 33045 29121 33057 29124
rect 33091 29121 33103 29155
rect 33045 29115 33103 29121
rect 34333 29155 34391 29161
rect 34333 29121 34345 29155
rect 34379 29152 34391 29155
rect 35437 29155 35495 29161
rect 35437 29152 35449 29155
rect 34379 29124 35449 29152
rect 34379 29121 34391 29124
rect 34333 29115 34391 29121
rect 35437 29121 35449 29124
rect 35483 29152 35495 29155
rect 36538 29152 36544 29164
rect 35483 29124 36544 29152
rect 35483 29121 35495 29124
rect 35437 29115 35495 29121
rect 23952 29056 24808 29084
rect 24949 29087 25007 29093
rect 23293 29047 23351 29053
rect 24949 29053 24961 29087
rect 24995 29084 25007 29087
rect 25409 29087 25467 29093
rect 25409 29084 25421 29087
rect 24995 29056 25421 29084
rect 24995 29053 25007 29056
rect 24949 29047 25007 29053
rect 25409 29053 25421 29056
rect 25455 29053 25467 29087
rect 26326 29084 26332 29096
rect 25409 29047 25467 29053
rect 25516 29056 26332 29084
rect 25516 29025 25544 29056
rect 26326 29044 26332 29056
rect 26384 29084 26390 29096
rect 27433 29087 27491 29093
rect 27433 29084 27445 29087
rect 26384 29056 27445 29084
rect 26384 29044 26390 29056
rect 27433 29053 27445 29056
rect 27479 29053 27491 29087
rect 30116 29084 30144 29112
rect 30929 29087 30987 29093
rect 30929 29084 30941 29087
rect 30116 29056 30941 29084
rect 27433 29047 27491 29053
rect 30929 29053 30941 29056
rect 30975 29053 30987 29087
rect 30929 29047 30987 29053
rect 25501 29019 25559 29025
rect 18095 28988 19196 29016
rect 19904 28988 20208 29016
rect 18095 28985 18107 28988
rect 18049 28979 18107 28985
rect 18325 28951 18383 28957
rect 18325 28917 18337 28951
rect 18371 28948 18383 28951
rect 19904 28948 19932 28988
rect 18371 28920 19932 28948
rect 18371 28917 18383 28920
rect 18325 28911 18383 28917
rect 19978 28908 19984 28960
rect 20036 28948 20042 28960
rect 20180 28948 20208 28988
rect 25501 28985 25513 29019
rect 25547 28985 25559 29019
rect 27890 29016 27896 29028
rect 27851 28988 27896 29016
rect 25501 28979 25559 28985
rect 27890 28976 27896 28988
rect 27948 28976 27954 29028
rect 31113 29019 31171 29025
rect 31113 29016 31125 29019
rect 30116 28988 31125 29016
rect 20530 28948 20536 28960
rect 20036 28920 20081 28948
rect 20180 28920 20536 28948
rect 20036 28908 20042 28920
rect 20530 28908 20536 28920
rect 20588 28948 20594 28960
rect 20809 28951 20867 28957
rect 20809 28948 20821 28951
rect 20588 28920 20821 28948
rect 20588 28908 20594 28920
rect 20809 28917 20821 28920
rect 20855 28917 20867 28951
rect 22370 28948 22376 28960
rect 22283 28920 22376 28948
rect 20809 28911 20867 28917
rect 22370 28908 22376 28920
rect 22428 28948 22434 28960
rect 22922 28948 22928 28960
rect 22428 28920 22928 28948
rect 22428 28908 22434 28920
rect 22922 28908 22928 28920
rect 22980 28948 22986 28960
rect 23109 28951 23167 28957
rect 23109 28948 23121 28951
rect 22980 28920 23121 28948
rect 22980 28908 22986 28920
rect 23109 28917 23121 28920
rect 23155 28917 23167 28951
rect 23109 28911 23167 28917
rect 24854 28908 24860 28960
rect 24912 28948 24918 28960
rect 25682 28948 25688 28960
rect 24912 28920 25688 28948
rect 24912 28908 24918 28920
rect 25682 28908 25688 28920
rect 25740 28908 25746 28960
rect 26421 28951 26479 28957
rect 26421 28917 26433 28951
rect 26467 28948 26479 28951
rect 26510 28948 26516 28960
rect 26467 28920 26516 28948
rect 26467 28917 26479 28920
rect 26421 28911 26479 28917
rect 26510 28908 26516 28920
rect 26568 28908 26574 28960
rect 30116 28957 30144 28988
rect 31113 28985 31125 28988
rect 31159 28985 31171 29019
rect 33060 29016 33088 29115
rect 36538 29112 36544 29124
rect 36596 29112 36602 29164
rect 33410 29044 33416 29096
rect 33468 29084 33474 29096
rect 34241 29087 34299 29093
rect 34241 29084 34253 29087
rect 33468 29056 34253 29084
rect 33468 29044 33474 29056
rect 34241 29053 34253 29056
rect 34287 29053 34299 29087
rect 34241 29047 34299 29053
rect 34425 29087 34483 29093
rect 34425 29053 34437 29087
rect 34471 29053 34483 29087
rect 34425 29047 34483 29053
rect 34330 29016 34336 29028
rect 33060 28988 34336 29016
rect 31113 28979 31171 28985
rect 34330 28976 34336 28988
rect 34388 28976 34394 29028
rect 34440 29016 34468 29047
rect 34514 29044 34520 29096
rect 34572 29084 34578 29096
rect 35345 29087 35403 29093
rect 34572 29056 34617 29084
rect 34572 29044 34578 29056
rect 35345 29053 35357 29087
rect 35391 29084 35403 29087
rect 37274 29084 37280 29096
rect 35391 29056 37280 29084
rect 35391 29053 35403 29056
rect 35345 29047 35403 29053
rect 35360 29016 35388 29047
rect 37274 29044 37280 29056
rect 37332 29044 37338 29096
rect 34440 28988 35388 29016
rect 29641 28951 29699 28957
rect 29641 28917 29653 28951
rect 29687 28948 29699 28951
rect 30101 28951 30159 28957
rect 30101 28948 30113 28951
rect 29687 28920 30113 28948
rect 29687 28917 29699 28920
rect 29641 28911 29699 28917
rect 30101 28917 30113 28920
rect 30147 28917 30159 28951
rect 30101 28911 30159 28917
rect 31938 28908 31944 28960
rect 31996 28948 32002 28960
rect 32125 28951 32183 28957
rect 32125 28948 32137 28951
rect 31996 28920 32137 28948
rect 31996 28908 32002 28920
rect 32125 28917 32137 28920
rect 32171 28917 32183 28951
rect 32125 28911 32183 28917
rect 34701 28951 34759 28957
rect 34701 28917 34713 28951
rect 34747 28948 34759 28951
rect 34790 28948 34796 28960
rect 34747 28920 34796 28948
rect 34747 28917 34759 28920
rect 34701 28911 34759 28917
rect 34790 28908 34796 28920
rect 34848 28908 34854 28960
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 15289 28747 15347 28753
rect 15289 28713 15301 28747
rect 15335 28744 15347 28747
rect 15378 28744 15384 28756
rect 15335 28716 15384 28744
rect 15335 28713 15347 28716
rect 15289 28707 15347 28713
rect 15378 28704 15384 28716
rect 15436 28704 15442 28756
rect 18049 28747 18107 28753
rect 18049 28713 18061 28747
rect 18095 28744 18107 28747
rect 18322 28744 18328 28756
rect 18095 28716 18328 28744
rect 18095 28713 18107 28716
rect 18049 28707 18107 28713
rect 18322 28704 18328 28716
rect 18380 28744 18386 28756
rect 18874 28744 18880 28756
rect 18380 28716 18880 28744
rect 18380 28704 18386 28716
rect 18874 28704 18880 28716
rect 18932 28704 18938 28756
rect 19058 28704 19064 28756
rect 19116 28744 19122 28756
rect 19429 28747 19487 28753
rect 19429 28744 19441 28747
rect 19116 28716 19441 28744
rect 19116 28704 19122 28716
rect 19429 28713 19441 28716
rect 19475 28713 19487 28747
rect 19429 28707 19487 28713
rect 20073 28747 20131 28753
rect 20073 28713 20085 28747
rect 20119 28744 20131 28747
rect 20438 28744 20444 28756
rect 20119 28716 20444 28744
rect 20119 28713 20131 28716
rect 20073 28707 20131 28713
rect 20438 28704 20444 28716
rect 20496 28704 20502 28756
rect 23385 28747 23443 28753
rect 23385 28713 23397 28747
rect 23431 28744 23443 28747
rect 23474 28744 23480 28756
rect 23431 28716 23480 28744
rect 23431 28713 23443 28716
rect 23385 28707 23443 28713
rect 23474 28704 23480 28716
rect 23532 28744 23538 28756
rect 24210 28744 24216 28756
rect 23532 28716 24216 28744
rect 23532 28704 23538 28716
rect 24210 28704 24216 28716
rect 24268 28704 24274 28756
rect 25038 28744 25044 28756
rect 24999 28716 25044 28744
rect 25038 28704 25044 28716
rect 25096 28704 25102 28756
rect 26326 28744 26332 28756
rect 26287 28716 26332 28744
rect 26326 28704 26332 28716
rect 26384 28704 26390 28756
rect 28166 28744 28172 28756
rect 28092 28716 28172 28744
rect 17770 28636 17776 28688
rect 17828 28676 17834 28688
rect 18601 28679 18659 28685
rect 18601 28676 18613 28679
rect 17828 28648 18613 28676
rect 17828 28636 17834 28648
rect 18601 28645 18613 28648
rect 18647 28676 18659 28679
rect 20346 28676 20352 28688
rect 18647 28648 20352 28676
rect 18647 28645 18659 28648
rect 18601 28639 18659 28645
rect 20346 28636 20352 28648
rect 20404 28636 20410 28688
rect 20993 28679 21051 28685
rect 20993 28645 21005 28679
rect 21039 28676 21051 28679
rect 22922 28676 22928 28688
rect 21039 28648 22928 28676
rect 21039 28645 21051 28648
rect 20993 28639 21051 28645
rect 22922 28636 22928 28648
rect 22980 28636 22986 28688
rect 25961 28679 26019 28685
rect 25961 28645 25973 28679
rect 26007 28676 26019 28679
rect 28092 28676 28120 28716
rect 28166 28704 28172 28716
rect 28224 28704 28230 28756
rect 29638 28744 29644 28756
rect 29599 28716 29644 28744
rect 29638 28704 29644 28716
rect 29696 28704 29702 28756
rect 30190 28704 30196 28756
rect 30248 28744 30254 28756
rect 30285 28747 30343 28753
rect 30285 28744 30297 28747
rect 30248 28716 30297 28744
rect 30248 28704 30254 28716
rect 30285 28713 30297 28716
rect 30331 28713 30343 28747
rect 30285 28707 30343 28713
rect 32953 28747 33011 28753
rect 32953 28713 32965 28747
rect 32999 28713 33011 28747
rect 32953 28707 33011 28713
rect 32030 28676 32036 28688
rect 26007 28648 28120 28676
rect 26007 28645 26019 28648
rect 25961 28639 26019 28645
rect 20530 28608 20536 28620
rect 20491 28580 20536 28608
rect 20530 28568 20536 28580
rect 20588 28568 20594 28620
rect 21082 28608 21088 28620
rect 21043 28580 21088 28608
rect 21082 28568 21088 28580
rect 21140 28608 21146 28620
rect 21637 28611 21695 28617
rect 21637 28608 21649 28611
rect 21140 28580 21649 28608
rect 21140 28568 21146 28580
rect 21637 28577 21649 28580
rect 21683 28577 21695 28611
rect 21637 28571 21695 28577
rect 22465 28611 22523 28617
rect 22465 28577 22477 28611
rect 22511 28608 22523 28611
rect 22738 28608 22744 28620
rect 22511 28580 22744 28608
rect 22511 28577 22523 28580
rect 22465 28571 22523 28577
rect 22738 28568 22744 28580
rect 22796 28568 22802 28620
rect 24578 28608 24584 28620
rect 24539 28580 24584 28608
rect 24578 28568 24584 28580
rect 24636 28568 24642 28620
rect 27890 28608 27896 28620
rect 27851 28580 27896 28608
rect 27890 28568 27896 28580
rect 27948 28568 27954 28620
rect 28092 28617 28120 28648
rect 30668 28648 32036 28676
rect 28077 28611 28135 28617
rect 28077 28577 28089 28611
rect 28123 28577 28135 28611
rect 28077 28571 28135 28577
rect 28169 28611 28227 28617
rect 28169 28577 28181 28611
rect 28215 28608 28227 28611
rect 28258 28608 28264 28620
rect 28215 28580 28264 28608
rect 28215 28577 28227 28580
rect 28169 28571 28227 28577
rect 28258 28568 28264 28580
rect 28316 28568 28322 28620
rect 28353 28611 28411 28617
rect 28353 28577 28365 28611
rect 28399 28608 28411 28611
rect 29362 28608 29368 28620
rect 28399 28580 29368 28608
rect 28399 28577 28411 28580
rect 28353 28571 28411 28577
rect 29362 28568 29368 28580
rect 29420 28608 29426 28620
rect 29420 28580 29592 28608
rect 29420 28568 29426 28580
rect 16666 28500 16672 28552
rect 16724 28540 16730 28552
rect 17586 28540 17592 28552
rect 16724 28512 17592 28540
rect 16724 28500 16730 28512
rect 17586 28500 17592 28512
rect 17644 28500 17650 28552
rect 17678 28500 17684 28552
rect 17736 28540 17742 28552
rect 17865 28543 17923 28549
rect 17736 28512 17781 28540
rect 17736 28500 17742 28512
rect 17865 28509 17877 28543
rect 17911 28540 17923 28543
rect 17954 28540 17960 28552
rect 17911 28512 17960 28540
rect 17911 28509 17923 28512
rect 17865 28503 17923 28509
rect 17954 28500 17960 28512
rect 18012 28500 18018 28552
rect 19334 28540 19340 28552
rect 19295 28512 19340 28540
rect 19334 28500 19340 28512
rect 19392 28500 19398 28552
rect 19521 28543 19579 28549
rect 19521 28509 19533 28543
rect 19567 28540 19579 28543
rect 20254 28540 20260 28552
rect 19567 28512 20260 28540
rect 19567 28509 19579 28512
rect 19521 28503 19579 28509
rect 20254 28500 20260 28512
rect 20312 28500 20318 28552
rect 20622 28500 20628 28552
rect 20680 28540 20686 28552
rect 20717 28543 20775 28549
rect 20717 28540 20729 28543
rect 20680 28512 20729 28540
rect 20680 28500 20686 28512
rect 20717 28509 20729 28512
rect 20763 28509 20775 28543
rect 20717 28503 20775 28509
rect 21910 28500 21916 28552
rect 21968 28540 21974 28552
rect 22005 28543 22063 28549
rect 22005 28540 22017 28543
rect 21968 28512 22017 28540
rect 21968 28500 21974 28512
rect 22005 28509 22017 28512
rect 22051 28509 22063 28543
rect 22005 28503 22063 28509
rect 22649 28543 22707 28549
rect 22649 28509 22661 28543
rect 22695 28540 22707 28543
rect 23106 28540 23112 28552
rect 22695 28512 23112 28540
rect 22695 28509 22707 28512
rect 22649 28503 22707 28509
rect 23106 28500 23112 28512
rect 23164 28500 23170 28552
rect 24673 28543 24731 28549
rect 24673 28509 24685 28543
rect 24719 28540 24731 28543
rect 24854 28540 24860 28552
rect 24719 28512 24860 28540
rect 24719 28509 24731 28512
rect 24673 28503 24731 28509
rect 24854 28500 24860 28512
rect 24912 28500 24918 28552
rect 26237 28543 26295 28549
rect 26237 28509 26249 28543
rect 26283 28509 26295 28543
rect 26237 28503 26295 28509
rect 21821 28475 21879 28481
rect 21821 28441 21833 28475
rect 21867 28472 21879 28475
rect 22094 28472 22100 28484
rect 21867 28444 22100 28472
rect 21867 28441 21879 28444
rect 21821 28435 21879 28441
rect 22094 28432 22100 28444
rect 22152 28472 22158 28484
rect 22833 28475 22891 28481
rect 22833 28472 22845 28475
rect 22152 28444 22845 28472
rect 22152 28432 22158 28444
rect 22833 28441 22845 28444
rect 22879 28472 22891 28475
rect 23014 28472 23020 28484
rect 22879 28444 23020 28472
rect 22879 28441 22891 28444
rect 22833 28435 22891 28441
rect 23014 28432 23020 28444
rect 23072 28432 23078 28484
rect 15746 28404 15752 28416
rect 15707 28376 15752 28404
rect 15746 28364 15752 28376
rect 15804 28404 15810 28416
rect 16114 28404 16120 28416
rect 15804 28376 16120 28404
rect 15804 28364 15810 28376
rect 16114 28364 16120 28376
rect 16172 28404 16178 28416
rect 16485 28407 16543 28413
rect 16485 28404 16497 28407
rect 16172 28376 16497 28404
rect 16172 28364 16178 28376
rect 16485 28373 16497 28376
rect 16531 28373 16543 28407
rect 16485 28367 16543 28373
rect 17129 28407 17187 28413
rect 17129 28373 17141 28407
rect 17175 28404 17187 28407
rect 17954 28404 17960 28416
rect 17175 28376 17960 28404
rect 17175 28373 17187 28376
rect 17129 28367 17187 28373
rect 17954 28364 17960 28376
rect 18012 28364 18018 28416
rect 26252 28404 26280 28503
rect 26326 28500 26332 28552
rect 26384 28540 26390 28552
rect 26973 28543 27031 28549
rect 26384 28512 26429 28540
rect 26384 28500 26390 28512
rect 26973 28509 26985 28543
rect 27019 28540 27031 28543
rect 27154 28540 27160 28552
rect 27019 28512 27160 28540
rect 27019 28509 27031 28512
rect 26973 28503 27031 28509
rect 27154 28500 27160 28512
rect 27212 28500 27218 28552
rect 27982 28540 27988 28552
rect 27943 28512 27988 28540
rect 27982 28500 27988 28512
rect 28040 28500 28046 28552
rect 29564 28549 29592 28580
rect 30374 28568 30380 28620
rect 30432 28608 30438 28620
rect 30668 28617 30696 28648
rect 32030 28636 32036 28648
rect 32088 28676 32094 28688
rect 32968 28676 32996 28707
rect 34514 28704 34520 28756
rect 34572 28744 34578 28756
rect 35805 28747 35863 28753
rect 35805 28744 35817 28747
rect 34572 28716 35817 28744
rect 34572 28704 34578 28716
rect 35805 28713 35817 28716
rect 35851 28713 35863 28747
rect 35805 28707 35863 28713
rect 34606 28676 34612 28688
rect 32088 28648 32904 28676
rect 32968 28648 34612 28676
rect 32088 28636 32094 28648
rect 30653 28611 30711 28617
rect 30653 28608 30665 28611
rect 30432 28580 30665 28608
rect 30432 28568 30438 28580
rect 30653 28577 30665 28580
rect 30699 28577 30711 28611
rect 32585 28611 32643 28617
rect 32585 28608 32597 28611
rect 30653 28571 30711 28577
rect 32048 28580 32597 28608
rect 29549 28543 29607 28549
rect 29549 28509 29561 28543
rect 29595 28509 29607 28543
rect 29730 28540 29736 28552
rect 29691 28512 29736 28540
rect 29549 28503 29607 28509
rect 29730 28500 29736 28512
rect 29788 28500 29794 28552
rect 30190 28500 30196 28552
rect 30248 28540 30254 28552
rect 30469 28543 30527 28549
rect 30469 28540 30481 28543
rect 30248 28512 30481 28540
rect 30248 28500 30254 28512
rect 30469 28509 30481 28512
rect 30515 28509 30527 28543
rect 30469 28503 30527 28509
rect 31711 28543 31769 28549
rect 31711 28509 31723 28543
rect 31757 28509 31769 28543
rect 31846 28540 31852 28552
rect 31807 28512 31852 28540
rect 31711 28503 31769 28509
rect 26786 28472 26792 28484
rect 26747 28444 26792 28472
rect 26786 28432 26792 28444
rect 26844 28432 26850 28484
rect 27062 28432 27068 28484
rect 27120 28472 27126 28484
rect 31481 28475 31539 28481
rect 31481 28472 31493 28475
rect 27120 28444 31493 28472
rect 27120 28432 27126 28444
rect 31481 28441 31493 28444
rect 31527 28441 31539 28475
rect 31726 28472 31754 28503
rect 31846 28500 31852 28512
rect 31904 28500 31910 28552
rect 31962 28543 32020 28549
rect 31962 28509 31974 28543
rect 32008 28540 32020 28543
rect 32048 28540 32076 28580
rect 32585 28577 32597 28580
rect 32631 28577 32643 28611
rect 32876 28608 32904 28648
rect 34606 28636 34612 28648
rect 34664 28636 34670 28688
rect 35253 28679 35311 28685
rect 35253 28645 35265 28679
rect 35299 28676 35311 28679
rect 35434 28676 35440 28688
rect 35299 28648 35440 28676
rect 35299 28645 35311 28648
rect 35253 28639 35311 28645
rect 35434 28636 35440 28648
rect 35492 28636 35498 28688
rect 34790 28608 34796 28620
rect 32876 28580 33640 28608
rect 34751 28580 34796 28608
rect 32585 28571 32643 28577
rect 32008 28512 32076 28540
rect 32125 28543 32183 28549
rect 32008 28509 32020 28512
rect 31962 28503 32020 28509
rect 32125 28509 32137 28543
rect 32171 28540 32183 28543
rect 32490 28540 32496 28552
rect 32171 28512 32496 28540
rect 32171 28509 32183 28512
rect 32125 28503 32183 28509
rect 32490 28500 32496 28512
rect 32548 28500 32554 28552
rect 33045 28543 33103 28549
rect 33045 28509 33057 28543
rect 33091 28540 33103 28543
rect 33410 28540 33416 28552
rect 33091 28512 33416 28540
rect 33091 28509 33103 28512
rect 33045 28503 33103 28509
rect 33410 28500 33416 28512
rect 33468 28500 33474 28552
rect 32306 28472 32312 28484
rect 31726 28444 32312 28472
rect 31481 28435 31539 28441
rect 32306 28432 32312 28444
rect 32364 28432 32370 28484
rect 33505 28475 33563 28481
rect 33505 28472 33517 28475
rect 32508 28444 33517 28472
rect 26878 28404 26884 28416
rect 26252 28376 26884 28404
rect 26878 28364 26884 28376
rect 26936 28404 26942 28416
rect 27157 28407 27215 28413
rect 27157 28404 27169 28407
rect 26936 28376 27169 28404
rect 26936 28364 26942 28376
rect 27157 28373 27169 28376
rect 27203 28373 27215 28407
rect 28810 28404 28816 28416
rect 28771 28376 28816 28404
rect 27157 28367 27215 28373
rect 28810 28364 28816 28376
rect 28868 28404 28874 28416
rect 29454 28404 29460 28416
rect 28868 28376 29460 28404
rect 28868 28364 28874 28376
rect 29454 28364 29460 28376
rect 29512 28364 29518 28416
rect 31018 28364 31024 28416
rect 31076 28404 31082 28416
rect 32508 28404 32536 28444
rect 33505 28441 33517 28444
rect 33551 28441 33563 28475
rect 33612 28472 33640 28580
rect 34790 28568 34796 28580
rect 34848 28568 34854 28620
rect 34054 28500 34060 28552
rect 34112 28540 34118 28552
rect 34885 28543 34943 28549
rect 34885 28540 34897 28543
rect 34112 28512 34897 28540
rect 34112 28500 34118 28512
rect 34885 28509 34897 28512
rect 34931 28509 34943 28543
rect 34885 28503 34943 28509
rect 35342 28500 35348 28552
rect 35400 28540 35406 28552
rect 35713 28543 35771 28549
rect 35713 28540 35725 28543
rect 35400 28512 35725 28540
rect 35400 28500 35406 28512
rect 35713 28509 35725 28512
rect 35759 28509 35771 28543
rect 35713 28503 35771 28509
rect 33612 28444 34192 28472
rect 33505 28435 33563 28441
rect 34164 28413 34192 28444
rect 31076 28376 32536 28404
rect 34149 28407 34207 28413
rect 31076 28364 31082 28376
rect 34149 28373 34161 28407
rect 34195 28404 34207 28407
rect 45278 28404 45284 28416
rect 34195 28376 45284 28404
rect 34195 28373 34207 28376
rect 34149 28367 34207 28373
rect 45278 28364 45284 28376
rect 45336 28364 45342 28416
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 18414 28200 18420 28212
rect 18375 28172 18420 28200
rect 18414 28160 18420 28172
rect 18472 28160 18478 28212
rect 19061 28203 19119 28209
rect 19061 28169 19073 28203
rect 19107 28200 19119 28203
rect 20622 28200 20628 28212
rect 19107 28172 20628 28200
rect 19107 28169 19119 28172
rect 19061 28163 19119 28169
rect 20622 28160 20628 28172
rect 20680 28160 20686 28212
rect 27062 28200 27068 28212
rect 20732 28172 27068 28200
rect 18322 28132 18328 28144
rect 18283 28104 18328 28132
rect 18322 28092 18328 28104
rect 18380 28092 18386 28144
rect 18509 28135 18567 28141
rect 18509 28101 18521 28135
rect 18555 28132 18567 28135
rect 18782 28132 18788 28144
rect 18555 28104 18788 28132
rect 18555 28101 18567 28104
rect 18509 28095 18567 28101
rect 18782 28092 18788 28104
rect 18840 28132 18846 28144
rect 20732 28132 20760 28172
rect 27062 28160 27068 28172
rect 27120 28160 27126 28212
rect 27890 28160 27896 28212
rect 27948 28200 27954 28212
rect 27985 28203 28043 28209
rect 27985 28200 27997 28203
rect 27948 28172 27997 28200
rect 27948 28160 27954 28172
rect 27985 28169 27997 28172
rect 28031 28169 28043 28203
rect 27985 28163 28043 28169
rect 28629 28203 28687 28209
rect 28629 28169 28641 28203
rect 28675 28200 28687 28203
rect 29730 28200 29736 28212
rect 28675 28172 29736 28200
rect 28675 28169 28687 28172
rect 28629 28163 28687 28169
rect 29730 28160 29736 28172
rect 29788 28160 29794 28212
rect 29914 28160 29920 28212
rect 29972 28200 29978 28212
rect 30285 28203 30343 28209
rect 30285 28200 30297 28203
rect 29972 28172 30297 28200
rect 29972 28160 29978 28172
rect 30285 28169 30297 28172
rect 30331 28169 30343 28203
rect 30285 28163 30343 28169
rect 30929 28203 30987 28209
rect 30929 28169 30941 28203
rect 30975 28200 30987 28203
rect 31846 28200 31852 28212
rect 30975 28172 31852 28200
rect 30975 28169 30987 28172
rect 30929 28163 30987 28169
rect 31846 28160 31852 28172
rect 31904 28160 31910 28212
rect 32214 28200 32220 28212
rect 32175 28172 32220 28200
rect 32214 28160 32220 28172
rect 32272 28160 32278 28212
rect 32490 28160 32496 28212
rect 32548 28200 32554 28212
rect 34057 28203 34115 28209
rect 32548 28172 34008 28200
rect 32548 28160 32554 28172
rect 18840 28104 19380 28132
rect 18840 28092 18846 28104
rect 1673 28067 1731 28073
rect 1673 28033 1685 28067
rect 1719 28064 1731 28067
rect 18230 28064 18236 28076
rect 1719 28036 2268 28064
rect 18191 28036 18236 28064
rect 1719 28033 1731 28036
rect 1673 28027 1731 28033
rect 1486 27928 1492 27940
rect 1447 27900 1492 27928
rect 1486 27888 1492 27900
rect 1544 27888 1550 27940
rect 2240 27937 2268 28036
rect 18230 28024 18236 28036
rect 18288 28064 18294 28076
rect 19352 28073 19380 28104
rect 19444 28104 20760 28132
rect 21269 28135 21327 28141
rect 19245 28067 19303 28073
rect 19245 28064 19257 28067
rect 18288 28036 19257 28064
rect 18288 28024 18294 28036
rect 19245 28033 19257 28036
rect 19291 28033 19303 28067
rect 19245 28027 19303 28033
rect 19337 28067 19395 28073
rect 19337 28033 19349 28067
rect 19383 28033 19395 28067
rect 19337 28027 19395 28033
rect 15286 27956 15292 28008
rect 15344 27996 15350 28008
rect 19444 27996 19472 28104
rect 21269 28101 21281 28135
rect 21315 28132 21327 28135
rect 23474 28132 23480 28144
rect 21315 28104 23480 28132
rect 21315 28101 21327 28104
rect 21269 28095 21327 28101
rect 19521 28067 19579 28073
rect 19521 28033 19533 28067
rect 19567 28033 19579 28067
rect 19702 28064 19708 28076
rect 19663 28036 19708 28064
rect 19521 28027 19579 28033
rect 15344 27968 19472 27996
rect 19536 27996 19564 28027
rect 19702 28024 19708 28036
rect 19760 28024 19766 28076
rect 19886 28024 19892 28076
rect 19944 28064 19950 28076
rect 20625 28067 20683 28073
rect 20625 28064 20637 28067
rect 19944 28036 20637 28064
rect 19944 28024 19950 28036
rect 20625 28033 20637 28036
rect 20671 28033 20683 28067
rect 22278 28064 22284 28076
rect 22239 28036 22284 28064
rect 20625 28027 20683 28033
rect 22278 28024 22284 28036
rect 22336 28024 22342 28076
rect 22848 28073 22876 28104
rect 23474 28092 23480 28104
rect 23532 28092 23538 28144
rect 25133 28135 25191 28141
rect 25133 28101 25145 28135
rect 25179 28132 25191 28135
rect 26050 28132 26056 28144
rect 25179 28104 26056 28132
rect 25179 28101 25191 28104
rect 25133 28095 25191 28101
rect 26050 28092 26056 28104
rect 26108 28092 26114 28144
rect 31481 28135 31539 28141
rect 31481 28132 31493 28135
rect 27632 28104 28672 28132
rect 22833 28067 22891 28073
rect 22833 28033 22845 28067
rect 22879 28033 22891 28067
rect 22833 28027 22891 28033
rect 23017 28067 23075 28073
rect 23017 28033 23029 28067
rect 23063 28064 23075 28067
rect 23661 28067 23719 28073
rect 23661 28064 23673 28067
rect 23063 28036 23673 28064
rect 23063 28033 23075 28036
rect 23017 28027 23075 28033
rect 23661 28033 23673 28036
rect 23707 28033 23719 28067
rect 23661 28027 23719 28033
rect 23845 28067 23903 28073
rect 23845 28033 23857 28067
rect 23891 28064 23903 28067
rect 24762 28064 24768 28076
rect 23891 28036 24768 28064
rect 23891 28033 23903 28036
rect 23845 28027 23903 28033
rect 20165 27999 20223 28005
rect 20165 27996 20177 27999
rect 19536 27968 20177 27996
rect 15344 27956 15350 27968
rect 20165 27965 20177 27968
rect 20211 27965 20223 27999
rect 22296 27996 22324 28024
rect 23032 27996 23060 28027
rect 24762 28024 24768 28036
rect 24820 28064 24826 28076
rect 24857 28067 24915 28073
rect 24857 28064 24869 28067
rect 24820 28036 24869 28064
rect 24820 28024 24826 28036
rect 24857 28033 24869 28036
rect 24903 28033 24915 28067
rect 25958 28064 25964 28076
rect 25919 28036 25964 28064
rect 24857 28027 24915 28033
rect 25958 28024 25964 28036
rect 26016 28024 26022 28076
rect 26237 28067 26295 28073
rect 26237 28033 26249 28067
rect 26283 28064 26295 28067
rect 26510 28064 26516 28076
rect 26283 28036 26516 28064
rect 26283 28033 26295 28036
rect 26237 28027 26295 28033
rect 26510 28024 26516 28036
rect 26568 28024 26574 28076
rect 27632 28073 27660 28104
rect 28644 28073 28672 28104
rect 30852 28104 31493 28132
rect 30852 28076 30880 28104
rect 31481 28101 31493 28104
rect 31527 28132 31539 28135
rect 31938 28132 31944 28144
rect 31527 28104 31944 28132
rect 31527 28101 31539 28104
rect 31481 28095 31539 28101
rect 31938 28092 31944 28104
rect 31996 28092 32002 28144
rect 32122 28092 32128 28144
rect 32180 28132 32186 28144
rect 33980 28141 34008 28172
rect 34057 28169 34069 28203
rect 34103 28200 34115 28203
rect 34606 28200 34612 28212
rect 34103 28172 34612 28200
rect 34103 28169 34115 28172
rect 34057 28163 34115 28169
rect 34606 28160 34612 28172
rect 34664 28160 34670 28212
rect 35161 28203 35219 28209
rect 35161 28169 35173 28203
rect 35207 28200 35219 28203
rect 37550 28200 37556 28212
rect 35207 28172 37556 28200
rect 35207 28169 35219 28172
rect 35161 28163 35219 28169
rect 33781 28135 33839 28141
rect 33781 28132 33793 28135
rect 32180 28104 33793 28132
rect 32180 28092 32186 28104
rect 33781 28101 33793 28104
rect 33827 28101 33839 28135
rect 33781 28095 33839 28101
rect 33965 28135 34023 28141
rect 33965 28101 33977 28135
rect 34011 28101 34023 28135
rect 34514 28132 34520 28144
rect 34427 28104 34520 28132
rect 33965 28095 34023 28101
rect 34514 28092 34520 28104
rect 34572 28132 34578 28144
rect 35176 28132 35204 28163
rect 37550 28160 37556 28172
rect 37608 28160 37614 28212
rect 34572 28104 35204 28132
rect 34572 28092 34578 28104
rect 27617 28067 27675 28073
rect 27617 28033 27629 28067
rect 27663 28033 27675 28067
rect 28445 28067 28503 28073
rect 28445 28064 28457 28067
rect 27617 28027 27675 28033
rect 27724 28036 28457 28064
rect 27724 28008 27752 28036
rect 28445 28033 28457 28036
rect 28491 28033 28503 28067
rect 28445 28027 28503 28033
rect 28629 28067 28687 28073
rect 28629 28033 28641 28067
rect 28675 28064 28687 28067
rect 28810 28064 28816 28076
rect 28675 28036 28816 28064
rect 28675 28033 28687 28036
rect 28629 28027 28687 28033
rect 28810 28024 28816 28036
rect 28868 28024 28874 28076
rect 30190 28064 30196 28076
rect 30151 28036 30196 28064
rect 30190 28024 30196 28036
rect 30248 28024 30254 28076
rect 30374 28064 30380 28076
rect 30335 28036 30380 28064
rect 30374 28024 30380 28036
rect 30432 28024 30438 28076
rect 30834 28064 30840 28076
rect 30795 28036 30840 28064
rect 30834 28024 30840 28036
rect 30892 28024 30898 28076
rect 31018 28064 31024 28076
rect 30979 28036 31024 28064
rect 31018 28024 31024 28036
rect 31076 28024 31082 28076
rect 32858 28064 32864 28076
rect 32819 28036 32864 28064
rect 32858 28024 32864 28036
rect 32916 28024 32922 28076
rect 33229 28067 33287 28073
rect 33229 28033 33241 28067
rect 33275 28064 33287 28067
rect 33502 28064 33508 28076
rect 33275 28036 33508 28064
rect 33275 28033 33287 28036
rect 33229 28027 33287 28033
rect 33502 28024 33508 28036
rect 33560 28024 33566 28076
rect 34054 28024 34060 28076
rect 34112 28064 34118 28076
rect 34112 28036 34157 28064
rect 34112 28024 34118 28036
rect 23474 27996 23480 28008
rect 22296 27968 23060 27996
rect 23435 27968 23480 27996
rect 20165 27959 20223 27965
rect 23474 27956 23480 27968
rect 23532 27956 23538 28008
rect 25133 27999 25191 28005
rect 25133 27965 25145 27999
rect 25179 27996 25191 27999
rect 25222 27996 25228 28008
rect 25179 27968 25228 27996
rect 25179 27965 25191 27968
rect 25133 27959 25191 27965
rect 25222 27956 25228 27968
rect 25280 27956 25286 28008
rect 27706 27996 27712 28008
rect 27667 27968 27712 27996
rect 27706 27956 27712 27968
rect 27764 27956 27770 28008
rect 29733 27999 29791 28005
rect 29733 27965 29745 27999
rect 29779 27996 29791 27999
rect 31036 27996 31064 28024
rect 29779 27968 31064 27996
rect 29779 27965 29791 27968
rect 29733 27959 29791 27965
rect 2225 27931 2283 27937
rect 2225 27897 2237 27931
rect 2271 27928 2283 27931
rect 17773 27931 17831 27937
rect 2271 27900 6914 27928
rect 2271 27897 2283 27900
rect 2225 27891 2283 27897
rect 6886 27860 6914 27900
rect 17773 27897 17785 27931
rect 17819 27928 17831 27931
rect 17954 27928 17960 27940
rect 17819 27900 17960 27928
rect 17819 27897 17831 27900
rect 17773 27891 17831 27897
rect 17954 27888 17960 27900
rect 18012 27928 18018 27940
rect 19242 27928 19248 27940
rect 18012 27900 19248 27928
rect 18012 27888 18018 27900
rect 19242 27888 19248 27900
rect 19300 27888 19306 27940
rect 19426 27928 19432 27940
rect 19387 27900 19432 27928
rect 19426 27888 19432 27900
rect 19484 27888 19490 27940
rect 24397 27931 24455 27937
rect 24397 27897 24409 27931
rect 24443 27928 24455 27931
rect 24854 27928 24860 27940
rect 24443 27900 24860 27928
rect 24443 27897 24455 27900
rect 24397 27891 24455 27897
rect 24854 27888 24860 27900
rect 24912 27928 24918 27940
rect 25498 27928 25504 27940
rect 24912 27900 25504 27928
rect 24912 27888 24918 27900
rect 25498 27888 25504 27900
rect 25556 27888 25562 27940
rect 26237 27931 26295 27937
rect 26237 27897 26249 27931
rect 26283 27928 26295 27931
rect 26786 27928 26792 27940
rect 26283 27900 26792 27928
rect 26283 27897 26295 27900
rect 26237 27891 26295 27897
rect 26786 27888 26792 27900
rect 26844 27888 26850 27940
rect 18598 27860 18604 27872
rect 6886 27832 18604 27860
rect 18598 27820 18604 27832
rect 18656 27820 18662 27872
rect 19334 27820 19340 27872
rect 19392 27860 19398 27872
rect 20349 27863 20407 27869
rect 20349 27860 20361 27863
rect 19392 27832 20361 27860
rect 19392 27820 19398 27832
rect 20349 27829 20361 27832
rect 20395 27829 20407 27863
rect 20349 27823 20407 27829
rect 23017 27863 23075 27869
rect 23017 27829 23029 27863
rect 23063 27860 23075 27863
rect 23566 27860 23572 27872
rect 23063 27832 23572 27860
rect 23063 27829 23075 27832
rect 23017 27823 23075 27829
rect 23566 27820 23572 27832
rect 23624 27820 23630 27872
rect 24946 27860 24952 27872
rect 24907 27832 24952 27860
rect 24946 27820 24952 27832
rect 25004 27820 25010 27872
rect 28810 27820 28816 27872
rect 28868 27860 28874 27872
rect 29089 27863 29147 27869
rect 29089 27860 29101 27863
rect 28868 27832 29101 27860
rect 28868 27820 28874 27832
rect 29089 27829 29101 27832
rect 29135 27829 29147 27863
rect 29089 27823 29147 27829
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 19426 27616 19432 27668
rect 19484 27656 19490 27668
rect 19797 27659 19855 27665
rect 19797 27656 19809 27659
rect 19484 27628 19809 27656
rect 19484 27616 19490 27628
rect 19797 27625 19809 27628
rect 19843 27656 19855 27659
rect 20070 27656 20076 27668
rect 19843 27628 20076 27656
rect 19843 27625 19855 27628
rect 19797 27619 19855 27625
rect 20070 27616 20076 27628
rect 20128 27616 20134 27668
rect 21821 27659 21879 27665
rect 21821 27625 21833 27659
rect 21867 27656 21879 27659
rect 22094 27656 22100 27668
rect 21867 27628 22100 27656
rect 21867 27625 21879 27628
rect 21821 27619 21879 27625
rect 22094 27616 22100 27628
rect 22152 27616 22158 27668
rect 26050 27616 26056 27668
rect 26108 27656 26114 27668
rect 26237 27659 26295 27665
rect 26237 27656 26249 27659
rect 26108 27628 26249 27656
rect 26108 27616 26114 27628
rect 26237 27625 26249 27628
rect 26283 27625 26295 27659
rect 26237 27619 26295 27625
rect 26421 27659 26479 27665
rect 26421 27625 26433 27659
rect 26467 27656 26479 27659
rect 27154 27656 27160 27668
rect 26467 27628 27160 27656
rect 26467 27625 26479 27628
rect 26421 27619 26479 27625
rect 27154 27616 27160 27628
rect 27212 27616 27218 27668
rect 27982 27616 27988 27668
rect 28040 27656 28046 27668
rect 28077 27659 28135 27665
rect 28077 27656 28089 27659
rect 28040 27628 28089 27656
rect 28040 27616 28046 27628
rect 28077 27625 28089 27628
rect 28123 27625 28135 27659
rect 28077 27619 28135 27625
rect 30561 27659 30619 27665
rect 30561 27625 30573 27659
rect 30607 27656 30619 27659
rect 30834 27656 30840 27668
rect 30607 27628 30840 27656
rect 30607 27625 30619 27628
rect 30561 27619 30619 27625
rect 30834 27616 30840 27628
rect 30892 27616 30898 27668
rect 32217 27659 32275 27665
rect 32217 27625 32229 27659
rect 32263 27656 32275 27659
rect 32858 27656 32864 27668
rect 32263 27628 32864 27656
rect 32263 27625 32275 27628
rect 32217 27619 32275 27625
rect 32858 27616 32864 27628
rect 32916 27616 32922 27668
rect 18598 27588 18604 27600
rect 18559 27560 18604 27588
rect 18598 27548 18604 27560
rect 18656 27548 18662 27600
rect 20990 27588 20996 27600
rect 20951 27560 20996 27588
rect 20990 27548 20996 27560
rect 21048 27548 21054 27600
rect 22005 27591 22063 27597
rect 22005 27557 22017 27591
rect 22051 27588 22063 27591
rect 22186 27588 22192 27600
rect 22051 27560 22192 27588
rect 22051 27557 22063 27560
rect 22005 27551 22063 27557
rect 22186 27548 22192 27560
rect 22244 27548 22250 27600
rect 23109 27591 23167 27597
rect 23109 27557 23121 27591
rect 23155 27588 23167 27591
rect 24946 27588 24952 27600
rect 23155 27560 24952 27588
rect 23155 27557 23167 27560
rect 23109 27551 23167 27557
rect 24946 27548 24952 27560
rect 25004 27548 25010 27600
rect 33502 27588 33508 27600
rect 33463 27560 33508 27588
rect 33502 27548 33508 27560
rect 33560 27548 33566 27600
rect 33594 27548 33600 27600
rect 33652 27588 33658 27600
rect 46382 27588 46388 27600
rect 33652 27560 46388 27588
rect 33652 27548 33658 27560
rect 46382 27548 46388 27560
rect 46440 27548 46446 27600
rect 22204 27520 22232 27548
rect 27525 27523 27583 27529
rect 22204 27492 22784 27520
rect 19702 27452 19708 27464
rect 19615 27424 19708 27452
rect 19702 27412 19708 27424
rect 19760 27412 19766 27464
rect 19886 27452 19892 27464
rect 19847 27424 19892 27452
rect 19886 27412 19892 27424
rect 19944 27412 19950 27464
rect 21542 27452 21548 27464
rect 21503 27424 21548 27452
rect 21542 27412 21548 27424
rect 21600 27412 21606 27464
rect 22278 27412 22284 27464
rect 22336 27452 22342 27464
rect 22756 27461 22784 27492
rect 27525 27489 27537 27523
rect 27571 27520 27583 27523
rect 27985 27523 28043 27529
rect 27985 27520 27997 27523
rect 27571 27492 27997 27520
rect 27571 27489 27583 27492
rect 27525 27483 27583 27489
rect 27985 27489 27997 27492
rect 28031 27489 28043 27523
rect 27985 27483 28043 27489
rect 33321 27523 33379 27529
rect 33321 27489 33333 27523
rect 33367 27520 33379 27523
rect 34790 27520 34796 27532
rect 33367 27492 34796 27520
rect 33367 27489 33379 27492
rect 33321 27483 33379 27489
rect 34790 27480 34796 27492
rect 34848 27480 34854 27532
rect 48130 27520 48136 27532
rect 48091 27492 48136 27520
rect 48130 27480 48136 27492
rect 48188 27480 48194 27532
rect 22465 27455 22523 27461
rect 22465 27452 22477 27455
rect 22336 27424 22477 27452
rect 22336 27412 22342 27424
rect 22465 27421 22477 27424
rect 22511 27421 22523 27455
rect 22465 27415 22523 27421
rect 22649 27455 22707 27461
rect 22649 27421 22661 27455
rect 22695 27421 22707 27455
rect 22649 27415 22707 27421
rect 22741 27455 22799 27461
rect 22741 27421 22753 27455
rect 22787 27421 22799 27455
rect 22741 27415 22799 27421
rect 22833 27455 22891 27461
rect 22833 27421 22845 27455
rect 22879 27452 22891 27455
rect 22922 27452 22928 27464
rect 22879 27424 22928 27452
rect 22879 27421 22891 27424
rect 22833 27415 22891 27421
rect 19720 27384 19748 27412
rect 20162 27384 20168 27396
rect 19720 27356 20168 27384
rect 20162 27344 20168 27356
rect 20220 27344 20226 27396
rect 22664 27384 22692 27415
rect 22922 27412 22928 27424
rect 22980 27412 22986 27464
rect 23566 27452 23572 27464
rect 23527 27424 23572 27452
rect 23566 27412 23572 27424
rect 23624 27412 23630 27464
rect 23753 27455 23811 27461
rect 23753 27421 23765 27455
rect 23799 27452 23811 27455
rect 24762 27452 24768 27464
rect 23799 27424 24768 27452
rect 23799 27421 23811 27424
rect 23753 27415 23811 27421
rect 24762 27412 24768 27424
rect 24820 27412 24826 27464
rect 25130 27452 25136 27464
rect 25091 27424 25136 27452
rect 25130 27412 25136 27424
rect 25188 27412 25194 27464
rect 25317 27455 25375 27461
rect 25317 27421 25329 27455
rect 25363 27452 25375 27455
rect 26234 27452 26240 27464
rect 25363 27424 26240 27452
rect 25363 27421 25375 27424
rect 25317 27415 25375 27421
rect 26234 27412 26240 27424
rect 26292 27412 26298 27464
rect 27065 27455 27123 27461
rect 27065 27421 27077 27455
rect 27111 27421 27123 27455
rect 27065 27415 27123 27421
rect 23014 27384 23020 27396
rect 22664 27356 23020 27384
rect 23014 27344 23020 27356
rect 23072 27384 23078 27396
rect 23661 27387 23719 27393
rect 23661 27384 23673 27387
rect 23072 27356 23673 27384
rect 23072 27344 23078 27356
rect 23661 27353 23673 27356
rect 23707 27353 23719 27387
rect 23661 27347 23719 27353
rect 24489 27387 24547 27393
rect 24489 27353 24501 27387
rect 24535 27384 24547 27387
rect 25148 27384 25176 27412
rect 24535 27356 25176 27384
rect 26053 27387 26111 27393
rect 24535 27353 24547 27356
rect 24489 27347 24547 27353
rect 26053 27353 26065 27387
rect 26099 27384 26111 27387
rect 26510 27384 26516 27396
rect 26099 27356 26516 27384
rect 26099 27353 26111 27356
rect 26053 27347 26111 27353
rect 26510 27344 26516 27356
rect 26568 27344 26574 27396
rect 27080 27384 27108 27415
rect 27154 27412 27160 27464
rect 27212 27452 27218 27464
rect 27341 27455 27399 27461
rect 27341 27452 27353 27455
rect 27212 27424 27353 27452
rect 27212 27412 27218 27424
rect 27341 27421 27353 27424
rect 27387 27421 27399 27455
rect 27341 27415 27399 27421
rect 28169 27455 28227 27461
rect 28169 27421 28181 27455
rect 28215 27421 28227 27455
rect 28169 27415 28227 27421
rect 28261 27455 28319 27461
rect 28261 27421 28273 27455
rect 28307 27452 28319 27455
rect 28721 27455 28779 27461
rect 28721 27452 28733 27455
rect 28307 27424 28733 27452
rect 28307 27421 28319 27424
rect 28261 27415 28319 27421
rect 28721 27421 28733 27424
rect 28767 27452 28779 27455
rect 28994 27452 29000 27464
rect 28767 27424 29000 27452
rect 28767 27421 28779 27424
rect 28721 27415 28779 27421
rect 28184 27384 28212 27415
rect 27080 27356 28212 27384
rect 27356 27328 27384 27356
rect 20530 27316 20536 27328
rect 20491 27288 20536 27316
rect 20530 27276 20536 27288
rect 20588 27276 20594 27328
rect 24946 27316 24952 27328
rect 24907 27288 24952 27316
rect 24946 27276 24952 27288
rect 25004 27276 25010 27328
rect 25958 27276 25964 27328
rect 26016 27316 26022 27328
rect 26253 27319 26311 27325
rect 26253 27316 26265 27319
rect 26016 27288 26265 27316
rect 26016 27276 26022 27288
rect 26253 27285 26265 27288
rect 26299 27285 26311 27319
rect 27154 27316 27160 27328
rect 27115 27288 27160 27316
rect 26253 27279 26311 27285
rect 27154 27276 27160 27288
rect 27212 27276 27218 27328
rect 27338 27276 27344 27328
rect 27396 27276 27402 27328
rect 27430 27276 27436 27328
rect 27488 27316 27494 27328
rect 28276 27316 28304 27415
rect 28994 27412 29000 27424
rect 29052 27452 29058 27464
rect 29549 27455 29607 27461
rect 29549 27452 29561 27455
rect 29052 27424 29561 27452
rect 29052 27412 29058 27424
rect 29549 27421 29561 27424
rect 29595 27421 29607 27455
rect 29549 27415 29607 27421
rect 30834 27412 30840 27464
rect 30892 27452 30898 27464
rect 31110 27452 31116 27464
rect 30892 27424 31116 27452
rect 30892 27412 30898 27424
rect 31110 27412 31116 27424
rect 31168 27452 31174 27464
rect 31205 27455 31263 27461
rect 31205 27452 31217 27455
rect 31168 27424 31217 27452
rect 31168 27412 31174 27424
rect 31205 27421 31217 27424
rect 31251 27421 31263 27455
rect 31205 27415 31263 27421
rect 31389 27455 31447 27461
rect 31389 27421 31401 27455
rect 31435 27452 31447 27455
rect 32122 27452 32128 27464
rect 31435 27424 32128 27452
rect 31435 27421 31447 27424
rect 31389 27415 31447 27421
rect 32122 27412 32128 27424
rect 32180 27412 32186 27464
rect 32309 27455 32367 27461
rect 32309 27421 32321 27455
rect 32355 27452 32367 27455
rect 32490 27452 32496 27464
rect 32355 27424 32496 27452
rect 32355 27421 32367 27424
rect 32309 27415 32367 27421
rect 30650 27344 30656 27396
rect 30708 27384 30714 27396
rect 31018 27384 31024 27396
rect 30708 27356 31024 27384
rect 30708 27344 30714 27356
rect 31018 27344 31024 27356
rect 31076 27344 31082 27396
rect 32030 27344 32036 27396
rect 32088 27384 32094 27396
rect 32324 27384 32352 27415
rect 32490 27412 32496 27424
rect 32548 27412 32554 27464
rect 33229 27455 33287 27461
rect 33229 27421 33241 27455
rect 33275 27452 33287 27455
rect 34054 27452 34060 27464
rect 33275 27424 34060 27452
rect 33275 27421 33287 27424
rect 33229 27415 33287 27421
rect 34054 27412 34060 27424
rect 34112 27412 34118 27464
rect 36538 27412 36544 27464
rect 36596 27452 36602 27464
rect 47857 27455 47915 27461
rect 47857 27452 47869 27455
rect 36596 27424 47869 27452
rect 36596 27412 36602 27424
rect 47857 27421 47869 27424
rect 47903 27421 47915 27455
rect 47857 27415 47915 27421
rect 32088 27356 32352 27384
rect 32088 27344 32094 27356
rect 27488 27288 28304 27316
rect 27488 27276 27494 27288
rect 32306 27276 32312 27328
rect 32364 27316 32370 27328
rect 32861 27319 32919 27325
rect 32861 27316 32873 27319
rect 32364 27288 32873 27316
rect 32364 27276 32370 27288
rect 32861 27285 32873 27288
rect 32907 27285 32919 27319
rect 33962 27316 33968 27328
rect 33923 27288 33968 27316
rect 32861 27279 32919 27285
rect 33962 27276 33968 27288
rect 34020 27276 34026 27328
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 18598 27072 18604 27124
rect 18656 27112 18662 27124
rect 18785 27115 18843 27121
rect 18785 27112 18797 27115
rect 18656 27084 18797 27112
rect 18656 27072 18662 27084
rect 18785 27081 18797 27084
rect 18831 27081 18843 27115
rect 18785 27075 18843 27081
rect 19978 27072 19984 27124
rect 20036 27112 20042 27124
rect 20165 27115 20223 27121
rect 20165 27112 20177 27115
rect 20036 27084 20177 27112
rect 20036 27072 20042 27084
rect 20165 27081 20177 27084
rect 20211 27081 20223 27115
rect 21818 27112 21824 27124
rect 20165 27075 20223 27081
rect 21100 27084 21824 27112
rect 19610 27004 19616 27056
rect 19668 27044 19674 27056
rect 19705 27047 19763 27053
rect 19705 27044 19717 27047
rect 19668 27016 19717 27044
rect 19668 27004 19674 27016
rect 19705 27013 19717 27016
rect 19751 27044 19763 27047
rect 20346 27044 20352 27056
rect 19751 27016 20352 27044
rect 19751 27013 19763 27016
rect 19705 27007 19763 27013
rect 20346 27004 20352 27016
rect 20404 27004 20410 27056
rect 21100 26988 21128 27084
rect 21818 27072 21824 27084
rect 21876 27072 21882 27124
rect 21913 27115 21971 27121
rect 21913 27081 21925 27115
rect 21959 27112 21971 27115
rect 22002 27112 22008 27124
rect 21959 27084 22008 27112
rect 21959 27081 21971 27084
rect 21913 27075 21971 27081
rect 22002 27072 22008 27084
rect 22060 27072 22066 27124
rect 23385 27115 23443 27121
rect 23385 27081 23397 27115
rect 23431 27112 23443 27115
rect 24578 27112 24584 27124
rect 23431 27084 24584 27112
rect 23431 27081 23443 27084
rect 23385 27075 23443 27081
rect 24578 27072 24584 27084
rect 24636 27072 24642 27124
rect 24762 27072 24768 27124
rect 24820 27112 24826 27124
rect 24820 27084 25820 27112
rect 24820 27072 24826 27084
rect 21177 27047 21235 27053
rect 21177 27013 21189 27047
rect 21223 27044 21235 27047
rect 21542 27044 21548 27056
rect 21223 27016 21548 27044
rect 21223 27013 21235 27016
rect 21177 27007 21235 27013
rect 21542 27004 21548 27016
rect 21600 27044 21606 27056
rect 24121 27047 24179 27053
rect 21600 27016 22140 27044
rect 21600 27004 21606 27016
rect 20530 26976 20536 26988
rect 20491 26948 20536 26976
rect 20530 26936 20536 26948
rect 20588 26936 20594 26988
rect 21082 26976 21088 26988
rect 20995 26948 21088 26976
rect 21082 26936 21088 26948
rect 21140 26936 21146 26988
rect 22112 26985 22140 27016
rect 24121 27013 24133 27047
rect 24167 27044 24179 27047
rect 25222 27044 25228 27056
rect 24167 27016 25228 27044
rect 24167 27013 24179 27016
rect 24121 27007 24179 27013
rect 25222 27004 25228 27016
rect 25280 27044 25286 27056
rect 25280 27016 25728 27044
rect 25280 27004 25286 27016
rect 21269 26979 21327 26985
rect 21269 26945 21281 26979
rect 21315 26945 21327 26979
rect 21269 26939 21327 26945
rect 22097 26979 22155 26985
rect 22097 26945 22109 26979
rect 22143 26945 22155 26979
rect 23014 26976 23020 26988
rect 22975 26948 23020 26976
rect 22097 26939 22155 26945
rect 21284 26840 21312 26939
rect 23014 26936 23020 26948
rect 23072 26936 23078 26988
rect 24026 26976 24032 26988
rect 23987 26948 24032 26976
rect 24026 26936 24032 26948
rect 24084 26936 24090 26988
rect 24213 26979 24271 26985
rect 24213 26945 24225 26979
rect 24259 26945 24271 26979
rect 24213 26939 24271 26945
rect 22278 26908 22284 26920
rect 22239 26880 22284 26908
rect 22278 26868 22284 26880
rect 22336 26868 22342 26920
rect 23106 26908 23112 26920
rect 23067 26880 23112 26908
rect 23106 26868 23112 26880
rect 23164 26868 23170 26920
rect 24228 26908 24256 26939
rect 24762 26936 24768 26988
rect 24820 26976 24826 26988
rect 24857 26979 24915 26985
rect 24857 26976 24869 26979
rect 24820 26948 24869 26976
rect 24820 26936 24826 26948
rect 24857 26945 24869 26948
rect 24903 26945 24915 26979
rect 24857 26939 24915 26945
rect 24946 26936 24952 26988
rect 25004 26936 25010 26988
rect 25038 26936 25044 26988
rect 25096 26976 25102 26988
rect 25700 26985 25728 27016
rect 25792 26985 25820 27084
rect 25958 27072 25964 27124
rect 26016 27112 26022 27124
rect 26053 27115 26111 27121
rect 26053 27112 26065 27115
rect 26016 27084 26065 27112
rect 26016 27072 26022 27084
rect 26053 27081 26065 27084
rect 26099 27081 26111 27115
rect 26053 27075 26111 27081
rect 26326 27072 26332 27124
rect 26384 27112 26390 27124
rect 27065 27115 27123 27121
rect 27065 27112 27077 27115
rect 26384 27084 27077 27112
rect 26384 27072 26390 27084
rect 27065 27081 27077 27084
rect 27111 27081 27123 27115
rect 27065 27075 27123 27081
rect 30466 27072 30472 27124
rect 30524 27072 30530 27124
rect 31113 27115 31171 27121
rect 31113 27081 31125 27115
rect 31159 27112 31171 27115
rect 32030 27112 32036 27124
rect 31159 27084 32036 27112
rect 31159 27081 31171 27084
rect 31113 27075 31171 27081
rect 32030 27072 32036 27084
rect 32088 27072 32094 27124
rect 32306 27112 32312 27124
rect 32267 27084 32312 27112
rect 32306 27072 32312 27084
rect 32364 27072 32370 27124
rect 48130 27112 48136 27124
rect 48091 27084 48136 27112
rect 48130 27072 48136 27084
rect 48188 27072 48194 27124
rect 30484 27044 30512 27072
rect 29288 27016 30512 27044
rect 25133 26979 25191 26985
rect 25133 26976 25145 26979
rect 25096 26948 25145 26976
rect 25096 26936 25102 26948
rect 25133 26945 25145 26948
rect 25179 26945 25191 26979
rect 25133 26939 25191 26945
rect 25685 26979 25743 26985
rect 25685 26945 25697 26979
rect 25731 26945 25743 26979
rect 25685 26939 25743 26945
rect 25777 26979 25835 26985
rect 25777 26945 25789 26979
rect 25823 26945 25835 26979
rect 25777 26939 25835 26945
rect 27154 26936 27160 26988
rect 27212 26976 27218 26988
rect 27430 26976 27436 26988
rect 27212 26948 27436 26976
rect 27212 26936 27218 26948
rect 27430 26936 27436 26948
rect 27488 26936 27494 26988
rect 28442 26976 28448 26988
rect 28403 26948 28448 26976
rect 28442 26936 28448 26948
rect 28500 26936 28506 26988
rect 24964 26908 24992 26936
rect 27338 26908 27344 26920
rect 24228 26880 25084 26908
rect 27299 26880 27344 26908
rect 22462 26840 22468 26852
rect 21284 26812 22468 26840
rect 22462 26800 22468 26812
rect 22520 26800 22526 26852
rect 24946 26840 24952 26852
rect 24907 26812 24952 26840
rect 24946 26800 24952 26812
rect 25004 26800 25010 26852
rect 25056 26849 25084 26880
rect 27338 26868 27344 26880
rect 27396 26868 27402 26920
rect 28537 26911 28595 26917
rect 28537 26877 28549 26911
rect 28583 26908 28595 26911
rect 29288 26908 29316 27016
rect 31202 27004 31208 27056
rect 31260 27044 31266 27056
rect 32766 27044 32772 27056
rect 31260 27016 32772 27044
rect 31260 27004 31266 27016
rect 29457 26979 29515 26985
rect 29457 26945 29469 26979
rect 29503 26976 29515 26979
rect 29822 26976 29828 26988
rect 29503 26948 29828 26976
rect 29503 26945 29515 26948
rect 29457 26939 29515 26945
rect 29822 26936 29828 26948
rect 29880 26936 29886 26988
rect 30282 26976 30288 26988
rect 30243 26948 30288 26976
rect 30282 26936 30288 26948
rect 30340 26936 30346 26988
rect 30466 26976 30472 26988
rect 30427 26948 30472 26976
rect 30466 26936 30472 26948
rect 30524 26936 30530 26988
rect 30650 26936 30656 26988
rect 30708 26976 30714 26988
rect 30929 26979 30987 26985
rect 30929 26976 30941 26979
rect 30708 26948 30941 26976
rect 30708 26936 30714 26948
rect 30929 26945 30941 26948
rect 30975 26945 30987 26979
rect 31110 26976 31116 26988
rect 31071 26948 31116 26976
rect 30929 26939 30987 26945
rect 31110 26936 31116 26948
rect 31168 26936 31174 26988
rect 32324 26985 32352 27016
rect 32766 27004 32772 27016
rect 32824 27004 32830 27056
rect 34054 27004 34060 27056
rect 34112 27044 34118 27056
rect 34149 27047 34207 27053
rect 34149 27044 34161 27047
rect 34112 27016 34161 27044
rect 34112 27004 34118 27016
rect 34149 27013 34161 27016
rect 34195 27013 34207 27047
rect 34149 27007 34207 27013
rect 32309 26979 32367 26985
rect 32309 26945 32321 26979
rect 32355 26945 32367 26979
rect 32309 26939 32367 26945
rect 32493 26979 32551 26985
rect 32493 26945 32505 26979
rect 32539 26976 32551 26979
rect 33042 26976 33048 26988
rect 32539 26948 33048 26976
rect 32539 26945 32551 26948
rect 32493 26939 32551 26945
rect 28583 26880 29316 26908
rect 29365 26911 29423 26917
rect 28583 26877 28595 26880
rect 28537 26871 28595 26877
rect 29365 26877 29377 26911
rect 29411 26877 29423 26911
rect 29365 26871 29423 26877
rect 25041 26843 25099 26849
rect 25041 26809 25053 26843
rect 25087 26809 25099 26843
rect 25041 26803 25099 26809
rect 28813 26843 28871 26849
rect 28813 26809 28825 26843
rect 28859 26840 28871 26843
rect 29380 26840 29408 26871
rect 32030 26868 32036 26920
rect 32088 26908 32094 26920
rect 32508 26908 32536 26939
rect 33042 26936 33048 26948
rect 33100 26976 33106 26988
rect 33100 26948 33258 26976
rect 33100 26936 33106 26948
rect 39574 26936 39580 26988
rect 39632 26936 39638 26988
rect 32088 26880 32536 26908
rect 32088 26868 32094 26880
rect 32766 26868 32772 26920
rect 32824 26908 32830 26920
rect 33321 26911 33379 26917
rect 33321 26908 33333 26911
rect 32824 26880 33333 26908
rect 32824 26868 32830 26880
rect 33321 26877 33333 26880
rect 33367 26908 33379 26911
rect 33367 26880 34744 26908
rect 33367 26877 33379 26880
rect 33321 26871 33379 26877
rect 28859 26812 29408 26840
rect 29825 26843 29883 26849
rect 28859 26809 28871 26812
rect 28813 26803 28871 26809
rect 29825 26809 29837 26843
rect 29871 26840 29883 26843
rect 30098 26840 30104 26852
rect 29871 26812 30104 26840
rect 29871 26809 29883 26812
rect 29825 26803 29883 26809
rect 30098 26800 30104 26812
rect 30156 26800 30162 26852
rect 24673 26775 24731 26781
rect 24673 26741 24685 26775
rect 24719 26772 24731 26775
rect 24854 26772 24860 26784
rect 24719 26744 24860 26772
rect 24719 26741 24731 26744
rect 24673 26735 24731 26741
rect 24854 26732 24860 26744
rect 24912 26732 24918 26784
rect 24964 26772 24992 26800
rect 25685 26775 25743 26781
rect 25685 26772 25697 26775
rect 24964 26744 25697 26772
rect 25685 26741 25697 26744
rect 25731 26741 25743 26775
rect 30374 26772 30380 26784
rect 30335 26744 30380 26772
rect 25685 26735 25743 26741
rect 30374 26732 30380 26744
rect 30432 26732 30438 26784
rect 34716 26781 34744 26880
rect 39592 26784 39620 26936
rect 34701 26775 34759 26781
rect 34701 26741 34713 26775
rect 34747 26772 34759 26775
rect 36354 26772 36360 26784
rect 34747 26744 36360 26772
rect 34747 26741 34759 26744
rect 34701 26735 34759 26741
rect 36354 26732 36360 26744
rect 36412 26732 36418 26784
rect 39574 26732 39580 26784
rect 39632 26732 39638 26784
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 19610 26568 19616 26580
rect 19571 26540 19616 26568
rect 19610 26528 19616 26540
rect 19668 26528 19674 26580
rect 20162 26568 20168 26580
rect 20123 26540 20168 26568
rect 20162 26528 20168 26540
rect 20220 26528 20226 26580
rect 20901 26571 20959 26577
rect 20901 26537 20913 26571
rect 20947 26568 20959 26571
rect 21082 26568 21088 26580
rect 20947 26540 21088 26568
rect 20947 26537 20959 26540
rect 20901 26531 20959 26537
rect 21082 26528 21088 26540
rect 21140 26528 21146 26580
rect 22186 26528 22192 26580
rect 22244 26568 22250 26580
rect 22925 26571 22983 26577
rect 22925 26568 22937 26571
rect 22244 26540 22937 26568
rect 22244 26528 22250 26540
rect 22925 26537 22937 26540
rect 22971 26537 22983 26571
rect 22925 26531 22983 26537
rect 23017 26571 23075 26577
rect 23017 26537 23029 26571
rect 23063 26568 23075 26571
rect 23106 26568 23112 26580
rect 23063 26540 23112 26568
rect 23063 26537 23075 26540
rect 23017 26531 23075 26537
rect 23106 26528 23112 26540
rect 23164 26528 23170 26580
rect 25038 26568 25044 26580
rect 24999 26540 25044 26568
rect 25038 26528 25044 26540
rect 25096 26528 25102 26580
rect 26510 26568 26516 26580
rect 26471 26540 26516 26568
rect 26510 26528 26516 26540
rect 26568 26528 26574 26580
rect 29822 26568 29828 26580
rect 29783 26540 29828 26568
rect 29822 26528 29828 26540
rect 29880 26528 29886 26580
rect 30650 26528 30656 26580
rect 30708 26568 30714 26580
rect 31941 26571 31999 26577
rect 31941 26568 31953 26571
rect 30708 26540 31953 26568
rect 30708 26528 30714 26540
rect 31941 26537 31953 26540
rect 31987 26537 31999 26571
rect 31941 26531 31999 26537
rect 33042 26528 33048 26580
rect 33100 26568 33106 26580
rect 33597 26571 33655 26577
rect 33597 26568 33609 26571
rect 33100 26540 33609 26568
rect 33100 26528 33106 26540
rect 33597 26537 33609 26540
rect 33643 26537 33655 26571
rect 33597 26531 33655 26537
rect 24026 26460 24032 26512
rect 24084 26500 24090 26512
rect 25869 26503 25927 26509
rect 25869 26500 25881 26503
rect 24084 26472 25881 26500
rect 24084 26460 24090 26472
rect 25869 26469 25881 26472
rect 25915 26469 25927 26503
rect 25869 26463 25927 26469
rect 27157 26503 27215 26509
rect 27157 26469 27169 26503
rect 27203 26500 27215 26503
rect 36538 26500 36544 26512
rect 27203 26472 36544 26500
rect 27203 26469 27215 26472
rect 27157 26463 27215 26469
rect 22278 26392 22284 26444
rect 22336 26432 22342 26444
rect 22373 26435 22431 26441
rect 22373 26432 22385 26435
rect 22336 26404 22385 26432
rect 22336 26392 22342 26404
rect 22373 26401 22385 26404
rect 22419 26432 22431 26435
rect 23109 26435 23167 26441
rect 23109 26432 23121 26435
rect 22419 26404 23121 26432
rect 22419 26401 22431 26404
rect 22373 26395 22431 26401
rect 23109 26401 23121 26404
rect 23155 26401 23167 26435
rect 27172 26432 27200 26463
rect 36538 26460 36544 26472
rect 36596 26460 36602 26512
rect 23109 26395 23167 26401
rect 25884 26404 27200 26432
rect 30101 26435 30159 26441
rect 19610 26324 19616 26376
rect 19668 26364 19674 26376
rect 20073 26367 20131 26373
rect 20073 26364 20085 26367
rect 19668 26336 20085 26364
rect 19668 26324 19674 26336
rect 20073 26333 20085 26336
rect 20119 26333 20131 26367
rect 20073 26327 20131 26333
rect 20257 26367 20315 26373
rect 20257 26333 20269 26367
rect 20303 26364 20315 26367
rect 20530 26364 20536 26376
rect 20303 26336 20536 26364
rect 20303 26333 20315 26336
rect 20257 26327 20315 26333
rect 20530 26324 20536 26336
rect 20588 26324 20594 26376
rect 21818 26324 21824 26376
rect 21876 26364 21882 26376
rect 22189 26367 22247 26373
rect 22189 26364 22201 26367
rect 21876 26336 22201 26364
rect 21876 26324 21882 26336
rect 22189 26333 22201 26336
rect 22235 26333 22247 26367
rect 22189 26327 22247 26333
rect 22833 26367 22891 26373
rect 22833 26333 22845 26367
rect 22879 26364 22891 26367
rect 22922 26364 22928 26376
rect 22879 26336 22928 26364
rect 22879 26333 22891 26336
rect 22833 26327 22891 26333
rect 22922 26324 22928 26336
rect 22980 26324 22986 26376
rect 25130 26324 25136 26376
rect 25188 26364 25194 26376
rect 25409 26367 25467 26373
rect 25409 26364 25421 26367
rect 25188 26336 25421 26364
rect 25188 26324 25194 26336
rect 25409 26333 25421 26336
rect 25455 26364 25467 26367
rect 25774 26364 25780 26376
rect 25455 26336 25780 26364
rect 25455 26333 25467 26336
rect 25409 26327 25467 26333
rect 25774 26324 25780 26336
rect 25832 26364 25838 26376
rect 25884 26373 25912 26404
rect 30101 26401 30113 26435
rect 30147 26432 30159 26435
rect 30282 26432 30288 26444
rect 30147 26404 30288 26432
rect 30147 26401 30159 26404
rect 30101 26395 30159 26401
rect 30282 26392 30288 26404
rect 30340 26432 30346 26444
rect 31113 26435 31171 26441
rect 31113 26432 31125 26435
rect 30340 26404 31125 26432
rect 30340 26392 30346 26404
rect 31113 26401 31125 26404
rect 31159 26401 31171 26435
rect 31570 26432 31576 26444
rect 31113 26395 31171 26401
rect 31496 26404 31576 26432
rect 25869 26367 25927 26373
rect 25869 26364 25881 26367
rect 25832 26336 25881 26364
rect 25832 26324 25838 26336
rect 25869 26333 25881 26336
rect 25915 26333 25927 26367
rect 25869 26327 25927 26333
rect 26053 26367 26111 26373
rect 26053 26333 26065 26367
rect 26099 26364 26111 26367
rect 26234 26364 26240 26376
rect 26099 26336 26240 26364
rect 26099 26333 26111 26336
rect 26053 26327 26111 26333
rect 1578 26256 1584 26308
rect 1636 26296 1642 26308
rect 1857 26299 1915 26305
rect 1857 26296 1869 26299
rect 1636 26268 1869 26296
rect 1636 26256 1642 26268
rect 1857 26265 1869 26268
rect 1903 26265 1915 26299
rect 1857 26259 1915 26265
rect 2041 26299 2099 26305
rect 2041 26265 2053 26299
rect 2087 26296 2099 26299
rect 10778 26296 10784 26308
rect 2087 26268 10784 26296
rect 2087 26265 2099 26268
rect 2041 26259 2099 26265
rect 10778 26256 10784 26268
rect 10836 26256 10842 26308
rect 21453 26299 21511 26305
rect 21453 26265 21465 26299
rect 21499 26296 21511 26299
rect 22005 26299 22063 26305
rect 22005 26296 22017 26299
rect 21499 26268 22017 26296
rect 21499 26265 21511 26268
rect 21453 26259 21511 26265
rect 22005 26265 22017 26268
rect 22051 26296 22063 26299
rect 22462 26296 22468 26308
rect 22051 26268 22468 26296
rect 22051 26265 22063 26268
rect 22005 26259 22063 26265
rect 22462 26256 22468 26268
rect 22520 26256 22526 26308
rect 24581 26299 24639 26305
rect 24581 26265 24593 26299
rect 24627 26296 24639 26299
rect 25225 26299 25283 26305
rect 25225 26296 25237 26299
rect 24627 26268 25237 26296
rect 24627 26265 24639 26268
rect 24581 26259 24639 26265
rect 25225 26265 25237 26268
rect 25271 26296 25283 26299
rect 26068 26296 26096 26327
rect 26234 26324 26240 26336
rect 26292 26324 26298 26376
rect 29822 26324 29828 26376
rect 29880 26364 29886 26376
rect 31496 26373 31524 26404
rect 31570 26392 31576 26404
rect 31628 26432 31634 26444
rect 33137 26435 33195 26441
rect 33137 26432 33149 26435
rect 31628 26404 33149 26432
rect 31628 26392 31634 26404
rect 33137 26401 33149 26404
rect 33183 26432 33195 26435
rect 33594 26432 33600 26444
rect 33183 26404 33600 26432
rect 33183 26401 33195 26404
rect 33137 26395 33195 26401
rect 33594 26392 33600 26404
rect 33652 26392 33658 26444
rect 30009 26367 30067 26373
rect 30009 26364 30021 26367
rect 29880 26336 30021 26364
rect 29880 26324 29886 26336
rect 30009 26333 30021 26336
rect 30055 26333 30067 26367
rect 30009 26327 30067 26333
rect 31481 26367 31539 26373
rect 31481 26333 31493 26367
rect 31527 26333 31539 26367
rect 32585 26367 32643 26373
rect 32585 26364 32597 26367
rect 31481 26327 31539 26333
rect 31726 26336 32597 26364
rect 25271 26268 26096 26296
rect 25271 26265 25283 26268
rect 25225 26259 25283 26265
rect 27430 26256 27436 26308
rect 27488 26296 27494 26308
rect 27709 26299 27767 26305
rect 27709 26296 27721 26299
rect 27488 26268 27721 26296
rect 27488 26256 27494 26268
rect 27709 26265 27721 26268
rect 27755 26265 27767 26299
rect 27709 26259 27767 26265
rect 28353 26299 28411 26305
rect 28353 26265 28365 26299
rect 28399 26296 28411 26299
rect 28442 26296 28448 26308
rect 28399 26268 28448 26296
rect 28399 26265 28411 26268
rect 28353 26259 28411 26265
rect 28442 26256 28448 26268
rect 28500 26256 28506 26308
rect 31110 26256 31116 26308
rect 31168 26296 31174 26308
rect 31297 26299 31355 26305
rect 31297 26296 31309 26299
rect 31168 26268 31309 26296
rect 31168 26256 31174 26268
rect 31297 26265 31309 26268
rect 31343 26296 31355 26299
rect 31726 26296 31754 26336
rect 32585 26333 32597 26336
rect 32631 26364 32643 26367
rect 33226 26364 33232 26376
rect 32631 26336 33232 26364
rect 32631 26333 32643 26336
rect 32585 26327 32643 26333
rect 33226 26324 33232 26336
rect 33284 26364 33290 26376
rect 47857 26367 47915 26373
rect 47857 26364 47869 26367
rect 33284 26336 47869 26364
rect 33284 26324 33290 26336
rect 47857 26333 47869 26336
rect 47903 26333 47915 26367
rect 48130 26364 48136 26376
rect 48091 26336 48136 26364
rect 47857 26327 47915 26333
rect 48130 26324 48136 26336
rect 48188 26324 48194 26376
rect 31343 26268 31754 26296
rect 31343 26265 31355 26268
rect 31297 26259 31355 26265
rect 30466 26228 30472 26240
rect 30379 26200 30472 26228
rect 30466 26188 30472 26200
rect 30524 26228 30530 26240
rect 31018 26228 31024 26240
rect 30524 26200 31024 26228
rect 30524 26188 30530 26200
rect 31018 26188 31024 26200
rect 31076 26188 31082 26240
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 21818 26024 21824 26036
rect 21779 25996 21824 26024
rect 21818 25984 21824 25996
rect 21876 25984 21882 26036
rect 30190 25984 30196 26036
rect 30248 26024 30254 26036
rect 30285 26027 30343 26033
rect 30285 26024 30297 26027
rect 30248 25996 30297 26024
rect 30248 25984 30254 25996
rect 30285 25993 30297 25996
rect 30331 25993 30343 26027
rect 31018 26024 31024 26036
rect 30979 25996 31024 26024
rect 30285 25987 30343 25993
rect 31018 25984 31024 25996
rect 31076 25984 31082 26036
rect 32766 26024 32772 26036
rect 32727 25996 32772 26024
rect 32766 25984 32772 25996
rect 32824 25984 32830 26036
rect 1578 25956 1584 25968
rect 1539 25928 1584 25956
rect 1578 25916 1584 25928
rect 1636 25916 1642 25968
rect 48130 25956 48136 25968
rect 48091 25928 48136 25956
rect 48130 25916 48136 25928
rect 48188 25916 48194 25968
rect 24578 25888 24584 25900
rect 24539 25860 24584 25888
rect 24578 25848 24584 25860
rect 24636 25848 24642 25900
rect 24762 25888 24768 25900
rect 24723 25860 24768 25888
rect 24762 25848 24768 25860
rect 24820 25848 24826 25900
rect 27249 25891 27307 25897
rect 27249 25857 27261 25891
rect 27295 25888 27307 25891
rect 28166 25888 28172 25900
rect 27295 25860 28172 25888
rect 27295 25857 27307 25860
rect 27249 25851 27307 25857
rect 28166 25848 28172 25860
rect 28224 25848 28230 25900
rect 29917 25891 29975 25897
rect 29917 25857 29929 25891
rect 29963 25888 29975 25891
rect 30374 25888 30380 25900
rect 29963 25860 30380 25888
rect 29963 25857 29975 25860
rect 29917 25851 29975 25857
rect 30374 25848 30380 25860
rect 30432 25848 30438 25900
rect 31021 25891 31079 25897
rect 31021 25857 31033 25891
rect 31067 25888 31079 25891
rect 31110 25888 31116 25900
rect 31067 25860 31116 25888
rect 31067 25857 31079 25860
rect 31021 25851 31079 25857
rect 31110 25848 31116 25860
rect 31168 25848 31174 25900
rect 31205 25891 31263 25897
rect 31205 25857 31217 25891
rect 31251 25888 31263 25891
rect 31570 25888 31576 25900
rect 31251 25860 31576 25888
rect 31251 25857 31263 25860
rect 31205 25851 31263 25857
rect 31570 25848 31576 25860
rect 31628 25848 31634 25900
rect 26142 25780 26148 25832
rect 26200 25820 26206 25832
rect 27157 25823 27215 25829
rect 27157 25820 27169 25823
rect 26200 25792 27169 25820
rect 26200 25780 26206 25792
rect 27157 25789 27169 25792
rect 27203 25789 27215 25823
rect 27157 25783 27215 25789
rect 27617 25823 27675 25829
rect 27617 25789 27629 25823
rect 27663 25820 27675 25823
rect 27706 25820 27712 25832
rect 27663 25792 27712 25820
rect 27663 25789 27675 25792
rect 27617 25783 27675 25789
rect 27706 25780 27712 25792
rect 27764 25780 27770 25832
rect 29822 25820 29828 25832
rect 29783 25792 29828 25820
rect 29822 25780 29828 25792
rect 29880 25780 29886 25832
rect 20530 25684 20536 25696
rect 20491 25656 20536 25684
rect 20530 25644 20536 25656
rect 20588 25644 20594 25696
rect 22462 25684 22468 25696
rect 22423 25656 22468 25684
rect 22462 25644 22468 25656
rect 22520 25644 22526 25696
rect 24673 25687 24731 25693
rect 24673 25653 24685 25687
rect 24719 25684 24731 25687
rect 24854 25684 24860 25696
rect 24719 25656 24860 25684
rect 24719 25653 24731 25656
rect 24673 25647 24731 25653
rect 24854 25644 24860 25656
rect 24912 25644 24918 25696
rect 25501 25687 25559 25693
rect 25501 25653 25513 25687
rect 25547 25684 25559 25687
rect 26234 25684 26240 25696
rect 25547 25656 26240 25684
rect 25547 25653 25559 25656
rect 25501 25647 25559 25653
rect 26234 25644 26240 25656
rect 26292 25644 26298 25696
rect 32030 25644 32036 25696
rect 32088 25684 32094 25696
rect 32125 25687 32183 25693
rect 32125 25684 32137 25687
rect 32088 25656 32137 25684
rect 32088 25644 32094 25656
rect 32125 25653 32137 25656
rect 32171 25653 32183 25687
rect 32125 25647 32183 25653
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 25133 25483 25191 25489
rect 25133 25449 25145 25483
rect 25179 25480 25191 25483
rect 27338 25480 27344 25492
rect 25179 25452 27344 25480
rect 25179 25449 25191 25452
rect 25133 25443 25191 25449
rect 27338 25440 27344 25452
rect 27396 25440 27402 25492
rect 28166 25480 28172 25492
rect 28127 25452 28172 25480
rect 28166 25440 28172 25452
rect 28224 25440 28230 25492
rect 28258 25440 28264 25492
rect 28316 25480 28322 25492
rect 28813 25483 28871 25489
rect 28813 25480 28825 25483
rect 28316 25452 28825 25480
rect 28316 25440 28322 25452
rect 28813 25449 28825 25452
rect 28859 25480 28871 25483
rect 29270 25480 29276 25492
rect 28859 25452 29276 25480
rect 28859 25449 28871 25452
rect 28813 25443 28871 25449
rect 29270 25440 29276 25452
rect 29328 25440 29334 25492
rect 31110 25440 31116 25492
rect 31168 25480 31174 25492
rect 31297 25483 31355 25489
rect 31297 25480 31309 25483
rect 31168 25452 31309 25480
rect 31168 25440 31174 25452
rect 31297 25449 31309 25452
rect 31343 25449 31355 25483
rect 31297 25443 31355 25449
rect 31570 25440 31576 25492
rect 31628 25480 31634 25492
rect 31849 25483 31907 25489
rect 31849 25480 31861 25483
rect 31628 25452 31861 25480
rect 31628 25440 31634 25452
rect 31849 25449 31861 25452
rect 31895 25449 31907 25483
rect 31849 25443 31907 25449
rect 25774 25412 25780 25424
rect 25735 25384 25780 25412
rect 25774 25372 25780 25384
rect 25832 25372 25838 25424
rect 26142 25372 26148 25424
rect 26200 25412 26206 25424
rect 27433 25415 27491 25421
rect 27433 25412 27445 25415
rect 26200 25384 27445 25412
rect 26200 25372 26206 25384
rect 27433 25381 27445 25384
rect 27479 25381 27491 25415
rect 27433 25375 27491 25381
rect 27525 25415 27583 25421
rect 27525 25381 27537 25415
rect 27571 25412 27583 25415
rect 29822 25412 29828 25424
rect 27571 25384 29828 25412
rect 27571 25381 27583 25384
rect 27525 25375 27583 25381
rect 29822 25372 29828 25384
rect 29880 25372 29886 25424
rect 24946 25344 24952 25356
rect 24907 25316 24952 25344
rect 24946 25304 24952 25316
rect 25004 25304 25010 25356
rect 26789 25347 26847 25353
rect 26789 25313 26801 25347
rect 26835 25344 26847 25347
rect 27617 25347 27675 25353
rect 26835 25316 27384 25344
rect 26835 25313 26847 25316
rect 26789 25307 26847 25313
rect 24854 25276 24860 25288
rect 24815 25248 24860 25276
rect 24854 25236 24860 25248
rect 24912 25236 24918 25288
rect 26694 25276 26700 25288
rect 26655 25248 26700 25276
rect 26694 25236 26700 25248
rect 26752 25236 26758 25288
rect 27356 25285 27384 25316
rect 27617 25313 27629 25347
rect 27663 25313 27675 25347
rect 27617 25307 27675 25313
rect 26881 25279 26939 25285
rect 26881 25245 26893 25279
rect 26927 25245 26939 25279
rect 26881 25239 26939 25245
rect 27341 25279 27399 25285
rect 27341 25245 27353 25279
rect 27387 25245 27399 25279
rect 27632 25276 27660 25307
rect 28074 25276 28080 25288
rect 27632 25248 28080 25276
rect 27341 25239 27399 25245
rect 26896 25208 26924 25239
rect 28074 25236 28080 25248
rect 28132 25236 28138 25288
rect 28258 25276 28264 25288
rect 28219 25248 28264 25276
rect 28258 25236 28264 25248
rect 28316 25236 28322 25288
rect 27982 25208 27988 25220
rect 26896 25180 27988 25208
rect 27982 25168 27988 25180
rect 28040 25168 28046 25220
rect 23477 25143 23535 25149
rect 23477 25109 23489 25143
rect 23523 25140 23535 25143
rect 23750 25140 23756 25152
rect 23523 25112 23756 25140
rect 23523 25109 23535 25112
rect 23477 25103 23535 25109
rect 23750 25100 23756 25112
rect 23808 25100 23814 25152
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 24857 24939 24915 24945
rect 24857 24905 24869 24939
rect 24903 24936 24915 24939
rect 26142 24936 26148 24948
rect 24903 24908 26148 24936
rect 24903 24905 24915 24908
rect 24857 24899 24915 24905
rect 26142 24896 26148 24908
rect 26200 24896 26206 24948
rect 28074 24936 28080 24948
rect 28035 24908 28080 24936
rect 28074 24896 28080 24908
rect 28132 24896 28138 24948
rect 27172 24840 28120 24868
rect 27172 24812 27200 24840
rect 23750 24800 23756 24812
rect 23711 24772 23756 24800
rect 23750 24760 23756 24772
rect 23808 24760 23814 24812
rect 23934 24800 23940 24812
rect 23895 24772 23940 24800
rect 23934 24760 23940 24772
rect 23992 24760 23998 24812
rect 24578 24800 24584 24812
rect 24539 24772 24584 24800
rect 24578 24760 24584 24772
rect 24636 24760 24642 24812
rect 24949 24803 25007 24809
rect 24949 24769 24961 24803
rect 24995 24769 25007 24803
rect 24949 24763 25007 24769
rect 23198 24692 23204 24744
rect 23256 24732 23262 24744
rect 23293 24735 23351 24741
rect 23293 24732 23305 24735
rect 23256 24704 23305 24732
rect 23256 24692 23262 24704
rect 23293 24701 23305 24704
rect 23339 24732 23351 24735
rect 23952 24732 23980 24760
rect 23339 24704 23980 24732
rect 24121 24735 24179 24741
rect 23339 24701 23351 24704
rect 23293 24695 23351 24701
rect 24121 24701 24133 24735
rect 24167 24732 24179 24735
rect 24762 24732 24768 24744
rect 24167 24704 24768 24732
rect 24167 24701 24179 24704
rect 24121 24695 24179 24701
rect 24762 24692 24768 24704
rect 24820 24732 24826 24744
rect 24964 24732 24992 24763
rect 25038 24760 25044 24812
rect 25096 24800 25102 24812
rect 26421 24803 26479 24809
rect 25096 24772 25141 24800
rect 25096 24760 25102 24772
rect 26421 24769 26433 24803
rect 26467 24800 26479 24803
rect 26694 24800 26700 24812
rect 26467 24772 26700 24800
rect 26467 24769 26479 24772
rect 26421 24763 26479 24769
rect 26694 24760 26700 24772
rect 26752 24800 26758 24812
rect 27154 24800 27160 24812
rect 26752 24772 27160 24800
rect 26752 24760 26758 24772
rect 27154 24760 27160 24772
rect 27212 24760 27218 24812
rect 27341 24803 27399 24809
rect 27341 24769 27353 24803
rect 27387 24800 27399 24803
rect 27982 24800 27988 24812
rect 27387 24772 27988 24800
rect 27387 24769 27399 24772
rect 27341 24763 27399 24769
rect 27982 24760 27988 24772
rect 28040 24760 28046 24812
rect 28092 24800 28120 24840
rect 28169 24803 28227 24809
rect 28169 24800 28181 24803
rect 28092 24772 28181 24800
rect 28169 24769 28181 24772
rect 28215 24800 28227 24803
rect 28629 24803 28687 24809
rect 28629 24800 28641 24803
rect 28215 24772 28641 24800
rect 28215 24769 28227 24772
rect 28169 24763 28227 24769
rect 28629 24769 28641 24772
rect 28675 24769 28687 24803
rect 28629 24763 28687 24769
rect 24820 24704 24992 24732
rect 27525 24735 27583 24741
rect 24820 24692 24826 24704
rect 27525 24701 27537 24735
rect 27571 24732 27583 24735
rect 28258 24732 28264 24744
rect 27571 24704 28264 24732
rect 27571 24701 27583 24704
rect 27525 24695 27583 24701
rect 28258 24692 28264 24704
rect 28316 24692 28322 24744
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 2225 24395 2283 24401
rect 2225 24361 2237 24395
rect 2271 24392 2283 24395
rect 8938 24392 8944 24404
rect 2271 24364 8944 24392
rect 2271 24361 2283 24364
rect 2225 24355 2283 24361
rect 1673 24191 1731 24197
rect 1673 24157 1685 24191
rect 1719 24188 1731 24191
rect 2240 24188 2268 24355
rect 8938 24352 8944 24364
rect 8996 24352 9002 24404
rect 24489 24395 24547 24401
rect 24489 24361 24501 24395
rect 24535 24392 24547 24395
rect 24578 24392 24584 24404
rect 24535 24364 24584 24392
rect 24535 24361 24547 24364
rect 24489 24355 24547 24361
rect 24578 24352 24584 24364
rect 24636 24352 24642 24404
rect 25133 24395 25191 24401
rect 25133 24361 25145 24395
rect 25179 24392 25191 24395
rect 26602 24392 26608 24404
rect 25179 24364 26608 24392
rect 25179 24361 25191 24364
rect 25133 24355 25191 24361
rect 23934 24216 23940 24268
rect 23992 24256 23998 24268
rect 23992 24228 24624 24256
rect 23992 24216 23998 24228
rect 1719 24160 2268 24188
rect 1719 24157 1731 24160
rect 1673 24151 1731 24157
rect 23750 24148 23756 24200
rect 23808 24188 23814 24200
rect 24596 24197 24624 24228
rect 24397 24191 24455 24197
rect 24397 24188 24409 24191
rect 23808 24160 24409 24188
rect 23808 24148 23814 24160
rect 24397 24157 24409 24160
rect 24443 24157 24455 24191
rect 24397 24151 24455 24157
rect 24581 24191 24639 24197
rect 24581 24157 24593 24191
rect 24627 24188 24639 24191
rect 25148 24188 25176 24355
rect 26602 24352 26608 24364
rect 26660 24352 26666 24404
rect 27709 24395 27767 24401
rect 27709 24361 27721 24395
rect 27755 24392 27767 24395
rect 27982 24392 27988 24404
rect 27755 24364 27988 24392
rect 27755 24361 27767 24364
rect 27709 24355 27767 24361
rect 27982 24352 27988 24364
rect 28040 24392 28046 24404
rect 28261 24395 28319 24401
rect 28261 24392 28273 24395
rect 28040 24364 28273 24392
rect 28040 24352 28046 24364
rect 28261 24361 28273 24364
rect 28307 24361 28319 24395
rect 28261 24355 28319 24361
rect 39758 24352 39764 24404
rect 39816 24392 39822 24404
rect 47765 24395 47823 24401
rect 47765 24392 47777 24395
rect 39816 24364 47777 24392
rect 39816 24352 39822 24364
rect 47765 24361 47777 24364
rect 47811 24361 47823 24395
rect 47765 24355 47823 24361
rect 24627 24160 25176 24188
rect 24627 24157 24639 24160
rect 24581 24151 24639 24157
rect 48041 24123 48099 24129
rect 48041 24089 48053 24123
rect 48087 24120 48099 24123
rect 48130 24120 48136 24132
rect 48087 24092 48136 24120
rect 48087 24089 48099 24092
rect 48041 24083 48099 24089
rect 48130 24080 48136 24092
rect 48188 24080 48194 24132
rect 1486 24052 1492 24064
rect 1447 24024 1492 24052
rect 1486 24012 1492 24024
rect 1544 24012 1550 24064
rect 23750 24052 23756 24064
rect 23711 24024 23756 24052
rect 23750 24012 23756 24024
rect 23808 24012 23814 24064
rect 27065 24055 27123 24061
rect 27065 24021 27077 24055
rect 27111 24052 27123 24055
rect 27154 24052 27160 24064
rect 27111 24024 27160 24052
rect 27111 24021 27123 24024
rect 27065 24015 27123 24021
rect 27154 24012 27160 24024
rect 27212 24012 27218 24064
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 48130 23848 48136 23860
rect 48091 23820 48136 23848
rect 48130 23808 48136 23820
rect 48188 23808 48194 23860
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 36998 21972 37004 22024
rect 37056 22012 37062 22024
rect 47305 22015 47363 22021
rect 47305 22012 47317 22015
rect 37056 21984 47317 22012
rect 37056 21972 37062 21984
rect 47305 21981 47317 21984
rect 47351 22012 47363 22015
rect 47857 22015 47915 22021
rect 47857 22012 47869 22015
rect 47351 21984 47869 22012
rect 47351 21981 47363 21984
rect 47305 21975 47363 21981
rect 47857 21981 47869 21984
rect 47903 21981 47915 22015
rect 47857 21975 47915 21981
rect 1578 21904 1584 21956
rect 1636 21944 1642 21956
rect 1857 21947 1915 21953
rect 1857 21944 1869 21947
rect 1636 21916 1869 21944
rect 1636 21904 1642 21916
rect 1857 21913 1869 21916
rect 1903 21913 1915 21947
rect 1857 21907 1915 21913
rect 1949 21879 2007 21885
rect 1949 21845 1961 21879
rect 1995 21876 2007 21879
rect 15746 21876 15752 21888
rect 1995 21848 15752 21876
rect 1995 21845 2007 21848
rect 1949 21839 2007 21845
rect 15746 21836 15752 21848
rect 15804 21836 15810 21888
rect 48038 21876 48044 21888
rect 47999 21848 48044 21876
rect 48038 21836 48044 21848
rect 48096 21836 48102 21888
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 1578 21672 1584 21684
rect 1539 21644 1584 21672
rect 1578 21632 1584 21644
rect 1636 21632 1642 21684
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 39390 20000 39396 20052
rect 39448 20040 39454 20052
rect 47305 20043 47363 20049
rect 47305 20040 47317 20043
rect 39448 20012 47317 20040
rect 39448 20000 39454 20012
rect 47305 20009 47317 20012
rect 47351 20009 47363 20043
rect 47305 20003 47363 20009
rect 47320 19836 47348 20003
rect 47857 19839 47915 19845
rect 47857 19836 47869 19839
rect 47320 19808 47869 19836
rect 47857 19805 47869 19808
rect 47903 19805 47915 19839
rect 47857 19799 47915 19805
rect 1854 19768 1860 19780
rect 1815 19740 1860 19768
rect 1854 19728 1860 19740
rect 1912 19728 1918 19780
rect 2133 19703 2191 19709
rect 2133 19669 2145 19703
rect 2179 19700 2191 19703
rect 13998 19700 14004 19712
rect 2179 19672 14004 19700
rect 2179 19669 2191 19672
rect 2133 19663 2191 19669
rect 13998 19660 14004 19672
rect 14056 19660 14062 19712
rect 48038 19700 48044 19712
rect 47999 19672 48044 19700
rect 48038 19660 48044 19672
rect 48096 19660 48102 19712
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 1673 19499 1731 19505
rect 1673 19465 1685 19499
rect 1719 19496 1731 19499
rect 1854 19496 1860 19508
rect 1719 19468 1860 19496
rect 1719 19465 1731 19468
rect 1673 19459 1731 19465
rect 1854 19456 1860 19468
rect 1912 19456 1918 19508
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 1578 18232 1584 18284
rect 1636 18272 1642 18284
rect 1857 18275 1915 18281
rect 1857 18272 1869 18275
rect 1636 18244 1869 18272
rect 1636 18232 1642 18244
rect 1857 18241 1869 18244
rect 1903 18241 1915 18275
rect 1857 18235 1915 18241
rect 41230 18232 41236 18284
rect 41288 18272 41294 18284
rect 47670 18272 47676 18284
rect 41288 18244 47676 18272
rect 41288 18232 41294 18244
rect 47670 18232 47676 18244
rect 47728 18272 47734 18284
rect 47857 18275 47915 18281
rect 47857 18272 47869 18275
rect 47728 18244 47869 18272
rect 47728 18232 47734 18244
rect 47857 18241 47869 18244
rect 47903 18241 47915 18275
rect 47857 18235 47915 18241
rect 1949 18071 2007 18077
rect 1949 18037 1961 18071
rect 1995 18068 2007 18071
rect 9858 18068 9864 18080
rect 1995 18040 9864 18068
rect 1995 18037 2007 18040
rect 1949 18031 2007 18037
rect 9858 18028 9864 18040
rect 9916 18028 9922 18080
rect 48038 18068 48044 18080
rect 47999 18040 48044 18068
rect 48038 18028 48044 18040
rect 48096 18028 48102 18080
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 47670 17864 47676 17876
rect 47631 17836 47676 17864
rect 47670 17824 47676 17836
rect 47728 17824 47734 17876
rect 1578 17796 1584 17808
rect 1539 17768 1584 17796
rect 1578 17756 1584 17768
rect 1636 17756 1642 17808
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 42058 16192 42064 16244
rect 42116 16232 42122 16244
rect 47949 16235 48007 16241
rect 47949 16232 47961 16235
rect 42116 16204 47961 16232
rect 42116 16192 42122 16204
rect 47949 16201 47961 16204
rect 47995 16201 48007 16235
rect 47949 16195 48007 16201
rect 1578 16056 1584 16108
rect 1636 16096 1642 16108
rect 1857 16099 1915 16105
rect 1857 16096 1869 16099
rect 1636 16068 1869 16096
rect 1636 16056 1642 16068
rect 1857 16065 1869 16068
rect 1903 16065 1915 16099
rect 48130 16096 48136 16108
rect 48091 16068 48136 16096
rect 1857 16059 1915 16065
rect 48130 16056 48136 16068
rect 48188 16056 48194 16108
rect 2133 15895 2191 15901
rect 2133 15861 2145 15895
rect 2179 15892 2191 15895
rect 39574 15892 39580 15904
rect 2179 15864 39580 15892
rect 2179 15861 2191 15864
rect 2133 15855 2191 15861
rect 39574 15852 39580 15864
rect 39632 15852 39638 15904
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 1578 15688 1584 15700
rect 1539 15660 1584 15688
rect 1578 15648 1584 15660
rect 1636 15648 1642 15700
rect 48130 15688 48136 15700
rect 48091 15660 48136 15688
rect 48130 15648 48136 15660
rect 48188 15648 48194 15700
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 1394 13920 1400 13932
rect 1355 13892 1400 13920
rect 1394 13880 1400 13892
rect 1452 13880 1458 13932
rect 47854 13920 47860 13932
rect 47815 13892 47860 13920
rect 47854 13880 47860 13892
rect 47912 13880 47918 13932
rect 35618 13852 35624 13864
rect 1596 13824 35624 13852
rect 1596 13793 1624 13824
rect 35618 13812 35624 13824
rect 35676 13812 35682 13864
rect 1581 13787 1639 13793
rect 1581 13753 1593 13787
rect 1627 13753 1639 13787
rect 1581 13747 1639 13753
rect 48038 13716 48044 13728
rect 47999 13688 48044 13716
rect 48038 13676 48044 13688
rect 48096 13676 48102 13728
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 1394 13512 1400 13524
rect 1355 13484 1400 13512
rect 1394 13472 1400 13484
rect 1452 13472 1458 13524
rect 47765 13515 47823 13521
rect 47765 13481 47777 13515
rect 47811 13512 47823 13515
rect 47854 13512 47860 13524
rect 47811 13484 47860 13512
rect 47811 13481 47823 13484
rect 47765 13475 47823 13481
rect 47854 13472 47860 13484
rect 47912 13472 47918 13524
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 47762 11840 47768 11892
rect 47820 11880 47826 11892
rect 47949 11883 48007 11889
rect 47949 11880 47961 11883
rect 47820 11852 47961 11880
rect 47820 11840 47826 11852
rect 47949 11849 47961 11852
rect 47995 11849 48007 11883
rect 47949 11843 48007 11849
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11744 1731 11747
rect 48130 11744 48136 11756
rect 1719 11716 2268 11744
rect 48091 11716 48136 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 1486 11608 1492 11620
rect 1447 11580 1492 11608
rect 1486 11568 1492 11580
rect 1544 11568 1550 11620
rect 2240 11617 2268 11716
rect 48130 11704 48136 11716
rect 48188 11704 48194 11756
rect 2225 11611 2283 11617
rect 2225 11577 2237 11611
rect 2271 11608 2283 11611
rect 27430 11608 27436 11620
rect 2271 11580 27436 11608
rect 2271 11577 2283 11580
rect 2225 11571 2283 11577
rect 27430 11568 27436 11580
rect 27488 11568 27494 11620
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 48130 11336 48136 11348
rect 48091 11308 48136 11336
rect 48130 11296 48136 11308
rect 48188 11296 48194 11348
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 31662 10004 31668 10056
rect 31720 10044 31726 10056
rect 47305 10047 47363 10053
rect 47305 10044 47317 10047
rect 31720 10016 47317 10044
rect 31720 10004 31726 10016
rect 47305 10013 47317 10016
rect 47351 10044 47363 10047
rect 47857 10047 47915 10053
rect 47857 10044 47869 10047
rect 47351 10016 47869 10044
rect 47351 10013 47363 10016
rect 47305 10007 47363 10013
rect 47857 10013 47869 10016
rect 47903 10013 47915 10047
rect 47857 10007 47915 10013
rect 1578 9936 1584 9988
rect 1636 9976 1642 9988
rect 1857 9979 1915 9985
rect 1857 9976 1869 9979
rect 1636 9948 1869 9976
rect 1636 9936 1642 9948
rect 1857 9945 1869 9948
rect 1903 9945 1915 9979
rect 1857 9939 1915 9945
rect 2133 9911 2191 9917
rect 2133 9877 2145 9911
rect 2179 9908 2191 9911
rect 31110 9908 31116 9920
rect 2179 9880 31116 9908
rect 2179 9877 2191 9880
rect 2133 9871 2191 9877
rect 31110 9868 31116 9880
rect 31168 9868 31174 9920
rect 48038 9908 48044 9920
rect 47999 9880 48044 9908
rect 48038 9868 48044 9880
rect 48096 9868 48102 9920
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 1578 9636 1584 9648
rect 1539 9608 1584 9636
rect 1578 9596 1584 9608
rect 1636 9596 1642 9648
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 47946 8072 47952 8084
rect 47907 8044 47952 8072
rect 47946 8032 47952 8044
rect 48004 8032 48010 8084
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7868 1731 7871
rect 2225 7871 2283 7877
rect 2225 7868 2237 7871
rect 1719 7840 2237 7868
rect 1719 7837 1731 7840
rect 1673 7831 1731 7837
rect 2225 7837 2237 7840
rect 2271 7868 2283 7871
rect 14918 7868 14924 7880
rect 2271 7840 14924 7868
rect 2271 7837 2283 7840
rect 2225 7831 2283 7837
rect 14918 7828 14924 7840
rect 14976 7828 14982 7880
rect 47397 7803 47455 7809
rect 47397 7769 47409 7803
rect 47443 7800 47455 7803
rect 48038 7800 48044 7812
rect 47443 7772 48044 7800
rect 47443 7769 47455 7772
rect 47397 7763 47455 7769
rect 48038 7760 48044 7772
rect 48096 7760 48102 7812
rect 1486 7732 1492 7744
rect 1447 7704 1492 7732
rect 1486 7692 1492 7704
rect 1544 7692 1550 7744
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 1578 5584 1584 5636
rect 1636 5624 1642 5636
rect 1857 5627 1915 5633
rect 1857 5624 1869 5627
rect 1636 5596 1869 5624
rect 1636 5584 1642 5596
rect 1857 5593 1869 5596
rect 1903 5593 1915 5627
rect 47857 5627 47915 5633
rect 47857 5624 47869 5627
rect 1857 5587 1915 5593
rect 26206 5596 47869 5624
rect 1949 5559 2007 5565
rect 1949 5525 1961 5559
rect 1995 5556 2007 5559
rect 11514 5556 11520 5568
rect 1995 5528 11520 5556
rect 1995 5525 2007 5528
rect 1949 5519 2007 5525
rect 11514 5516 11520 5528
rect 11572 5516 11578 5568
rect 22462 5516 22468 5568
rect 22520 5556 22526 5568
rect 26206 5556 26234 5596
rect 47857 5593 47869 5596
rect 47903 5593 47915 5627
rect 48038 5624 48044 5636
rect 47999 5596 48044 5624
rect 47857 5587 47915 5593
rect 48038 5584 48044 5596
rect 48096 5584 48102 5636
rect 22520 5528 26234 5556
rect 47397 5559 47455 5565
rect 22520 5516 22526 5528
rect 47397 5525 47409 5559
rect 47443 5556 47455 5559
rect 48056 5556 48084 5584
rect 47443 5528 48084 5556
rect 47443 5525 47455 5528
rect 47397 5519 47455 5525
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 1578 5352 1584 5364
rect 1539 5324 1584 5352
rect 1578 5312 1584 5324
rect 1636 5312 1642 5364
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 39482 4088 39488 4140
rect 39540 4128 39546 4140
rect 47581 4131 47639 4137
rect 47581 4128 47593 4131
rect 39540 4100 47593 4128
rect 39540 4088 39546 4100
rect 47581 4097 47593 4100
rect 47627 4128 47639 4131
rect 47762 4128 47768 4140
rect 47627 4100 47768 4128
rect 47627 4097 47639 4100
rect 47581 4091 47639 4097
rect 47762 4088 47768 4100
rect 47820 4088 47826 4140
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 47302 3584 47308 3596
rect 47263 3556 47308 3584
rect 47302 3544 47308 3556
rect 47360 3544 47366 3596
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3485 1731 3519
rect 47320 3516 47348 3544
rect 47857 3519 47915 3525
rect 47857 3516 47869 3519
rect 47320 3488 47869 3516
rect 1673 3479 1731 3485
rect 47857 3485 47869 3488
rect 47903 3485 47915 3519
rect 47857 3479 47915 3485
rect 1688 3448 1716 3479
rect 2225 3451 2283 3457
rect 2225 3448 2237 3451
rect 1688 3420 2237 3448
rect 2225 3417 2237 3420
rect 2271 3448 2283 3451
rect 15470 3448 15476 3460
rect 2271 3420 15476 3448
rect 2271 3417 2283 3420
rect 2225 3411 2283 3417
rect 15470 3408 15476 3420
rect 15528 3408 15534 3460
rect 46845 3451 46903 3457
rect 46845 3417 46857 3451
rect 46891 3448 46903 3451
rect 48314 3448 48320 3460
rect 46891 3420 48320 3448
rect 46891 3417 46903 3420
rect 46845 3411 46903 3417
rect 48314 3408 48320 3420
rect 48372 3408 48378 3460
rect 1486 3380 1492 3392
rect 1447 3352 1492 3380
rect 1486 3340 1492 3352
rect 1544 3340 1550 3392
rect 48038 3380 48044 3392
rect 47999 3352 48044 3380
rect 48038 3340 48044 3352
rect 48096 3340 48102 3392
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 32217 3179 32275 3185
rect 32217 3145 32229 3179
rect 32263 3176 32275 3179
rect 32582 3176 32588 3188
rect 32263 3148 32588 3176
rect 32263 3145 32275 3148
rect 32217 3139 32275 3145
rect 32582 3136 32588 3148
rect 32640 3136 32646 3188
rect 1394 3040 1400 3052
rect 1355 3012 1400 3040
rect 1394 3000 1400 3012
rect 1452 3040 1458 3052
rect 2685 3043 2743 3049
rect 2685 3040 2697 3043
rect 1452 3012 2697 3040
rect 1452 3000 1458 3012
rect 2685 3009 2697 3012
rect 2731 3009 2743 3043
rect 2685 3003 2743 3009
rect 48133 3043 48191 3049
rect 48133 3009 48145 3043
rect 48179 3040 48191 3043
rect 48314 3040 48320 3052
rect 48179 3012 48320 3040
rect 48179 3009 48191 3012
rect 48133 3003 48191 3009
rect 48314 3000 48320 3012
rect 48372 3040 48378 3052
rect 49602 3040 49608 3052
rect 48372 3012 49608 3040
rect 48372 3000 48378 3012
rect 49602 3000 49608 3012
rect 49660 3000 49666 3052
rect 4249 2975 4307 2981
rect 4249 2941 4261 2975
rect 4295 2972 4307 2975
rect 4614 2972 4620 2984
rect 4295 2944 4620 2972
rect 4295 2941 4307 2944
rect 4249 2935 4307 2941
rect 4614 2932 4620 2944
rect 4672 2972 4678 2984
rect 28810 2972 28816 2984
rect 4672 2944 28816 2972
rect 4672 2932 4678 2944
rect 28810 2932 28816 2944
rect 28868 2932 28874 2984
rect 46566 2972 46572 2984
rect 46527 2944 46572 2972
rect 46566 2932 46572 2944
rect 46624 2932 46630 2984
rect 1581 2907 1639 2913
rect 1581 2873 1593 2907
rect 1627 2904 1639 2907
rect 10962 2904 10968 2916
rect 1627 2876 10968 2904
rect 1627 2873 1639 2876
rect 1581 2867 1639 2873
rect 10962 2864 10968 2876
rect 11020 2864 11026 2916
rect 11974 2904 11980 2916
rect 11935 2876 11980 2904
rect 11974 2864 11980 2876
rect 12032 2864 12038 2916
rect 36078 2864 36084 2916
rect 36136 2904 36142 2916
rect 47949 2907 48007 2913
rect 47949 2904 47961 2907
rect 36136 2876 47961 2904
rect 36136 2864 36142 2876
rect 47949 2873 47961 2876
rect 47995 2873 48007 2907
rect 47949 2867 48007 2873
rect 14 2796 20 2848
rect 72 2836 78 2848
rect 2130 2836 2136 2848
rect 72 2808 2136 2836
rect 72 2796 78 2808
rect 2130 2796 2136 2808
rect 2188 2796 2194 2848
rect 9030 2796 9036 2848
rect 9088 2836 9094 2848
rect 9125 2839 9183 2845
rect 9125 2836 9137 2839
rect 9088 2808 9137 2836
rect 9088 2796 9094 2808
rect 9125 2805 9137 2808
rect 9171 2805 9183 2839
rect 9125 2799 9183 2805
rect 16758 2796 16764 2848
rect 16816 2836 16822 2848
rect 16853 2839 16911 2845
rect 16853 2836 16865 2839
rect 16816 2808 16865 2836
rect 16816 2796 16822 2808
rect 16853 2805 16865 2808
rect 16899 2805 16911 2839
rect 16853 2799 16911 2805
rect 18690 2796 18696 2848
rect 18748 2836 18754 2848
rect 19429 2839 19487 2845
rect 19429 2836 19441 2839
rect 18748 2808 19441 2836
rect 18748 2796 18754 2808
rect 19429 2805 19441 2808
rect 19475 2836 19487 2839
rect 19702 2836 19708 2848
rect 19475 2808 19708 2836
rect 19475 2805 19487 2808
rect 19429 2799 19487 2805
rect 19702 2796 19708 2808
rect 19760 2796 19766 2848
rect 20625 2839 20683 2845
rect 20625 2805 20637 2839
rect 20671 2836 20683 2839
rect 20714 2836 20720 2848
rect 20671 2808 20720 2836
rect 20671 2805 20683 2808
rect 20625 2799 20683 2805
rect 20714 2796 20720 2808
rect 20772 2796 20778 2848
rect 24486 2796 24492 2848
rect 24544 2836 24550 2848
rect 24581 2839 24639 2845
rect 24581 2836 24593 2839
rect 24544 2808 24593 2836
rect 24544 2796 24550 2808
rect 24581 2805 24593 2808
rect 24627 2805 24639 2839
rect 28350 2836 28356 2848
rect 28311 2808 28356 2836
rect 24581 2799 24639 2805
rect 28350 2796 28356 2808
rect 28408 2796 28414 2848
rect 39945 2839 40003 2845
rect 39945 2805 39957 2839
rect 39991 2836 40003 2839
rect 40034 2836 40040 2848
rect 39991 2808 40040 2836
rect 39991 2805 40003 2808
rect 39945 2799 40003 2805
rect 40034 2796 40040 2808
rect 40092 2796 40098 2848
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 9766 2632 9772 2644
rect 6886 2604 9772 2632
rect 5445 2567 5503 2573
rect 5445 2533 5457 2567
rect 5491 2564 5503 2567
rect 6886 2564 6914 2604
rect 9766 2592 9772 2604
rect 9824 2592 9830 2644
rect 20898 2632 20904 2644
rect 20859 2604 20904 2632
rect 20898 2592 20904 2604
rect 20956 2592 20962 2644
rect 23198 2632 23204 2644
rect 21468 2604 23204 2632
rect 5491 2536 6914 2564
rect 7469 2567 7527 2573
rect 5491 2533 5503 2536
rect 5445 2527 5503 2533
rect 7469 2533 7481 2567
rect 7515 2564 7527 2567
rect 9490 2564 9496 2576
rect 7515 2536 9496 2564
rect 7515 2533 7527 2536
rect 7469 2527 7527 2533
rect 9490 2524 9496 2536
rect 9548 2524 9554 2576
rect 13265 2567 13323 2573
rect 13265 2533 13277 2567
rect 13311 2564 13323 2567
rect 14550 2564 14556 2576
rect 13311 2536 14556 2564
rect 13311 2533 13323 2536
rect 13265 2527 13323 2533
rect 14550 2524 14556 2536
rect 14608 2524 14614 2576
rect 19889 2567 19947 2573
rect 19889 2533 19901 2567
rect 19935 2564 19947 2567
rect 21468 2564 21496 2604
rect 23198 2592 23204 2604
rect 23256 2592 23262 2644
rect 26234 2592 26240 2644
rect 26292 2632 26298 2644
rect 28537 2635 28595 2641
rect 28537 2632 28549 2635
rect 26292 2604 28549 2632
rect 26292 2592 26298 2604
rect 28537 2601 28549 2604
rect 28583 2601 28595 2635
rect 36354 2632 36360 2644
rect 28537 2595 28595 2601
rect 31726 2604 35848 2632
rect 36315 2604 36360 2632
rect 19935 2536 21496 2564
rect 19935 2533 19947 2536
rect 19889 2527 19947 2533
rect 22554 2524 22560 2576
rect 22612 2564 22618 2576
rect 22612 2536 23060 2564
rect 22612 2524 22618 2536
rect 1673 2499 1731 2505
rect 1673 2465 1685 2499
rect 1719 2496 1731 2499
rect 9585 2499 9643 2505
rect 1719 2468 9536 2496
rect 1719 2465 1731 2468
rect 1673 2459 1731 2465
rect 2130 2428 2136 2440
rect 2091 2400 2136 2428
rect 2130 2388 2136 2400
rect 2188 2388 2194 2440
rect 4065 2431 4123 2437
rect 4065 2397 4077 2431
rect 4111 2428 4123 2431
rect 4614 2428 4620 2440
rect 4111 2400 4620 2428
rect 4111 2397 4123 2400
rect 4065 2391 4123 2397
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 4801 2431 4859 2437
rect 4801 2397 4813 2431
rect 4847 2428 4859 2431
rect 5166 2428 5172 2440
rect 4847 2400 5172 2428
rect 4847 2397 4859 2400
rect 4801 2391 4859 2397
rect 5166 2388 5172 2400
rect 5224 2428 5230 2440
rect 5261 2431 5319 2437
rect 5261 2428 5273 2431
rect 5224 2400 5273 2428
rect 5224 2388 5230 2400
rect 5261 2397 5273 2400
rect 5307 2397 5319 2431
rect 5261 2391 5319 2397
rect 1302 2320 1308 2372
rect 1360 2360 1366 2372
rect 1489 2363 1547 2369
rect 1489 2360 1501 2363
rect 1360 2332 1501 2360
rect 1360 2320 1366 2332
rect 1489 2329 1501 2332
rect 1535 2360 1547 2363
rect 2869 2363 2927 2369
rect 2869 2360 2881 2363
rect 1535 2332 2881 2360
rect 1535 2329 1547 2332
rect 1489 2323 1547 2329
rect 2869 2329 2881 2332
rect 2915 2329 2927 2363
rect 2869 2323 2927 2329
rect 6733 2363 6791 2369
rect 6733 2329 6745 2363
rect 6779 2360 6791 2363
rect 7098 2360 7104 2372
rect 6779 2332 7104 2360
rect 6779 2329 6791 2332
rect 6733 2323 6791 2329
rect 7098 2320 7104 2332
rect 7156 2360 7162 2372
rect 7285 2363 7343 2369
rect 7285 2360 7297 2363
rect 7156 2332 7297 2360
rect 7156 2320 7162 2332
rect 7285 2329 7297 2332
rect 7331 2329 7343 2363
rect 7285 2323 7343 2329
rect 9030 2320 9036 2372
rect 9088 2360 9094 2372
rect 9401 2363 9459 2369
rect 9401 2360 9413 2363
rect 9088 2332 9413 2360
rect 9088 2320 9094 2332
rect 9401 2329 9413 2332
rect 9447 2329 9459 2363
rect 9508 2360 9536 2468
rect 9585 2465 9597 2499
rect 9631 2496 9643 2499
rect 9631 2468 20208 2496
rect 9631 2465 9643 2468
rect 9585 2459 9643 2465
rect 11793 2431 11851 2437
rect 11793 2397 11805 2431
rect 11839 2428 11851 2431
rect 11974 2428 11980 2440
rect 11839 2400 11980 2428
rect 11839 2397 11851 2400
rect 11793 2391 11851 2397
rect 11974 2388 11980 2400
rect 12032 2388 12038 2440
rect 14826 2428 14832 2440
rect 12084 2400 14832 2428
rect 12084 2360 12112 2400
rect 14826 2388 14832 2400
rect 14884 2388 14890 2440
rect 15194 2428 15200 2440
rect 15155 2400 15200 2428
rect 15194 2388 15200 2400
rect 15252 2428 15258 2440
rect 15657 2431 15715 2437
rect 15657 2428 15669 2431
rect 15252 2400 15669 2428
rect 15252 2388 15258 2400
rect 15657 2397 15669 2400
rect 15703 2397 15715 2431
rect 19702 2428 19708 2440
rect 19663 2400 19708 2428
rect 15657 2391 15715 2397
rect 19702 2388 19708 2400
rect 19760 2388 19766 2440
rect 9508 2332 12112 2360
rect 12529 2363 12587 2369
rect 9401 2323 9459 2329
rect 12529 2329 12541 2363
rect 12575 2360 12587 2363
rect 12894 2360 12900 2372
rect 12575 2332 12900 2360
rect 12575 2329 12587 2332
rect 12529 2323 12587 2329
rect 12894 2320 12900 2332
rect 12952 2360 12958 2372
rect 13081 2363 13139 2369
rect 13081 2360 13093 2363
rect 12952 2332 13093 2360
rect 12952 2320 12958 2332
rect 13081 2329 13093 2332
rect 13127 2329 13139 2363
rect 13081 2323 13139 2329
rect 16758 2320 16764 2372
rect 16816 2360 16822 2372
rect 17129 2363 17187 2369
rect 17129 2360 17141 2363
rect 16816 2332 17141 2360
rect 16816 2320 16822 2332
rect 17129 2329 17141 2332
rect 17175 2329 17187 2363
rect 20180 2360 20208 2468
rect 20530 2456 20536 2508
rect 20588 2496 20594 2508
rect 22925 2499 22983 2505
rect 22925 2496 22937 2499
rect 20588 2468 22937 2496
rect 20588 2456 20594 2468
rect 22925 2465 22937 2468
rect 22971 2465 22983 2499
rect 23032 2496 23060 2536
rect 25498 2524 25504 2576
rect 25556 2564 25562 2576
rect 31726 2564 31754 2604
rect 25556 2536 31754 2564
rect 34885 2567 34943 2573
rect 25556 2524 25562 2536
rect 34885 2533 34897 2567
rect 34931 2533 34943 2567
rect 35820 2564 35848 2604
rect 36354 2592 36360 2604
rect 36412 2592 36418 2644
rect 45278 2632 45284 2644
rect 45239 2604 45284 2632
rect 45278 2592 45284 2604
rect 45336 2592 45342 2644
rect 37553 2567 37611 2573
rect 37553 2564 37565 2567
rect 35820 2536 37565 2564
rect 34885 2527 34943 2533
rect 37553 2533 37565 2536
rect 37599 2533 37611 2567
rect 44174 2564 44180 2576
rect 44135 2536 44180 2564
rect 37553 2527 37611 2533
rect 27249 2499 27307 2505
rect 23032 2468 27200 2496
rect 22925 2459 22983 2465
rect 20714 2428 20720 2440
rect 20675 2400 20720 2428
rect 20714 2388 20720 2400
rect 20772 2388 20778 2440
rect 22189 2431 22247 2437
rect 22189 2397 22201 2431
rect 22235 2428 22247 2431
rect 22554 2428 22560 2440
rect 22235 2400 22560 2428
rect 22235 2397 22247 2400
rect 22189 2391 22247 2397
rect 22554 2388 22560 2400
rect 22612 2428 22618 2440
rect 22649 2431 22707 2437
rect 22649 2428 22661 2431
rect 22612 2400 22661 2428
rect 22612 2388 22618 2400
rect 22649 2397 22661 2400
rect 22695 2397 22707 2431
rect 26973 2431 27031 2437
rect 26973 2428 26985 2431
rect 22649 2391 22707 2397
rect 26436 2400 26985 2428
rect 23750 2360 23756 2372
rect 20180 2332 23756 2360
rect 17129 2323 17187 2329
rect 23750 2320 23756 2332
rect 23808 2320 23814 2372
rect 24486 2320 24492 2372
rect 24544 2360 24550 2372
rect 24857 2363 24915 2369
rect 24857 2360 24869 2363
rect 24544 2332 24869 2360
rect 24544 2320 24550 2332
rect 24857 2329 24869 2332
rect 24903 2329 24915 2363
rect 24857 2323 24915 2329
rect 26436 2304 26464 2400
rect 26973 2397 26985 2400
rect 27019 2397 27031 2431
rect 27172 2428 27200 2468
rect 27249 2465 27261 2499
rect 27295 2496 27307 2499
rect 28442 2496 28448 2508
rect 27295 2468 28448 2496
rect 27295 2465 27307 2468
rect 27249 2459 27307 2465
rect 28442 2456 28448 2468
rect 28500 2456 28506 2508
rect 30650 2496 30656 2508
rect 30611 2468 30656 2496
rect 30650 2456 30656 2468
rect 30708 2456 30714 2508
rect 34900 2496 34928 2527
rect 30760 2468 34928 2496
rect 29917 2431 29975 2437
rect 27172 2400 28764 2428
rect 26973 2391 27031 2397
rect 28350 2320 28356 2372
rect 28408 2360 28414 2372
rect 28629 2363 28687 2369
rect 28629 2360 28641 2363
rect 28408 2332 28641 2360
rect 28408 2320 28414 2332
rect 28629 2329 28641 2332
rect 28675 2329 28687 2363
rect 28736 2360 28764 2400
rect 29917 2397 29929 2431
rect 29963 2428 29975 2431
rect 30282 2428 30288 2440
rect 29963 2400 30288 2428
rect 29963 2397 29975 2400
rect 29917 2391 29975 2397
rect 30282 2388 30288 2400
rect 30340 2428 30346 2440
rect 30377 2431 30435 2437
rect 30377 2428 30389 2431
rect 30340 2400 30389 2428
rect 30340 2388 30346 2400
rect 30377 2397 30389 2400
rect 30423 2397 30435 2431
rect 30377 2391 30435 2397
rect 30760 2360 30788 2468
rect 32582 2428 32588 2440
rect 32543 2400 32588 2428
rect 32582 2388 32588 2400
rect 32640 2388 32646 2440
rect 34701 2431 34759 2437
rect 34701 2428 34713 2431
rect 34164 2400 34713 2428
rect 28736 2332 30788 2360
rect 28629 2323 28687 2329
rect 34164 2304 34192 2400
rect 34701 2397 34713 2400
rect 34747 2397 34759 2431
rect 37568 2428 37596 2527
rect 44174 2524 44180 2536
rect 44232 2524 44238 2576
rect 38105 2431 38163 2437
rect 38105 2428 38117 2431
rect 37568 2400 38117 2428
rect 34701 2391 34759 2397
rect 38105 2397 38117 2400
rect 38151 2397 38163 2431
rect 40034 2428 40040 2440
rect 39995 2400 40040 2428
rect 38105 2391 38163 2397
rect 40034 2388 40040 2400
rect 40092 2388 40098 2440
rect 42429 2431 42487 2437
rect 42429 2428 42441 2431
rect 41892 2400 42441 2428
rect 35713 2363 35771 2369
rect 35713 2329 35725 2363
rect 35759 2360 35771 2363
rect 36078 2360 36084 2372
rect 35759 2332 36084 2360
rect 35759 2329 35771 2332
rect 35713 2323 35771 2329
rect 36078 2320 36084 2332
rect 36136 2360 36142 2372
rect 36265 2363 36323 2369
rect 36265 2360 36277 2363
rect 36136 2332 36277 2360
rect 36136 2320 36142 2332
rect 36265 2329 36277 2332
rect 36311 2329 36323 2363
rect 36265 2323 36323 2329
rect 41892 2304 41920 2400
rect 42429 2397 42441 2400
rect 42475 2397 42487 2431
rect 42429 2391 42487 2397
rect 45278 2388 45284 2440
rect 45336 2428 45342 2440
rect 45833 2431 45891 2437
rect 45833 2428 45845 2431
rect 45336 2400 45845 2428
rect 45336 2388 45342 2400
rect 45833 2397 45845 2400
rect 45879 2397 45891 2431
rect 45833 2391 45891 2397
rect 46566 2388 46572 2440
rect 46624 2428 46630 2440
rect 46753 2431 46811 2437
rect 46753 2428 46765 2431
rect 46624 2400 46765 2428
rect 46624 2388 46630 2400
rect 46753 2397 46765 2400
rect 46799 2397 46811 2431
rect 47762 2428 47768 2440
rect 47723 2400 47768 2428
rect 46753 2391 46811 2397
rect 47762 2388 47768 2400
rect 47820 2388 47826 2440
rect 43441 2363 43499 2369
rect 43441 2329 43453 2363
rect 43487 2360 43499 2363
rect 43806 2360 43812 2372
rect 43487 2332 43812 2360
rect 43487 2329 43499 2332
rect 43441 2323 43499 2329
rect 43806 2320 43812 2332
rect 43864 2360 43870 2372
rect 43993 2363 44051 2369
rect 43993 2360 44005 2363
rect 43864 2332 44005 2360
rect 43864 2320 43870 2332
rect 43993 2329 44005 2332
rect 44039 2329 44051 2363
rect 43993 2323 44051 2329
rect 2314 2292 2320 2304
rect 2275 2264 2320 2292
rect 2314 2252 2320 2264
rect 2372 2252 2378 2304
rect 3234 2252 3240 2304
rect 3292 2292 3298 2304
rect 3881 2295 3939 2301
rect 3881 2292 3893 2295
rect 3292 2264 3893 2292
rect 3292 2252 3298 2264
rect 3881 2261 3893 2264
rect 3927 2261 3939 2295
rect 3881 2255 3939 2261
rect 10962 2252 10968 2304
rect 11020 2292 11026 2304
rect 11609 2295 11667 2301
rect 11609 2292 11621 2295
rect 11020 2264 11621 2292
rect 11020 2252 11026 2264
rect 11609 2261 11621 2264
rect 11655 2261 11667 2295
rect 11609 2255 11667 2261
rect 14826 2252 14832 2304
rect 14884 2292 14890 2304
rect 15013 2295 15071 2301
rect 15013 2292 15025 2295
rect 14884 2264 15025 2292
rect 14884 2252 14890 2264
rect 15013 2261 15025 2264
rect 15059 2261 15071 2295
rect 17218 2292 17224 2304
rect 17179 2264 17224 2292
rect 15013 2255 15071 2261
rect 17218 2252 17224 2264
rect 17276 2252 17282 2304
rect 24946 2292 24952 2304
rect 24907 2264 24952 2292
rect 24946 2252 24952 2264
rect 25004 2252 25010 2304
rect 26418 2292 26424 2304
rect 26379 2264 26424 2292
rect 26418 2252 26424 2264
rect 26476 2252 26482 2304
rect 32214 2252 32220 2304
rect 32272 2292 32278 2304
rect 32401 2295 32459 2301
rect 32401 2292 32413 2295
rect 32272 2264 32413 2292
rect 32272 2252 32278 2264
rect 32401 2261 32413 2264
rect 32447 2261 32459 2295
rect 34146 2292 34152 2304
rect 34107 2264 34152 2292
rect 32401 2255 32459 2261
rect 34146 2252 34152 2264
rect 34204 2252 34210 2304
rect 38010 2252 38016 2304
rect 38068 2292 38074 2304
rect 38289 2295 38347 2301
rect 38289 2292 38301 2295
rect 38068 2264 38301 2292
rect 38068 2252 38074 2264
rect 38289 2261 38301 2264
rect 38335 2261 38347 2295
rect 40218 2292 40224 2304
rect 40179 2264 40224 2292
rect 38289 2255 38347 2261
rect 40218 2252 40224 2264
rect 40276 2252 40282 2304
rect 41874 2292 41880 2304
rect 41835 2264 41880 2292
rect 41874 2252 41880 2264
rect 41932 2252 41938 2304
rect 42610 2292 42616 2304
rect 42571 2264 42616 2292
rect 42610 2252 42616 2264
rect 42668 2252 42674 2304
rect 45738 2252 45744 2304
rect 45796 2292 45802 2304
rect 46017 2295 46075 2301
rect 46017 2292 46029 2295
rect 45796 2264 46029 2292
rect 45796 2252 45802 2264
rect 46017 2261 46029 2264
rect 46063 2261 46075 2295
rect 46017 2255 46075 2261
rect 46842 2252 46848 2304
rect 46900 2292 46906 2304
rect 46937 2295 46995 2301
rect 46937 2292 46949 2295
rect 46900 2264 46949 2292
rect 46900 2252 46906 2264
rect 46937 2261 46949 2264
rect 46983 2261 46995 2295
rect 46937 2255 46995 2261
rect 47670 2252 47676 2304
rect 47728 2292 47734 2304
rect 47949 2295 48007 2301
rect 47949 2292 47961 2295
rect 47728 2264 47961 2292
rect 47728 2252 47734 2264
rect 47949 2261 47961 2264
rect 47995 2261 48007 2295
rect 47949 2255 48007 2261
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 2314 2048 2320 2100
rect 2372 2088 2378 2100
rect 32030 2088 32036 2100
rect 2372 2060 32036 2088
rect 2372 2048 2378 2060
rect 32030 2048 32036 2060
rect 32088 2048 32094 2100
rect 17218 1980 17224 2032
rect 17276 2020 17282 2032
rect 27154 2020 27160 2032
rect 17276 1992 27160 2020
rect 17276 1980 17282 1992
rect 27154 1980 27160 1992
rect 27212 1980 27218 2032
rect 42610 2020 42616 2032
rect 41386 1992 42616 2020
rect 24946 1912 24952 1964
rect 25004 1952 25010 1964
rect 33962 1952 33968 1964
rect 25004 1924 33968 1952
rect 25004 1912 25010 1924
rect 33962 1912 33968 1924
rect 34020 1912 34026 1964
rect 13354 1844 13360 1896
rect 13412 1884 13418 1896
rect 40218 1884 40224 1896
rect 13412 1856 40224 1884
rect 13412 1844 13418 1856
rect 40218 1844 40224 1856
rect 40276 1844 40282 1896
rect 20346 1776 20352 1828
rect 20404 1816 20410 1828
rect 41386 1816 41414 1992
rect 42610 1980 42616 1992
rect 42668 1980 42674 2032
rect 20404 1788 41414 1816
rect 20404 1776 20410 1788
<< via1 >>
rect 21088 47744 21140 47796
rect 30840 47744 30892 47796
rect 19156 47676 19208 47728
rect 29828 47676 29880 47728
rect 21180 47608 21232 47660
rect 26240 47608 26292 47660
rect 26424 47608 26476 47660
rect 32496 47608 32548 47660
rect 19616 47540 19668 47592
rect 37372 47608 37424 47660
rect 17224 47472 17276 47524
rect 22008 47472 22060 47524
rect 26240 47472 26292 47524
rect 26884 47472 26936 47524
rect 14280 47404 14332 47456
rect 40776 47404 40828 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 5816 47200 5868 47252
rect 13544 47200 13596 47252
rect 15476 47200 15528 47252
rect 15752 47200 15804 47252
rect 19616 47243 19668 47252
rect 9588 47132 9640 47184
rect 17224 47132 17276 47184
rect 19616 47209 19625 47243
rect 19625 47209 19659 47243
rect 19659 47209 19668 47243
rect 19616 47200 19668 47209
rect 21180 47243 21232 47252
rect 21180 47209 21189 47243
rect 21189 47209 21223 47243
rect 21223 47209 21232 47243
rect 21180 47200 21232 47209
rect 23204 47200 23256 47252
rect 26424 47243 26476 47252
rect 21088 47132 21140 47184
rect 9128 47064 9180 47116
rect 9772 47107 9824 47116
rect 9772 47073 9781 47107
rect 9781 47073 9815 47107
rect 9815 47073 9824 47107
rect 9772 47064 9824 47073
rect 12348 47064 12400 47116
rect 12532 47064 12584 47116
rect 14188 47064 14240 47116
rect 20 46860 72 46912
rect 2688 46996 2740 47048
rect 3976 47039 4028 47048
rect 3976 47005 3985 47039
rect 3985 47005 4019 47039
rect 4019 47005 4028 47039
rect 3976 46996 4028 47005
rect 6828 46996 6880 47048
rect 7840 47039 7892 47048
rect 7840 47005 7849 47039
rect 7849 47005 7883 47039
rect 7883 47005 7892 47039
rect 7840 46996 7892 47005
rect 11612 46996 11664 47048
rect 1952 46860 2004 46912
rect 2504 46860 2556 46912
rect 2872 46928 2924 46980
rect 9864 46928 9916 46980
rect 10876 46928 10928 46980
rect 14280 47039 14332 47048
rect 14280 47005 14289 47039
rect 14289 47005 14323 47039
rect 14323 47005 14332 47039
rect 14280 46996 14332 47005
rect 14740 47064 14792 47116
rect 16856 47064 16908 47116
rect 20260 47064 20312 47116
rect 15752 47039 15804 47048
rect 15752 47005 15761 47039
rect 15761 47005 15795 47039
rect 15795 47005 15804 47039
rect 15752 46996 15804 47005
rect 17040 47039 17092 47048
rect 8024 46903 8076 46912
rect 8024 46869 8033 46903
rect 8033 46869 8067 46903
rect 8067 46869 8076 46903
rect 8024 46860 8076 46869
rect 10416 46860 10468 46912
rect 14096 46903 14148 46912
rect 14096 46869 14105 46903
rect 14105 46869 14139 46903
rect 14139 46869 14148 46903
rect 14096 46860 14148 46869
rect 15292 46928 15344 46980
rect 17040 47005 17049 47039
rect 17049 47005 17083 47039
rect 17083 47005 17092 47039
rect 17040 46996 17092 47005
rect 19432 47039 19484 47048
rect 17408 46928 17460 46980
rect 19432 47005 19441 47039
rect 19441 47005 19475 47039
rect 19475 47005 19484 47039
rect 19432 46996 19484 47005
rect 21732 46996 21784 47048
rect 22192 47039 22244 47048
rect 22192 47005 22201 47039
rect 22201 47005 22235 47039
rect 22235 47005 22244 47039
rect 22192 46996 22244 47005
rect 26424 47209 26433 47243
rect 26433 47209 26467 47243
rect 26467 47209 26476 47243
rect 26424 47200 26476 47209
rect 34336 47200 34388 47252
rect 30840 47132 30892 47184
rect 33876 47132 33928 47184
rect 37280 47200 37332 47252
rect 38660 47200 38712 47252
rect 40592 47200 40644 47252
rect 40776 47243 40828 47252
rect 40776 47209 40785 47243
rect 40785 47209 40819 47243
rect 40819 47209 40828 47243
rect 40776 47200 40828 47209
rect 42800 47243 42852 47252
rect 42800 47209 42809 47243
rect 42809 47209 42843 47243
rect 42843 47209 42852 47243
rect 42800 47200 42852 47209
rect 46664 47243 46716 47252
rect 46664 47209 46673 47243
rect 46673 47209 46707 47243
rect 46707 47209 46716 47243
rect 46664 47200 46716 47209
rect 24400 47039 24452 47048
rect 24400 47005 24409 47039
rect 24409 47005 24443 47039
rect 24443 47005 24452 47039
rect 24400 46996 24452 47005
rect 24584 47039 24636 47048
rect 24584 47005 24593 47039
rect 24593 47005 24627 47039
rect 24627 47005 24636 47039
rect 24584 46996 24636 47005
rect 24952 46996 25004 47048
rect 28356 47064 28408 47116
rect 42432 47064 42484 47116
rect 29828 47039 29880 47048
rect 29828 47005 29837 47039
rect 29837 47005 29871 47039
rect 29871 47005 29880 47039
rect 29828 46996 29880 47005
rect 32128 47039 32180 47048
rect 32128 47005 32137 47039
rect 32137 47005 32171 47039
rect 32171 47005 32180 47039
rect 32128 46996 32180 47005
rect 20352 46971 20404 46980
rect 20352 46937 20361 46971
rect 20361 46937 20395 46971
rect 20395 46937 20404 46971
rect 20352 46928 20404 46937
rect 20996 46928 21048 46980
rect 21272 46928 21324 46980
rect 16488 46860 16540 46912
rect 20812 46860 20864 46912
rect 22284 46928 22336 46980
rect 28816 46928 28868 46980
rect 29184 46928 29236 46980
rect 31944 46928 31996 46980
rect 32496 46928 32548 46980
rect 38660 46996 38712 47048
rect 40592 46996 40644 47048
rect 46204 46996 46256 47048
rect 48320 46996 48372 47048
rect 35900 46928 35952 46980
rect 45468 46928 45520 46980
rect 26148 46860 26200 46912
rect 38752 46903 38804 46912
rect 38752 46869 38761 46903
rect 38761 46869 38795 46903
rect 38795 46869 38804 46903
rect 38752 46860 38804 46869
rect 44456 46860 44508 46912
rect 45192 46860 45244 46912
rect 47124 46928 47176 46980
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 2504 46699 2556 46708
rect 2504 46665 2513 46699
rect 2513 46665 2547 46699
rect 2547 46665 2556 46699
rect 2504 46656 2556 46665
rect 2688 46656 2740 46708
rect 10416 46699 10468 46708
rect 10416 46665 10425 46699
rect 10425 46665 10459 46699
rect 10459 46665 10468 46699
rect 10416 46656 10468 46665
rect 9588 46588 9640 46640
rect 12716 46588 12768 46640
rect 1400 46563 1452 46572
rect 1400 46529 1409 46563
rect 1409 46529 1443 46563
rect 1443 46529 1452 46563
rect 1400 46520 1452 46529
rect 19432 46656 19484 46708
rect 20904 46656 20956 46708
rect 24400 46699 24452 46708
rect 12992 46631 13044 46640
rect 12992 46597 13001 46631
rect 13001 46597 13035 46631
rect 13035 46597 13044 46631
rect 12992 46588 13044 46597
rect 10876 46452 10928 46504
rect 9864 46427 9916 46436
rect 9864 46393 9873 46427
rect 9873 46393 9907 46427
rect 9907 46393 9916 46427
rect 9864 46384 9916 46393
rect 10784 46384 10836 46436
rect 13176 46520 13228 46572
rect 13728 46563 13780 46572
rect 13728 46529 13737 46563
rect 13737 46529 13771 46563
rect 13771 46529 13780 46563
rect 13728 46520 13780 46529
rect 13820 46520 13872 46572
rect 14280 46520 14332 46572
rect 14740 46563 14792 46572
rect 14740 46529 14749 46563
rect 14749 46529 14783 46563
rect 14783 46529 14792 46563
rect 14740 46520 14792 46529
rect 15752 46588 15804 46640
rect 16948 46588 17000 46640
rect 12992 46452 13044 46504
rect 15292 46495 15344 46504
rect 14096 46384 14148 46436
rect 2688 46316 2740 46368
rect 6828 46359 6880 46368
rect 6828 46325 6837 46359
rect 6837 46325 6871 46359
rect 6871 46325 6880 46359
rect 6828 46316 6880 46325
rect 9312 46359 9364 46368
rect 9312 46325 9321 46359
rect 9321 46325 9355 46359
rect 9355 46325 9364 46359
rect 9312 46316 9364 46325
rect 12440 46359 12492 46368
rect 12440 46325 12449 46359
rect 12449 46325 12483 46359
rect 12483 46325 12492 46359
rect 12440 46316 12492 46325
rect 13452 46316 13504 46368
rect 15292 46461 15301 46495
rect 15301 46461 15335 46495
rect 15335 46461 15344 46495
rect 15292 46452 15344 46461
rect 16672 46520 16724 46572
rect 18052 46563 18104 46572
rect 18052 46529 18061 46563
rect 18061 46529 18095 46563
rect 18095 46529 18104 46563
rect 18052 46520 18104 46529
rect 18696 46520 18748 46572
rect 19340 46588 19392 46640
rect 21640 46588 21692 46640
rect 16764 46495 16816 46504
rect 16764 46461 16773 46495
rect 16773 46461 16807 46495
rect 16807 46461 16816 46495
rect 16764 46452 16816 46461
rect 18512 46452 18564 46504
rect 20076 46520 20128 46572
rect 20720 46520 20772 46572
rect 21180 46520 21232 46572
rect 21824 46520 21876 46572
rect 22100 46588 22152 46640
rect 24400 46665 24409 46699
rect 24409 46665 24443 46699
rect 24443 46665 24452 46699
rect 24400 46656 24452 46665
rect 24400 46520 24452 46572
rect 25964 46588 26016 46640
rect 24952 46563 25004 46572
rect 24952 46529 24961 46563
rect 24961 46529 24995 46563
rect 24995 46529 25004 46563
rect 24952 46520 25004 46529
rect 25228 46563 25280 46572
rect 25228 46529 25262 46563
rect 25262 46529 25280 46563
rect 25228 46520 25280 46529
rect 25504 46520 25556 46572
rect 22928 46495 22980 46504
rect 22928 46461 22937 46495
rect 22937 46461 22971 46495
rect 22971 46461 22980 46495
rect 22928 46452 22980 46461
rect 23572 46452 23624 46504
rect 26608 46520 26660 46572
rect 32864 46656 32916 46708
rect 42432 46699 42484 46708
rect 42432 46665 42441 46699
rect 42441 46665 42475 46699
rect 42475 46665 42484 46699
rect 42432 46656 42484 46665
rect 45192 46699 45244 46708
rect 45192 46665 45201 46699
rect 45201 46665 45235 46699
rect 45235 46665 45244 46699
rect 45192 46656 45244 46665
rect 18236 46384 18288 46436
rect 19984 46427 20036 46436
rect 19984 46393 19993 46427
rect 19993 46393 20027 46427
rect 20027 46393 20036 46427
rect 19984 46384 20036 46393
rect 22192 46384 22244 46436
rect 28356 46563 28408 46572
rect 28356 46529 28365 46563
rect 28365 46529 28399 46563
rect 28399 46529 28408 46563
rect 28356 46520 28408 46529
rect 34796 46588 34848 46640
rect 47216 46588 47268 46640
rect 49608 46588 49660 46640
rect 30932 46520 30984 46572
rect 31484 46520 31536 46572
rect 32128 46563 32180 46572
rect 32128 46529 32137 46563
rect 32137 46529 32171 46563
rect 32171 46529 32180 46563
rect 32128 46520 32180 46529
rect 33968 46520 34020 46572
rect 34060 46563 34112 46572
rect 34060 46529 34069 46563
rect 34069 46529 34103 46563
rect 34103 46529 34112 46563
rect 34060 46520 34112 46529
rect 48136 46520 48188 46572
rect 27988 46452 28040 46504
rect 43260 46452 43312 46504
rect 18420 46316 18472 46368
rect 20996 46316 21048 46368
rect 24584 46316 24636 46368
rect 26424 46316 26476 46368
rect 27436 46316 27488 46368
rect 31024 46384 31076 46436
rect 34704 46384 34756 46436
rect 46756 46427 46808 46436
rect 46756 46393 46765 46427
rect 46765 46393 46799 46427
rect 46799 46393 46808 46427
rect 46756 46384 46808 46393
rect 31300 46316 31352 46368
rect 31576 46359 31628 46368
rect 31576 46325 31585 46359
rect 31585 46325 31619 46359
rect 31619 46325 31628 46359
rect 31576 46316 31628 46325
rect 34428 46316 34480 46368
rect 35900 46359 35952 46368
rect 35900 46325 35909 46359
rect 35909 46325 35943 46359
rect 35943 46325 35952 46359
rect 35900 46316 35952 46325
rect 36820 46316 36872 46368
rect 46204 46359 46256 46368
rect 46204 46325 46213 46359
rect 46213 46325 46247 46359
rect 46247 46325 46256 46359
rect 46204 46316 46256 46325
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 1400 46112 1452 46164
rect 11612 46112 11664 46164
rect 12716 46112 12768 46164
rect 13452 46155 13504 46164
rect 13452 46121 13461 46155
rect 13461 46121 13495 46155
rect 13495 46121 13504 46155
rect 13452 46112 13504 46121
rect 9312 46044 9364 46096
rect 14188 46112 14240 46164
rect 18512 46112 18564 46164
rect 18696 46155 18748 46164
rect 18696 46121 18705 46155
rect 18705 46121 18739 46155
rect 18739 46121 18748 46155
rect 18696 46112 18748 46121
rect 23388 46112 23440 46164
rect 25964 46112 26016 46164
rect 31668 46112 31720 46164
rect 18420 46044 18472 46096
rect 13728 45976 13780 46028
rect 1676 45908 1728 45960
rect 2780 45908 2832 45960
rect 14096 45951 14148 45960
rect 14096 45917 14105 45951
rect 14105 45917 14139 45951
rect 14139 45917 14148 45951
rect 14096 45908 14148 45917
rect 14280 45951 14332 45960
rect 14280 45917 14289 45951
rect 14289 45917 14323 45951
rect 14323 45917 14332 45951
rect 14280 45908 14332 45917
rect 16488 45951 16540 45960
rect 16488 45917 16497 45951
rect 16497 45917 16531 45951
rect 16531 45917 16540 45951
rect 16488 45908 16540 45917
rect 16764 45951 16816 45960
rect 16764 45917 16773 45951
rect 16773 45917 16807 45951
rect 16807 45917 16816 45951
rect 16764 45908 16816 45917
rect 20904 46019 20956 46028
rect 20904 45985 20913 46019
rect 20913 45985 20947 46019
rect 20947 45985 20956 46019
rect 20904 45976 20956 45985
rect 22008 46019 22060 46028
rect 22008 45985 22017 46019
rect 22017 45985 22051 46019
rect 22051 45985 22060 46019
rect 22008 45976 22060 45985
rect 22192 45976 22244 46028
rect 13912 45840 13964 45892
rect 14464 45883 14516 45892
rect 14464 45849 14473 45883
rect 14473 45849 14507 45883
rect 14507 45849 14516 45883
rect 14464 45840 14516 45849
rect 16672 45883 16724 45892
rect 1952 45815 2004 45824
rect 1952 45781 1961 45815
rect 1961 45781 1995 45815
rect 1995 45781 2004 45815
rect 1952 45772 2004 45781
rect 10232 45815 10284 45824
rect 10232 45781 10241 45815
rect 10241 45781 10275 45815
rect 10275 45781 10284 45815
rect 10232 45772 10284 45781
rect 11704 45772 11756 45824
rect 11888 45815 11940 45824
rect 11888 45781 11897 45815
rect 11897 45781 11931 45815
rect 11931 45781 11940 45815
rect 11888 45772 11940 45781
rect 16028 45772 16080 45824
rect 16672 45849 16681 45883
rect 16681 45849 16715 45883
rect 16715 45849 16724 45883
rect 16672 45840 16724 45849
rect 18420 45840 18472 45892
rect 21916 45951 21968 45960
rect 21916 45917 21925 45951
rect 21925 45917 21959 45951
rect 21959 45917 21968 45951
rect 21916 45908 21968 45917
rect 22100 45908 22152 45960
rect 24492 45951 24544 45960
rect 24492 45917 24501 45951
rect 24501 45917 24535 45951
rect 24535 45917 24544 45951
rect 24492 45908 24544 45917
rect 18880 45840 18932 45892
rect 20168 45840 20220 45892
rect 23572 45883 23624 45892
rect 17684 45772 17736 45824
rect 18052 45772 18104 45824
rect 21456 45772 21508 45824
rect 22192 45815 22244 45824
rect 22192 45781 22201 45815
rect 22201 45781 22235 45815
rect 22235 45781 22244 45815
rect 22192 45772 22244 45781
rect 23572 45849 23581 45883
rect 23581 45849 23615 45883
rect 23615 45849 23624 45883
rect 23572 45840 23624 45849
rect 24492 45772 24544 45824
rect 31024 46044 31076 46096
rect 24952 45976 25004 46028
rect 28632 45976 28684 46028
rect 34060 46155 34112 46164
rect 24768 45908 24820 45960
rect 27068 45908 27120 45960
rect 29092 45908 29144 45960
rect 30288 45951 30340 45960
rect 30288 45917 30297 45951
rect 30297 45917 30331 45951
rect 30331 45917 30340 45951
rect 30288 45908 30340 45917
rect 32128 45951 32180 45960
rect 32128 45917 32137 45951
rect 32137 45917 32171 45951
rect 32171 45917 32180 45951
rect 32128 45908 32180 45917
rect 25136 45840 25188 45892
rect 31760 45840 31812 45892
rect 34060 46121 34069 46155
rect 34069 46121 34103 46155
rect 34103 46121 34112 46155
rect 34060 46112 34112 46121
rect 34796 46112 34848 46164
rect 48136 46112 48188 46164
rect 47216 46087 47268 46096
rect 47216 46053 47225 46087
rect 47225 46053 47259 46087
rect 47259 46053 47268 46087
rect 47216 46044 47268 46053
rect 48044 45951 48096 45960
rect 48044 45917 48053 45951
rect 48053 45917 48087 45951
rect 48087 45917 48096 45951
rect 48044 45908 48096 45917
rect 26148 45772 26200 45824
rect 26976 45815 27028 45824
rect 26976 45781 26985 45815
rect 26985 45781 27019 45815
rect 27019 45781 27028 45815
rect 26976 45772 27028 45781
rect 28540 45772 28592 45824
rect 30012 45772 30064 45824
rect 47032 45840 47084 45892
rect 46204 45772 46256 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 1676 45611 1728 45620
rect 1676 45577 1685 45611
rect 1685 45577 1719 45611
rect 1719 45577 1728 45611
rect 1676 45568 1728 45577
rect 1952 45568 2004 45620
rect 11152 45568 11204 45620
rect 9680 45543 9732 45552
rect 9680 45509 9689 45543
rect 9689 45509 9723 45543
rect 9723 45509 9732 45543
rect 9680 45500 9732 45509
rect 11888 45543 11940 45552
rect 11888 45509 11897 45543
rect 11897 45509 11931 45543
rect 11931 45509 11940 45543
rect 11888 45500 11940 45509
rect 12532 45543 12584 45552
rect 12532 45509 12541 45543
rect 12541 45509 12575 45543
rect 12575 45509 12584 45543
rect 12532 45500 12584 45509
rect 13912 45568 13964 45620
rect 16764 45568 16816 45620
rect 17684 45568 17736 45620
rect 12808 45432 12860 45484
rect 13268 45475 13320 45484
rect 13268 45441 13277 45475
rect 13277 45441 13311 45475
rect 13311 45441 13320 45475
rect 14464 45500 14516 45552
rect 13268 45432 13320 45441
rect 13912 45475 13964 45484
rect 13912 45441 13921 45475
rect 13921 45441 13955 45475
rect 13955 45441 13964 45475
rect 13912 45432 13964 45441
rect 16488 45432 16540 45484
rect 12992 45339 13044 45348
rect 12992 45305 13001 45339
rect 13001 45305 13035 45339
rect 13035 45305 13044 45339
rect 12992 45296 13044 45305
rect 17592 45475 17644 45484
rect 17592 45441 17601 45475
rect 17601 45441 17635 45475
rect 17635 45441 17644 45475
rect 17592 45432 17644 45441
rect 18236 45475 18288 45484
rect 18236 45441 18245 45475
rect 18245 45441 18279 45475
rect 18279 45441 18288 45475
rect 18236 45432 18288 45441
rect 18328 45475 18380 45484
rect 18328 45441 18337 45475
rect 18337 45441 18371 45475
rect 18371 45441 18380 45475
rect 18328 45432 18380 45441
rect 18604 45432 18656 45484
rect 18420 45364 18472 45416
rect 21732 45568 21784 45620
rect 22100 45568 22152 45620
rect 26148 45611 26200 45620
rect 20720 45500 20772 45552
rect 20996 45500 21048 45552
rect 21640 45500 21692 45552
rect 22192 45543 22244 45552
rect 22192 45509 22201 45543
rect 22201 45509 22235 45543
rect 22235 45509 22244 45543
rect 22192 45500 22244 45509
rect 22928 45500 22980 45552
rect 20812 45432 20864 45484
rect 21088 45475 21140 45484
rect 21088 45441 21097 45475
rect 21097 45441 21131 45475
rect 21131 45441 21140 45475
rect 21088 45432 21140 45441
rect 22284 45475 22336 45484
rect 22284 45441 22293 45475
rect 22293 45441 22327 45475
rect 22327 45441 22336 45475
rect 26148 45577 26157 45611
rect 26157 45577 26191 45611
rect 26191 45577 26200 45611
rect 26148 45568 26200 45577
rect 26792 45568 26844 45620
rect 28632 45568 28684 45620
rect 29000 45568 29052 45620
rect 30380 45568 30432 45620
rect 31484 45611 31536 45620
rect 23204 45500 23256 45552
rect 31484 45577 31493 45611
rect 31493 45577 31527 45611
rect 31527 45577 31536 45611
rect 31484 45568 31536 45577
rect 31668 45568 31720 45620
rect 38752 45568 38804 45620
rect 48044 45611 48096 45620
rect 48044 45577 48053 45611
rect 48053 45577 48087 45611
rect 48087 45577 48096 45611
rect 48044 45568 48096 45577
rect 22284 45432 22336 45441
rect 23572 45432 23624 45484
rect 24492 45432 24544 45484
rect 20996 45364 21048 45416
rect 21824 45407 21876 45416
rect 21824 45373 21833 45407
rect 21833 45373 21867 45407
rect 21867 45373 21876 45407
rect 21824 45364 21876 45373
rect 22008 45364 22060 45416
rect 24032 45407 24084 45416
rect 24032 45373 24041 45407
rect 24041 45373 24075 45407
rect 24075 45373 24084 45407
rect 24032 45364 24084 45373
rect 24400 45364 24452 45416
rect 25044 45364 25096 45416
rect 14464 45296 14516 45348
rect 16580 45296 16632 45348
rect 19156 45296 19208 45348
rect 19340 45296 19392 45348
rect 10416 45271 10468 45280
rect 10416 45237 10425 45271
rect 10425 45237 10459 45271
rect 10459 45237 10468 45271
rect 10416 45228 10468 45237
rect 12164 45228 12216 45280
rect 12624 45228 12676 45280
rect 16028 45228 16080 45280
rect 20444 45271 20496 45280
rect 20444 45237 20453 45271
rect 20453 45237 20487 45271
rect 20487 45237 20496 45271
rect 20444 45228 20496 45237
rect 21180 45296 21232 45348
rect 24860 45296 24912 45348
rect 23204 45228 23256 45280
rect 23480 45271 23532 45280
rect 23480 45237 23489 45271
rect 23489 45237 23523 45271
rect 23523 45237 23532 45271
rect 23480 45228 23532 45237
rect 23940 45228 23992 45280
rect 25964 45475 26016 45484
rect 25964 45441 25973 45475
rect 25973 45441 26007 45475
rect 26007 45441 26016 45475
rect 25964 45432 26016 45441
rect 26240 45475 26292 45484
rect 26240 45441 26249 45475
rect 26249 45441 26283 45475
rect 26283 45441 26292 45475
rect 26240 45432 26292 45441
rect 26976 45432 27028 45484
rect 29644 45475 29696 45484
rect 29644 45441 29653 45475
rect 29653 45441 29687 45475
rect 29687 45441 29696 45475
rect 29644 45432 29696 45441
rect 32128 45432 32180 45484
rect 33232 45475 33284 45484
rect 33876 45500 33928 45552
rect 33232 45441 33250 45475
rect 33250 45441 33284 45475
rect 33232 45432 33284 45441
rect 34612 45475 34664 45484
rect 34612 45441 34621 45475
rect 34621 45441 34655 45475
rect 34655 45441 34664 45475
rect 34612 45432 34664 45441
rect 31024 45364 31076 45416
rect 35532 45364 35584 45416
rect 27160 45296 27212 45348
rect 28356 45271 28408 45280
rect 28356 45237 28365 45271
rect 28365 45237 28399 45271
rect 28399 45237 28408 45271
rect 28356 45228 28408 45237
rect 32036 45296 32088 45348
rect 43260 45296 43312 45348
rect 33876 45228 33928 45280
rect 34060 45271 34112 45280
rect 34060 45237 34069 45271
rect 34069 45237 34103 45271
rect 34103 45237 34112 45271
rect 34060 45228 34112 45237
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 13268 45024 13320 45076
rect 14280 45024 14332 45076
rect 17040 45024 17092 45076
rect 20536 45024 20588 45076
rect 21640 45024 21692 45076
rect 22100 45067 22152 45076
rect 22100 45033 22109 45067
rect 22109 45033 22143 45067
rect 22143 45033 22152 45067
rect 22100 45024 22152 45033
rect 24032 45024 24084 45076
rect 24584 45024 24636 45076
rect 25964 45024 26016 45076
rect 22192 44956 22244 45008
rect 23480 44956 23532 45008
rect 14004 44888 14056 44940
rect 16580 44931 16632 44940
rect 10232 44820 10284 44872
rect 12808 44863 12860 44872
rect 6828 44752 6880 44804
rect 10876 44752 10928 44804
rect 12440 44752 12492 44804
rect 12808 44829 12817 44863
rect 12817 44829 12851 44863
rect 12851 44829 12860 44863
rect 12808 44820 12860 44829
rect 13268 44820 13320 44872
rect 13360 44820 13412 44872
rect 16580 44897 16589 44931
rect 16589 44897 16623 44931
rect 16623 44897 16632 44931
rect 16580 44888 16632 44897
rect 17040 44931 17092 44940
rect 17040 44897 17049 44931
rect 17049 44897 17083 44931
rect 17083 44897 17092 44931
rect 17040 44888 17092 44897
rect 20444 44888 20496 44940
rect 21640 44931 21692 44940
rect 14740 44820 14792 44872
rect 15108 44820 15160 44872
rect 15476 44863 15528 44872
rect 15476 44829 15485 44863
rect 15485 44829 15519 44863
rect 15519 44829 15528 44863
rect 15476 44820 15528 44829
rect 13820 44752 13872 44804
rect 14648 44752 14700 44804
rect 16488 44820 16540 44872
rect 19248 44863 19300 44872
rect 19248 44829 19257 44863
rect 19257 44829 19291 44863
rect 19291 44829 19300 44863
rect 19248 44820 19300 44829
rect 20536 44863 20588 44872
rect 20536 44829 20545 44863
rect 20545 44829 20579 44863
rect 20579 44829 20588 44863
rect 20536 44820 20588 44829
rect 20904 44863 20956 44872
rect 20904 44829 20913 44863
rect 20913 44829 20947 44863
rect 20947 44829 20956 44863
rect 20904 44820 20956 44829
rect 21640 44897 21649 44931
rect 21649 44897 21683 44931
rect 21683 44897 21692 44931
rect 21640 44888 21692 44897
rect 22008 44888 22060 44940
rect 25780 44956 25832 45008
rect 27068 44931 27120 44940
rect 21732 44863 21784 44872
rect 21732 44829 21741 44863
rect 21741 44829 21775 44863
rect 21775 44829 21784 44863
rect 21732 44820 21784 44829
rect 22284 44820 22336 44872
rect 9864 44684 9916 44736
rect 11244 44727 11296 44736
rect 11244 44693 11253 44727
rect 11253 44693 11287 44727
rect 11287 44693 11296 44727
rect 11244 44684 11296 44693
rect 16028 44684 16080 44736
rect 17960 44684 18012 44736
rect 19156 44684 19208 44736
rect 19340 44727 19392 44736
rect 19340 44693 19349 44727
rect 19349 44693 19383 44727
rect 19383 44693 19392 44727
rect 19340 44684 19392 44693
rect 20720 44684 20772 44736
rect 23204 44752 23256 44804
rect 25044 44863 25096 44872
rect 25044 44829 25053 44863
rect 25053 44829 25087 44863
rect 25087 44829 25096 44863
rect 25044 44820 25096 44829
rect 26056 44820 26108 44872
rect 27068 44897 27077 44931
rect 27077 44897 27111 44931
rect 27111 44897 27120 44931
rect 27068 44888 27120 44897
rect 30932 45024 30984 45076
rect 31024 45024 31076 45076
rect 47952 45024 48004 45076
rect 48136 45067 48188 45076
rect 48136 45033 48145 45067
rect 48145 45033 48179 45067
rect 48179 45033 48188 45067
rect 48136 45024 48188 45033
rect 20996 44684 21048 44736
rect 22008 44684 22060 44736
rect 23480 44684 23532 44736
rect 23756 44727 23808 44736
rect 23756 44693 23765 44727
rect 23765 44693 23799 44727
rect 23799 44693 23808 44727
rect 23756 44684 23808 44693
rect 25780 44684 25832 44736
rect 27528 44752 27580 44804
rect 28080 44684 28132 44736
rect 30656 44820 30708 44872
rect 32036 44888 32088 44940
rect 34704 44888 34756 44940
rect 33784 44820 33836 44872
rect 34060 44820 34112 44872
rect 29276 44752 29328 44804
rect 34612 44752 34664 44804
rect 32312 44684 32364 44736
rect 33876 44684 33928 44736
rect 35440 44684 35492 44736
rect 36084 44727 36136 44736
rect 36084 44693 36093 44727
rect 36093 44693 36127 44727
rect 36127 44693 36136 44727
rect 36084 44684 36136 44693
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 10416 44480 10468 44532
rect 12624 44480 12676 44532
rect 12808 44480 12860 44532
rect 13268 44523 13320 44532
rect 13268 44489 13277 44523
rect 13277 44489 13311 44523
rect 13311 44489 13320 44523
rect 13268 44480 13320 44489
rect 16028 44523 16080 44532
rect 16028 44489 16037 44523
rect 16037 44489 16071 44523
rect 16071 44489 16080 44523
rect 16028 44480 16080 44489
rect 16304 44412 16356 44464
rect 19248 44480 19300 44532
rect 21732 44480 21784 44532
rect 22284 44480 22336 44532
rect 23756 44480 23808 44532
rect 33968 44480 34020 44532
rect 34428 44480 34480 44532
rect 47952 44523 48004 44532
rect 1400 44387 1452 44396
rect 1400 44353 1409 44387
rect 1409 44353 1443 44387
rect 1443 44353 1452 44387
rect 1400 44344 1452 44353
rect 9864 44344 9916 44396
rect 13268 44344 13320 44396
rect 12164 44276 12216 44328
rect 14004 44344 14056 44396
rect 15108 44344 15160 44396
rect 15292 44344 15344 44396
rect 15476 44344 15528 44396
rect 17500 44387 17552 44396
rect 17500 44353 17509 44387
rect 17509 44353 17543 44387
rect 17543 44353 17552 44387
rect 17500 44344 17552 44353
rect 18052 44387 18104 44396
rect 18052 44353 18061 44387
rect 18061 44353 18095 44387
rect 18095 44353 18104 44387
rect 18052 44344 18104 44353
rect 18144 44387 18196 44396
rect 18144 44353 18153 44387
rect 18153 44353 18187 44387
rect 18187 44353 18196 44387
rect 18144 44344 18196 44353
rect 19248 44387 19300 44396
rect 13452 44276 13504 44328
rect 15016 44276 15068 44328
rect 16488 44276 16540 44328
rect 18972 44319 19024 44328
rect 18972 44285 18981 44319
rect 18981 44285 19015 44319
rect 19015 44285 19024 44319
rect 18972 44276 19024 44285
rect 19248 44353 19257 44387
rect 19257 44353 19291 44387
rect 19291 44353 19300 44387
rect 19248 44344 19300 44353
rect 24768 44412 24820 44464
rect 25320 44412 25372 44464
rect 20168 44344 20220 44396
rect 20720 44387 20772 44396
rect 20720 44353 20729 44387
rect 20729 44353 20763 44387
rect 20763 44353 20772 44387
rect 20720 44344 20772 44353
rect 12440 44208 12492 44260
rect 20352 44276 20404 44328
rect 21180 44344 21232 44396
rect 21824 44387 21876 44396
rect 21824 44353 21833 44387
rect 21833 44353 21867 44387
rect 21867 44353 21876 44387
rect 21824 44344 21876 44353
rect 22008 44387 22060 44396
rect 22008 44353 22017 44387
rect 22017 44353 22051 44387
rect 22051 44353 22060 44387
rect 22008 44344 22060 44353
rect 23756 44387 23808 44396
rect 23756 44353 23765 44387
rect 23765 44353 23799 44387
rect 23799 44353 23808 44387
rect 23756 44344 23808 44353
rect 23940 44387 23992 44396
rect 23940 44353 23949 44387
rect 23949 44353 23983 44387
rect 23983 44353 23992 44387
rect 23940 44344 23992 44353
rect 24860 44344 24912 44396
rect 27896 44344 27948 44396
rect 32036 44412 32088 44464
rect 33324 44387 33376 44396
rect 22284 44319 22336 44328
rect 22284 44285 22293 44319
rect 22293 44285 22327 44319
rect 22327 44285 22336 44319
rect 22284 44276 22336 44285
rect 23112 44276 23164 44328
rect 23480 44276 23532 44328
rect 24768 44319 24820 44328
rect 24768 44285 24777 44319
rect 24777 44285 24811 44319
rect 24811 44285 24820 44319
rect 24768 44276 24820 44285
rect 25504 44208 25556 44260
rect 25596 44208 25648 44260
rect 1676 44140 1728 44192
rect 9864 44140 9916 44192
rect 10968 44183 11020 44192
rect 10968 44149 10977 44183
rect 10977 44149 11011 44183
rect 11011 44149 11020 44183
rect 10968 44140 11020 44149
rect 14096 44183 14148 44192
rect 14096 44149 14105 44183
rect 14105 44149 14139 44183
rect 14139 44149 14148 44183
rect 14096 44140 14148 44149
rect 18236 44140 18288 44192
rect 20812 44183 20864 44192
rect 20812 44149 20821 44183
rect 20821 44149 20855 44183
rect 20855 44149 20864 44183
rect 20812 44140 20864 44149
rect 21640 44140 21692 44192
rect 22928 44140 22980 44192
rect 23940 44183 23992 44192
rect 23940 44149 23949 44183
rect 23949 44149 23983 44183
rect 23983 44149 23992 44183
rect 23940 44140 23992 44149
rect 24400 44183 24452 44192
rect 24400 44149 24409 44183
rect 24409 44149 24443 44183
rect 24443 44149 24452 44183
rect 24400 44140 24452 44149
rect 25044 44140 25096 44192
rect 26056 44183 26108 44192
rect 26056 44149 26065 44183
rect 26065 44149 26099 44183
rect 26099 44149 26108 44183
rect 26056 44140 26108 44149
rect 33324 44353 33342 44387
rect 33342 44353 33376 44387
rect 33324 44344 33376 44353
rect 34704 44344 34756 44396
rect 35440 44387 35492 44396
rect 35440 44353 35449 44387
rect 35449 44353 35483 44387
rect 35483 44353 35492 44387
rect 35440 44344 35492 44353
rect 35532 44387 35584 44396
rect 35532 44353 35541 44387
rect 35541 44353 35575 44387
rect 35575 44353 35584 44387
rect 35532 44344 35584 44353
rect 29000 44319 29052 44328
rect 29000 44285 29009 44319
rect 29009 44285 29043 44319
rect 29043 44285 29052 44319
rect 29000 44276 29052 44285
rect 31484 44276 31536 44328
rect 34796 44319 34848 44328
rect 34796 44285 34805 44319
rect 34805 44285 34839 44319
rect 34839 44285 34848 44319
rect 34796 44276 34848 44285
rect 35900 44208 35952 44260
rect 47952 44489 47961 44523
rect 47961 44489 47995 44523
rect 47995 44489 48004 44523
rect 47952 44480 48004 44489
rect 48044 44387 48096 44396
rect 48044 44353 48053 44387
rect 48053 44353 48087 44387
rect 48087 44353 48096 44387
rect 48044 44344 48096 44353
rect 29000 44140 29052 44192
rect 30472 44140 30524 44192
rect 33600 44140 33652 44192
rect 35348 44140 35400 44192
rect 36728 44183 36780 44192
rect 36728 44149 36737 44183
rect 36737 44149 36771 44183
rect 36771 44149 36780 44183
rect 36728 44140 36780 44149
rect 37280 44140 37332 44192
rect 37740 44140 37792 44192
rect 37924 44183 37976 44192
rect 37924 44149 37933 44183
rect 37933 44149 37967 44183
rect 37967 44149 37976 44183
rect 37924 44140 37976 44149
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 1400 43979 1452 43988
rect 1400 43945 1409 43979
rect 1409 43945 1443 43979
rect 1443 43945 1452 43979
rect 1400 43936 1452 43945
rect 11704 43936 11756 43988
rect 14096 43936 14148 43988
rect 14464 43979 14516 43988
rect 14464 43945 14473 43979
rect 14473 43945 14507 43979
rect 14507 43945 14516 43979
rect 14464 43936 14516 43945
rect 16028 43936 16080 43988
rect 17960 43936 18012 43988
rect 18972 43936 19024 43988
rect 15108 43868 15160 43920
rect 13084 43843 13136 43852
rect 13084 43809 13093 43843
rect 13093 43809 13127 43843
rect 13127 43809 13136 43843
rect 13084 43800 13136 43809
rect 14832 43800 14884 43852
rect 17868 43800 17920 43852
rect 20536 43936 20588 43988
rect 20628 43936 20680 43988
rect 10876 43775 10928 43784
rect 10876 43741 10885 43775
rect 10885 43741 10919 43775
rect 10919 43741 10928 43775
rect 10876 43732 10928 43741
rect 10968 43664 11020 43716
rect 12808 43732 12860 43784
rect 12900 43732 12952 43784
rect 14924 43775 14976 43784
rect 14924 43741 14933 43775
rect 14933 43741 14967 43775
rect 14967 43741 14976 43775
rect 14924 43732 14976 43741
rect 15200 43732 15252 43784
rect 16304 43775 16356 43784
rect 16304 43741 16313 43775
rect 16313 43741 16347 43775
rect 16347 43741 16356 43775
rect 16304 43732 16356 43741
rect 16488 43775 16540 43784
rect 16488 43741 16497 43775
rect 16497 43741 16531 43775
rect 16531 43741 16540 43775
rect 16488 43732 16540 43741
rect 16580 43732 16632 43784
rect 18236 43775 18288 43784
rect 18236 43741 18245 43775
rect 18245 43741 18279 43775
rect 18279 43741 18288 43775
rect 18236 43732 18288 43741
rect 20812 43868 20864 43920
rect 24768 43911 24820 43920
rect 21180 43800 21232 43852
rect 22008 43800 22060 43852
rect 21548 43775 21600 43784
rect 15660 43664 15712 43716
rect 21548 43741 21557 43775
rect 21557 43741 21591 43775
rect 21591 43741 21600 43775
rect 21548 43732 21600 43741
rect 22284 43775 22336 43784
rect 18696 43707 18748 43716
rect 18696 43673 18705 43707
rect 18705 43673 18739 43707
rect 18739 43673 18748 43707
rect 18696 43664 18748 43673
rect 19432 43664 19484 43716
rect 9864 43596 9916 43648
rect 11796 43596 11848 43648
rect 15568 43596 15620 43648
rect 19984 43596 20036 43648
rect 20720 43596 20772 43648
rect 21272 43664 21324 43716
rect 22284 43741 22293 43775
rect 22293 43741 22327 43775
rect 22327 43741 22336 43775
rect 22284 43732 22336 43741
rect 22744 43732 22796 43784
rect 23388 43732 23440 43784
rect 24768 43877 24777 43911
rect 24777 43877 24811 43911
rect 24811 43877 24820 43911
rect 24768 43868 24820 43877
rect 25504 43936 25556 43988
rect 26976 43868 27028 43920
rect 34796 43936 34848 43988
rect 48044 43979 48096 43988
rect 48044 43945 48053 43979
rect 48053 43945 48087 43979
rect 48087 43945 48096 43979
rect 48044 43936 48096 43945
rect 24492 43800 24544 43852
rect 27068 43800 27120 43852
rect 24952 43732 25004 43784
rect 26976 43732 27028 43784
rect 34060 43800 34112 43852
rect 29368 43732 29420 43784
rect 34612 43732 34664 43784
rect 22192 43664 22244 43716
rect 22836 43664 22888 43716
rect 24124 43664 24176 43716
rect 24860 43664 24912 43716
rect 21456 43596 21508 43648
rect 22100 43596 22152 43648
rect 22468 43596 22520 43648
rect 23204 43596 23256 43648
rect 23756 43596 23808 43648
rect 29184 43664 29236 43716
rect 35348 43800 35400 43852
rect 36176 43800 36228 43852
rect 35164 43775 35216 43784
rect 35164 43741 35173 43775
rect 35173 43741 35207 43775
rect 35207 43741 35216 43775
rect 35164 43732 35216 43741
rect 35624 43775 35676 43784
rect 35624 43741 35633 43775
rect 35633 43741 35667 43775
rect 35667 43741 35676 43775
rect 35624 43732 35676 43741
rect 35532 43664 35584 43716
rect 35992 43664 36044 43716
rect 36268 43732 36320 43784
rect 37924 43732 37976 43784
rect 27620 43596 27672 43648
rect 28724 43639 28776 43648
rect 28724 43605 28733 43639
rect 28733 43605 28767 43639
rect 28767 43605 28776 43639
rect 28724 43596 28776 43605
rect 30564 43596 30616 43648
rect 32036 43596 32088 43648
rect 33140 43596 33192 43648
rect 34060 43596 34112 43648
rect 36452 43707 36504 43716
rect 36452 43673 36461 43707
rect 36461 43673 36495 43707
rect 36495 43673 36504 43707
rect 36636 43707 36688 43716
rect 36452 43664 36504 43673
rect 36636 43673 36645 43707
rect 36645 43673 36679 43707
rect 36679 43673 36688 43707
rect 36636 43664 36688 43673
rect 37740 43707 37792 43716
rect 37740 43673 37749 43707
rect 37749 43673 37783 43707
rect 37783 43673 37792 43707
rect 37740 43664 37792 43673
rect 37832 43596 37884 43648
rect 38384 43639 38436 43648
rect 38384 43605 38393 43639
rect 38393 43605 38427 43639
rect 38427 43605 38436 43639
rect 38384 43596 38436 43605
rect 38568 43596 38620 43648
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 10784 43392 10836 43444
rect 12900 43435 12952 43444
rect 12900 43401 12909 43435
rect 12909 43401 12943 43435
rect 12943 43401 12952 43435
rect 12900 43392 12952 43401
rect 13084 43392 13136 43444
rect 13912 43435 13964 43444
rect 10968 43324 11020 43376
rect 12992 43256 13044 43308
rect 13912 43401 13921 43435
rect 13921 43401 13955 43435
rect 13955 43401 13964 43435
rect 13912 43392 13964 43401
rect 15200 43392 15252 43444
rect 13452 43231 13504 43240
rect 12624 43120 12676 43172
rect 13452 43197 13461 43231
rect 13461 43197 13495 43231
rect 13495 43197 13504 43231
rect 13452 43188 13504 43197
rect 13360 43120 13412 43172
rect 14924 43188 14976 43240
rect 15660 43231 15712 43240
rect 15660 43197 15669 43231
rect 15669 43197 15703 43231
rect 15703 43197 15712 43231
rect 15660 43188 15712 43197
rect 16764 43256 16816 43308
rect 16948 43256 17000 43308
rect 17040 43256 17092 43308
rect 17960 43324 18012 43376
rect 19248 43392 19300 43444
rect 21548 43392 21600 43444
rect 28080 43435 28132 43444
rect 17684 43299 17736 43308
rect 17684 43265 17693 43299
rect 17693 43265 17727 43299
rect 17727 43265 17736 43299
rect 17684 43256 17736 43265
rect 18328 43299 18380 43308
rect 18328 43265 18337 43299
rect 18337 43265 18371 43299
rect 18371 43265 18380 43299
rect 18328 43256 18380 43265
rect 18512 43299 18564 43308
rect 18512 43265 18521 43299
rect 18521 43265 18555 43299
rect 18555 43265 18564 43299
rect 18512 43256 18564 43265
rect 17868 43231 17920 43240
rect 17868 43197 17877 43231
rect 17877 43197 17911 43231
rect 17911 43197 17920 43231
rect 17868 43188 17920 43197
rect 20628 43324 20680 43376
rect 20812 43324 20864 43376
rect 20720 43299 20772 43308
rect 20720 43265 20729 43299
rect 20729 43265 20763 43299
rect 20763 43265 20772 43299
rect 20720 43256 20772 43265
rect 22008 43299 22060 43308
rect 19432 43188 19484 43240
rect 15844 43120 15896 43172
rect 17960 43120 18012 43172
rect 18604 43120 18656 43172
rect 19984 43188 20036 43240
rect 20352 43188 20404 43240
rect 22008 43265 22017 43299
rect 22017 43265 22051 43299
rect 22051 43265 22060 43299
rect 22008 43256 22060 43265
rect 23756 43324 23808 43376
rect 23388 43299 23440 43308
rect 23388 43265 23397 43299
rect 23397 43265 23431 43299
rect 23431 43265 23440 43299
rect 23388 43256 23440 43265
rect 24032 43299 24084 43308
rect 24032 43265 24041 43299
rect 24041 43265 24075 43299
rect 24075 43265 24084 43299
rect 24032 43256 24084 43265
rect 24768 43324 24820 43376
rect 27252 43324 27304 43376
rect 28080 43401 28089 43435
rect 28089 43401 28123 43435
rect 28123 43401 28132 43435
rect 28080 43392 28132 43401
rect 29000 43392 29052 43444
rect 29184 43392 29236 43444
rect 33324 43392 33376 43444
rect 34520 43392 34572 43444
rect 35900 43392 35952 43444
rect 30380 43367 30432 43376
rect 30380 43333 30389 43367
rect 30389 43333 30423 43367
rect 30423 43333 30432 43367
rect 30380 43324 30432 43333
rect 32036 43324 32088 43376
rect 26332 43256 26384 43308
rect 27068 43256 27120 43308
rect 33324 43299 33376 43308
rect 33692 43324 33744 43376
rect 35532 43324 35584 43376
rect 33324 43265 33342 43299
rect 33342 43265 33376 43299
rect 33324 43256 33376 43265
rect 35624 43256 35676 43308
rect 37832 43256 37884 43308
rect 38292 43256 38344 43308
rect 38384 43299 38436 43308
rect 38384 43265 38393 43299
rect 38393 43265 38427 43299
rect 38427 43265 38436 43299
rect 38384 43256 38436 43265
rect 38568 43299 38620 43308
rect 38568 43265 38577 43299
rect 38577 43265 38611 43299
rect 38611 43265 38620 43299
rect 38568 43256 38620 43265
rect 24492 43188 24544 43240
rect 26976 43231 27028 43240
rect 26976 43197 26985 43231
rect 26985 43197 27019 43231
rect 27019 43197 27028 43231
rect 26976 43188 27028 43197
rect 35992 43188 36044 43240
rect 36728 43188 36780 43240
rect 24400 43120 24452 43172
rect 14188 43052 14240 43104
rect 16672 43052 16724 43104
rect 19984 43052 20036 43104
rect 21916 43052 21968 43104
rect 25412 43052 25464 43104
rect 27620 43095 27672 43104
rect 27620 43061 27629 43095
rect 27629 43061 27663 43095
rect 27663 43061 27672 43095
rect 27620 43052 27672 43061
rect 30840 43095 30892 43104
rect 30840 43061 30849 43095
rect 30849 43061 30883 43095
rect 30883 43061 30892 43095
rect 30840 43052 30892 43061
rect 32220 43095 32272 43104
rect 32220 43061 32229 43095
rect 32229 43061 32263 43095
rect 32263 43061 32272 43095
rect 32220 43052 32272 43061
rect 35164 43052 35216 43104
rect 35900 43120 35952 43172
rect 36636 43120 36688 43172
rect 39948 43120 40000 43172
rect 38016 43052 38068 43104
rect 38292 43052 38344 43104
rect 39120 43095 39172 43104
rect 39120 43061 39129 43095
rect 39129 43061 39163 43095
rect 39163 43061 39172 43095
rect 39120 43052 39172 43061
rect 40224 43052 40276 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 10968 42848 11020 42900
rect 13084 42848 13136 42900
rect 15660 42848 15712 42900
rect 18512 42848 18564 42900
rect 19524 42848 19576 42900
rect 12624 42780 12676 42832
rect 16580 42780 16632 42832
rect 9588 42712 9640 42764
rect 10784 42644 10836 42696
rect 11244 42644 11296 42696
rect 12256 42644 12308 42696
rect 12900 42712 12952 42764
rect 12992 42644 13044 42696
rect 13544 42755 13596 42764
rect 13544 42721 13553 42755
rect 13553 42721 13587 42755
rect 13587 42721 13596 42755
rect 15844 42755 15896 42764
rect 13544 42712 13596 42721
rect 14832 42687 14884 42696
rect 14832 42653 14841 42687
rect 14841 42653 14875 42687
rect 14875 42653 14884 42687
rect 14832 42644 14884 42653
rect 15568 42687 15620 42696
rect 15568 42653 15577 42687
rect 15577 42653 15611 42687
rect 15611 42653 15620 42687
rect 15568 42644 15620 42653
rect 15844 42721 15853 42755
rect 15853 42721 15887 42755
rect 15887 42721 15896 42755
rect 15844 42712 15896 42721
rect 16764 42712 16816 42764
rect 20720 42848 20772 42900
rect 21640 42891 21692 42900
rect 21640 42857 21649 42891
rect 21649 42857 21683 42891
rect 21683 42857 21692 42891
rect 21640 42848 21692 42857
rect 23204 42848 23256 42900
rect 31484 42848 31536 42900
rect 34060 42848 34112 42900
rect 39948 42848 40000 42900
rect 20352 42755 20404 42764
rect 20352 42721 20361 42755
rect 20361 42721 20395 42755
rect 20395 42721 20404 42755
rect 20352 42712 20404 42721
rect 16856 42644 16908 42696
rect 17960 42687 18012 42696
rect 17960 42653 17969 42687
rect 17969 42653 18003 42687
rect 18003 42653 18012 42687
rect 17960 42644 18012 42653
rect 18144 42687 18196 42696
rect 18144 42653 18153 42687
rect 18153 42653 18187 42687
rect 18187 42653 18196 42687
rect 18144 42644 18196 42653
rect 19340 42687 19392 42696
rect 19340 42653 19349 42687
rect 19349 42653 19383 42687
rect 19383 42653 19392 42687
rect 19340 42644 19392 42653
rect 1492 42551 1544 42560
rect 1492 42517 1501 42551
rect 1501 42517 1535 42551
rect 1535 42517 1544 42551
rect 1492 42508 1544 42517
rect 9588 42551 9640 42560
rect 9588 42517 9597 42551
rect 9597 42517 9631 42551
rect 9631 42517 9640 42551
rect 9588 42508 9640 42517
rect 10784 42508 10836 42560
rect 11796 42551 11848 42560
rect 11796 42517 11805 42551
rect 11805 42517 11839 42551
rect 11839 42517 11848 42551
rect 11796 42508 11848 42517
rect 14924 42576 14976 42628
rect 12900 42508 12952 42560
rect 13820 42508 13872 42560
rect 17132 42619 17184 42628
rect 17132 42585 17141 42619
rect 17141 42585 17175 42619
rect 17175 42585 17184 42619
rect 17132 42576 17184 42585
rect 18512 42576 18564 42628
rect 15660 42508 15712 42560
rect 16948 42508 17000 42560
rect 17960 42508 18012 42560
rect 18788 42508 18840 42560
rect 21916 42712 21968 42764
rect 22100 42712 22152 42764
rect 23480 42755 23532 42764
rect 23480 42721 23489 42755
rect 23489 42721 23523 42755
rect 23523 42721 23532 42755
rect 23480 42712 23532 42721
rect 21548 42687 21600 42696
rect 21548 42653 21557 42687
rect 21557 42653 21591 42687
rect 21591 42653 21600 42687
rect 21548 42644 21600 42653
rect 21824 42644 21876 42696
rect 22008 42619 22060 42628
rect 22008 42585 22017 42619
rect 22017 42585 22051 42619
rect 22051 42585 22060 42619
rect 22008 42576 22060 42585
rect 22744 42619 22796 42628
rect 22744 42585 22753 42619
rect 22753 42585 22787 42619
rect 22787 42585 22796 42619
rect 22744 42576 22796 42585
rect 22836 42576 22888 42628
rect 26332 42780 26384 42832
rect 34612 42780 34664 42832
rect 24032 42712 24084 42764
rect 24492 42712 24544 42764
rect 23756 42644 23808 42696
rect 24676 42644 24728 42696
rect 25780 42712 25832 42764
rect 27068 42712 27120 42764
rect 32036 42712 32088 42764
rect 34428 42712 34480 42764
rect 34704 42755 34756 42764
rect 34704 42721 34713 42755
rect 34713 42721 34747 42755
rect 34747 42721 34756 42755
rect 34704 42712 34756 42721
rect 24860 42687 24912 42696
rect 24860 42653 24869 42687
rect 24869 42653 24903 42687
rect 24903 42653 24912 42687
rect 24860 42644 24912 42653
rect 25688 42687 25740 42696
rect 24032 42576 24084 42628
rect 25688 42653 25697 42687
rect 25697 42653 25731 42687
rect 25731 42653 25740 42687
rect 25688 42644 25740 42653
rect 29828 42687 29880 42696
rect 29828 42653 29837 42687
rect 29837 42653 29871 42687
rect 29871 42653 29880 42687
rect 29828 42644 29880 42653
rect 22192 42508 22244 42560
rect 22560 42551 22612 42560
rect 22560 42517 22569 42551
rect 22569 42517 22603 42551
rect 22603 42517 22612 42551
rect 22560 42508 22612 42517
rect 24584 42508 24636 42560
rect 24860 42508 24912 42560
rect 26056 42508 26108 42560
rect 26700 42551 26752 42560
rect 26700 42517 26709 42551
rect 26709 42517 26743 42551
rect 26743 42517 26752 42551
rect 26700 42508 26752 42517
rect 28632 42508 28684 42560
rect 28908 42508 28960 42560
rect 33784 42644 33836 42696
rect 33876 42644 33928 42696
rect 37280 42755 37332 42764
rect 37280 42721 37289 42755
rect 37289 42721 37323 42755
rect 37323 42721 37332 42755
rect 37280 42712 37332 42721
rect 38292 42755 38344 42764
rect 38292 42721 38301 42755
rect 38301 42721 38335 42755
rect 38335 42721 38344 42755
rect 38292 42712 38344 42721
rect 35164 42687 35216 42696
rect 35164 42653 35173 42687
rect 35173 42653 35207 42687
rect 35207 42653 35216 42687
rect 35164 42644 35216 42653
rect 35440 42687 35492 42696
rect 31392 42576 31444 42628
rect 31024 42508 31076 42560
rect 31760 42551 31812 42560
rect 31760 42517 31769 42551
rect 31769 42517 31803 42551
rect 31803 42517 31812 42551
rect 31760 42508 31812 42517
rect 34244 42576 34296 42628
rect 35440 42653 35449 42687
rect 35449 42653 35483 42687
rect 35483 42653 35492 42687
rect 35440 42644 35492 42653
rect 35992 42644 36044 42696
rect 36268 42687 36320 42696
rect 36268 42653 36277 42687
rect 36277 42653 36311 42687
rect 36311 42653 36320 42687
rect 36268 42644 36320 42653
rect 35348 42576 35400 42628
rect 37464 42644 37516 42696
rect 38016 42687 38068 42696
rect 38016 42653 38025 42687
rect 38025 42653 38059 42687
rect 38059 42653 38068 42687
rect 38016 42644 38068 42653
rect 48136 42687 48188 42696
rect 48136 42653 48145 42687
rect 48145 42653 48179 42687
rect 48179 42653 48188 42687
rect 48136 42644 48188 42653
rect 37188 42576 37240 42628
rect 35624 42508 35676 42560
rect 35900 42508 35952 42560
rect 36452 42508 36504 42560
rect 36544 42551 36596 42560
rect 36544 42517 36553 42551
rect 36553 42517 36587 42551
rect 36587 42517 36596 42551
rect 36544 42508 36596 42517
rect 37740 42508 37792 42560
rect 38568 42508 38620 42560
rect 40040 42508 40092 42560
rect 47952 42551 48004 42560
rect 47952 42517 47961 42551
rect 47961 42517 47995 42551
rect 47995 42517 48004 42551
rect 47952 42508 48004 42517
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 11060 42304 11112 42356
rect 12072 42304 12124 42356
rect 12440 42304 12492 42356
rect 13452 42304 13504 42356
rect 14096 42347 14148 42356
rect 14096 42313 14105 42347
rect 14105 42313 14139 42347
rect 14139 42313 14148 42347
rect 14096 42304 14148 42313
rect 15200 42347 15252 42356
rect 15200 42313 15209 42347
rect 15209 42313 15243 42347
rect 15243 42313 15252 42347
rect 15200 42304 15252 42313
rect 20536 42347 20588 42356
rect 18144 42236 18196 42288
rect 19984 42236 20036 42288
rect 20536 42313 20545 42347
rect 20545 42313 20579 42347
rect 20579 42313 20588 42347
rect 20536 42304 20588 42313
rect 21180 42347 21232 42356
rect 21180 42313 21189 42347
rect 21189 42313 21223 42347
rect 21223 42313 21232 42347
rect 21180 42304 21232 42313
rect 21824 42347 21876 42356
rect 21824 42313 21833 42347
rect 21833 42313 21867 42347
rect 21867 42313 21876 42347
rect 21824 42304 21876 42313
rect 24032 42347 24084 42356
rect 24032 42313 24041 42347
rect 24041 42313 24075 42347
rect 24075 42313 24084 42347
rect 24032 42304 24084 42313
rect 24860 42347 24912 42356
rect 24860 42313 24869 42347
rect 24869 42313 24903 42347
rect 24903 42313 24912 42347
rect 24860 42304 24912 42313
rect 20996 42236 21048 42288
rect 21732 42236 21784 42288
rect 12256 42168 12308 42220
rect 12992 42211 13044 42220
rect 12992 42177 13001 42211
rect 13001 42177 13035 42211
rect 13035 42177 13044 42211
rect 12992 42168 13044 42177
rect 15660 42211 15712 42220
rect 15660 42177 15669 42211
rect 15669 42177 15703 42211
rect 15703 42177 15712 42211
rect 15660 42168 15712 42177
rect 16672 42211 16724 42220
rect 16672 42177 16681 42211
rect 16681 42177 16715 42211
rect 16715 42177 16724 42211
rect 16672 42168 16724 42177
rect 17132 42168 17184 42220
rect 17960 42211 18012 42220
rect 17960 42177 17969 42211
rect 17969 42177 18003 42211
rect 18003 42177 18012 42211
rect 17960 42168 18012 42177
rect 19340 42168 19392 42220
rect 20904 42168 20956 42220
rect 21180 42168 21232 42220
rect 21456 42168 21508 42220
rect 21548 42168 21600 42220
rect 22008 42211 22060 42220
rect 22008 42177 22017 42211
rect 22017 42177 22051 42211
rect 22051 42177 22060 42211
rect 22008 42168 22060 42177
rect 22284 42211 22336 42220
rect 22284 42177 22293 42211
rect 22293 42177 22327 42211
rect 22327 42177 22336 42211
rect 22284 42168 22336 42177
rect 22468 42211 22520 42220
rect 22468 42177 22477 42211
rect 22477 42177 22511 42211
rect 22511 42177 22520 42211
rect 22468 42168 22520 42177
rect 22560 42168 22612 42220
rect 23296 42236 23348 42288
rect 30472 42304 30524 42356
rect 30656 42304 30708 42356
rect 31760 42304 31812 42356
rect 35348 42347 35400 42356
rect 35348 42313 35357 42347
rect 35357 42313 35391 42347
rect 35391 42313 35400 42347
rect 35348 42304 35400 42313
rect 35532 42304 35584 42356
rect 35992 42347 36044 42356
rect 35992 42313 36001 42347
rect 36001 42313 36035 42347
rect 36035 42313 36044 42347
rect 35992 42304 36044 42313
rect 31852 42236 31904 42288
rect 34152 42236 34204 42288
rect 15936 42143 15988 42152
rect 15936 42109 15945 42143
rect 15945 42109 15979 42143
rect 15979 42109 15988 42143
rect 15936 42100 15988 42109
rect 16764 42100 16816 42152
rect 18328 42100 18380 42152
rect 18420 42100 18472 42152
rect 21916 42100 21968 42152
rect 24400 42168 24452 42220
rect 24584 42211 24636 42220
rect 24584 42177 24593 42211
rect 24593 42177 24627 42211
rect 24627 42177 24636 42211
rect 25504 42211 25556 42220
rect 24584 42168 24636 42177
rect 25504 42177 25513 42211
rect 25513 42177 25547 42211
rect 25547 42177 25556 42211
rect 25504 42168 25556 42177
rect 18788 42032 18840 42084
rect 19340 42032 19392 42084
rect 19984 42075 20036 42084
rect 19984 42041 19993 42075
rect 19993 42041 20027 42075
rect 20027 42041 20036 42075
rect 19984 42032 20036 42041
rect 10784 41964 10836 42016
rect 15752 42007 15804 42016
rect 15752 41973 15761 42007
rect 15761 41973 15795 42007
rect 15795 41973 15804 42007
rect 15752 41964 15804 41973
rect 16856 41964 16908 42016
rect 20720 41964 20772 42016
rect 21640 41964 21692 42016
rect 21916 41964 21968 42016
rect 29092 42168 29144 42220
rect 30656 42168 30708 42220
rect 35348 42168 35400 42220
rect 37464 42211 37516 42220
rect 29276 42143 29328 42152
rect 25964 41964 26016 42016
rect 27160 42007 27212 42016
rect 27160 41973 27169 42007
rect 27169 41973 27203 42007
rect 27203 41973 27212 42007
rect 27160 41964 27212 41973
rect 29276 42109 29285 42143
rect 29285 42109 29319 42143
rect 29319 42109 29328 42143
rect 29276 42100 29328 42109
rect 30748 42100 30800 42152
rect 30932 42100 30984 42152
rect 31852 42100 31904 42152
rect 32128 42143 32180 42152
rect 32128 42109 32137 42143
rect 32137 42109 32171 42143
rect 32171 42109 32180 42143
rect 32128 42100 32180 42109
rect 33600 42100 33652 42152
rect 35440 42100 35492 42152
rect 37464 42177 37473 42211
rect 37473 42177 37507 42211
rect 37507 42177 37516 42211
rect 37464 42168 37516 42177
rect 38292 42211 38344 42220
rect 36360 42143 36412 42152
rect 36360 42109 36369 42143
rect 36369 42109 36403 42143
rect 36403 42109 36412 42143
rect 36360 42100 36412 42109
rect 37280 42100 37332 42152
rect 38292 42177 38301 42211
rect 38301 42177 38335 42211
rect 38335 42177 38344 42211
rect 38292 42168 38344 42177
rect 38476 42211 38528 42220
rect 38476 42177 38485 42211
rect 38485 42177 38519 42211
rect 38519 42177 38528 42211
rect 38476 42168 38528 42177
rect 38568 42211 38620 42220
rect 38568 42177 38577 42211
rect 38577 42177 38611 42211
rect 38611 42177 38620 42211
rect 38568 42168 38620 42177
rect 32036 42032 32088 42084
rect 33876 42032 33928 42084
rect 37188 42032 37240 42084
rect 37648 42075 37700 42084
rect 37648 42041 37657 42075
rect 37657 42041 37691 42075
rect 37691 42041 37700 42075
rect 39120 42100 39172 42152
rect 37648 42032 37700 42041
rect 30380 42007 30432 42016
rect 30380 41973 30389 42007
rect 30389 41973 30423 42007
rect 30423 41973 30432 42007
rect 30380 41964 30432 41973
rect 33140 41964 33192 42016
rect 35164 41964 35216 42016
rect 35808 41964 35860 42016
rect 37924 41964 37976 42016
rect 39304 41964 39356 42016
rect 40040 41964 40092 42016
rect 40224 42007 40276 42016
rect 40224 41973 40233 42007
rect 40233 41973 40267 42007
rect 40267 41973 40276 42007
rect 40224 41964 40276 41973
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 13544 41760 13596 41812
rect 14188 41803 14240 41812
rect 14188 41769 14197 41803
rect 14197 41769 14231 41803
rect 14231 41769 14240 41803
rect 14188 41760 14240 41769
rect 15568 41803 15620 41812
rect 15568 41769 15577 41803
rect 15577 41769 15611 41803
rect 15611 41769 15620 41803
rect 15568 41760 15620 41769
rect 15752 41760 15804 41812
rect 17684 41760 17736 41812
rect 18420 41803 18472 41812
rect 18420 41769 18429 41803
rect 18429 41769 18463 41803
rect 18463 41769 18472 41803
rect 18420 41760 18472 41769
rect 19432 41760 19484 41812
rect 20720 41803 20772 41812
rect 20720 41769 20729 41803
rect 20729 41769 20763 41803
rect 20763 41769 20772 41803
rect 20720 41760 20772 41769
rect 22284 41760 22336 41812
rect 25964 41760 26016 41812
rect 27068 41760 27120 41812
rect 27712 41760 27764 41812
rect 28080 41760 28132 41812
rect 14740 41599 14792 41608
rect 14740 41565 14752 41599
rect 14752 41565 14786 41599
rect 14786 41565 14792 41599
rect 14740 41556 14792 41565
rect 11060 41488 11112 41540
rect 12164 41488 12216 41540
rect 15660 41556 15712 41608
rect 15936 41556 15988 41608
rect 16764 41599 16816 41608
rect 16764 41565 16773 41599
rect 16773 41565 16807 41599
rect 16807 41565 16816 41599
rect 16764 41556 16816 41565
rect 16948 41599 17000 41608
rect 16948 41565 16957 41599
rect 16957 41565 16991 41599
rect 16991 41565 17000 41599
rect 16948 41556 17000 41565
rect 18788 41624 18840 41676
rect 19156 41624 19208 41676
rect 20536 41624 20588 41676
rect 21364 41624 21416 41676
rect 18512 41599 18564 41608
rect 16120 41488 16172 41540
rect 18512 41565 18521 41599
rect 18521 41565 18555 41599
rect 18555 41565 18564 41599
rect 18512 41556 18564 41565
rect 19432 41599 19484 41608
rect 19432 41565 19441 41599
rect 19441 41565 19475 41599
rect 19475 41565 19484 41599
rect 19432 41556 19484 41565
rect 20352 41556 20404 41608
rect 21732 41556 21784 41608
rect 17224 41488 17276 41540
rect 18420 41488 18472 41540
rect 9588 41420 9640 41472
rect 13544 41420 13596 41472
rect 15108 41420 15160 41472
rect 16764 41420 16816 41472
rect 17960 41420 18012 41472
rect 21088 41420 21140 41472
rect 23112 41692 23164 41744
rect 24492 41667 24544 41676
rect 24492 41633 24501 41667
rect 24501 41633 24535 41667
rect 24535 41633 24544 41667
rect 24492 41624 24544 41633
rect 25412 41692 25464 41744
rect 27344 41692 27396 41744
rect 34244 41760 34296 41812
rect 35348 41760 35400 41812
rect 36360 41803 36412 41812
rect 36360 41769 36369 41803
rect 36369 41769 36403 41803
rect 36403 41769 36412 41803
rect 36360 41760 36412 41769
rect 38292 41803 38344 41812
rect 38292 41769 38301 41803
rect 38301 41769 38335 41803
rect 38335 41769 38344 41803
rect 38292 41760 38344 41769
rect 34520 41692 34572 41744
rect 34888 41692 34940 41744
rect 36176 41692 36228 41744
rect 40040 41760 40092 41812
rect 29092 41624 29144 41676
rect 31208 41667 31260 41676
rect 31208 41633 31217 41667
rect 31217 41633 31251 41667
rect 31251 41633 31260 41667
rect 31208 41624 31260 41633
rect 22560 41556 22612 41608
rect 23940 41556 23992 41608
rect 24676 41556 24728 41608
rect 29000 41556 29052 41608
rect 29920 41556 29972 41608
rect 30196 41556 30248 41608
rect 33692 41624 33744 41676
rect 36544 41624 36596 41676
rect 32404 41599 32456 41608
rect 32404 41565 32413 41599
rect 32413 41565 32447 41599
rect 32447 41565 32456 41599
rect 32404 41556 32456 41565
rect 33416 41556 33468 41608
rect 33600 41599 33652 41608
rect 33600 41565 33609 41599
rect 33609 41565 33643 41599
rect 33643 41565 33652 41599
rect 33600 41556 33652 41565
rect 33876 41556 33928 41608
rect 35716 41556 35768 41608
rect 38568 41692 38620 41744
rect 40224 41692 40276 41744
rect 37740 41667 37792 41676
rect 37740 41633 37749 41667
rect 37749 41633 37783 41667
rect 37783 41633 37792 41667
rect 37740 41624 37792 41633
rect 37648 41599 37700 41608
rect 23112 41420 23164 41472
rect 23480 41420 23532 41472
rect 24216 41420 24268 41472
rect 25320 41420 25372 41472
rect 25780 41420 25832 41472
rect 27712 41420 27764 41472
rect 28908 41463 28960 41472
rect 28908 41429 28917 41463
rect 28917 41429 28951 41463
rect 28951 41429 28960 41463
rect 28908 41420 28960 41429
rect 30472 41420 30524 41472
rect 32496 41420 32548 41472
rect 33324 41463 33376 41472
rect 33324 41429 33333 41463
rect 33333 41429 33367 41463
rect 33367 41429 33376 41463
rect 33324 41420 33376 41429
rect 33784 41463 33836 41472
rect 33784 41429 33793 41463
rect 33793 41429 33827 41463
rect 33827 41429 33836 41463
rect 34336 41488 34388 41540
rect 33784 41420 33836 41429
rect 34612 41420 34664 41472
rect 37648 41565 37657 41599
rect 37657 41565 37691 41599
rect 37691 41565 37700 41599
rect 37648 41556 37700 41565
rect 38752 41556 38804 41608
rect 39304 41599 39356 41608
rect 39304 41565 39313 41599
rect 39313 41565 39347 41599
rect 39347 41565 39356 41599
rect 39304 41556 39356 41565
rect 37004 41420 37056 41472
rect 38016 41420 38068 41472
rect 38292 41420 38344 41472
rect 40500 41463 40552 41472
rect 40500 41429 40509 41463
rect 40509 41429 40543 41463
rect 40543 41429 40552 41463
rect 40500 41420 40552 41429
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 13544 41216 13596 41268
rect 13820 41216 13872 41268
rect 14740 41216 14792 41268
rect 15108 41259 15160 41268
rect 15108 41225 15117 41259
rect 15117 41225 15151 41259
rect 15151 41225 15160 41259
rect 16120 41259 16172 41268
rect 15108 41216 15160 41225
rect 11060 41080 11112 41132
rect 15660 41148 15712 41200
rect 15200 41080 15252 41132
rect 16120 41225 16129 41259
rect 16129 41225 16163 41259
rect 16163 41225 16172 41259
rect 16120 41216 16172 41225
rect 16948 41216 17000 41268
rect 18144 41216 18196 41268
rect 17592 41148 17644 41200
rect 15936 41123 15988 41132
rect 15936 41089 15945 41123
rect 15945 41089 15979 41123
rect 15979 41089 15988 41123
rect 16856 41123 16908 41132
rect 15936 41080 15988 41089
rect 16856 41089 16865 41123
rect 16865 41089 16899 41123
rect 16899 41089 16908 41123
rect 16856 41080 16908 41089
rect 15660 41055 15712 41064
rect 15660 41021 15669 41055
rect 15669 41021 15703 41055
rect 15703 41021 15712 41055
rect 15660 41012 15712 41021
rect 16764 41055 16816 41064
rect 16764 41021 16773 41055
rect 16773 41021 16807 41055
rect 16807 41021 16816 41055
rect 16764 41012 16816 41021
rect 18144 41080 18196 41132
rect 18420 41123 18472 41132
rect 18420 41089 18429 41123
rect 18429 41089 18463 41123
rect 18463 41089 18472 41123
rect 18420 41080 18472 41089
rect 18880 41148 18932 41200
rect 19708 41216 19760 41268
rect 20076 41216 20128 41268
rect 20352 41259 20404 41268
rect 20352 41225 20361 41259
rect 20361 41225 20395 41259
rect 20395 41225 20404 41259
rect 20352 41216 20404 41225
rect 22008 41216 22060 41268
rect 23020 41216 23072 41268
rect 24308 41216 24360 41268
rect 27436 41216 27488 41268
rect 27804 41259 27856 41268
rect 27804 41225 27813 41259
rect 27813 41225 27847 41259
rect 27847 41225 27856 41259
rect 27804 41216 27856 41225
rect 29092 41259 29144 41268
rect 29092 41225 29101 41259
rect 29101 41225 29135 41259
rect 29135 41225 29144 41259
rect 29092 41216 29144 41225
rect 33784 41216 33836 41268
rect 36544 41259 36596 41268
rect 36544 41225 36553 41259
rect 36553 41225 36587 41259
rect 36587 41225 36596 41259
rect 36544 41216 36596 41225
rect 38752 41216 38804 41268
rect 40224 41216 40276 41268
rect 19064 41080 19116 41132
rect 11060 40876 11112 40928
rect 12716 40876 12768 40928
rect 13544 40876 13596 40928
rect 18328 41012 18380 41064
rect 19248 41123 19300 41132
rect 19248 41089 19258 41123
rect 19258 41089 19292 41123
rect 19292 41089 19300 41123
rect 19984 41148 20036 41200
rect 19248 41080 19300 41089
rect 19616 41123 19668 41132
rect 19616 41089 19649 41123
rect 19649 41089 19668 41123
rect 19616 41080 19668 41089
rect 18512 40944 18564 40996
rect 19432 41012 19484 41064
rect 23480 41148 23532 41200
rect 25964 41148 26016 41200
rect 29000 41148 29052 41200
rect 30840 41148 30892 41200
rect 34152 41148 34204 41200
rect 36268 41148 36320 41200
rect 38476 41191 38528 41200
rect 38476 41157 38485 41191
rect 38485 41157 38519 41191
rect 38519 41157 38528 41191
rect 38476 41148 38528 41157
rect 20444 41123 20496 41132
rect 20076 40944 20128 40996
rect 20444 41089 20453 41123
rect 20453 41089 20487 41123
rect 20487 41089 20496 41123
rect 20444 41080 20496 41089
rect 21824 41123 21876 41132
rect 21824 41089 21833 41123
rect 21833 41089 21867 41123
rect 21867 41089 21876 41123
rect 21824 41080 21876 41089
rect 21272 41012 21324 41064
rect 21732 41012 21784 41064
rect 22744 41080 22796 41132
rect 24400 41123 24452 41132
rect 24400 41089 24409 41123
rect 24409 41089 24443 41123
rect 24443 41089 24452 41123
rect 24400 41080 24452 41089
rect 24492 41123 24544 41132
rect 24492 41089 24501 41123
rect 24501 41089 24535 41123
rect 24535 41089 24544 41123
rect 24492 41080 24544 41089
rect 24952 41080 25004 41132
rect 25228 41080 25280 41132
rect 25780 41080 25832 41132
rect 29092 41080 29144 41132
rect 32128 41123 32180 41132
rect 32128 41089 32137 41123
rect 32137 41089 32171 41123
rect 32171 41089 32180 41123
rect 32128 41080 32180 41089
rect 32680 41080 32732 41132
rect 34704 41080 34756 41132
rect 23848 41012 23900 41064
rect 25504 41012 25556 41064
rect 34520 41012 34572 41064
rect 34888 41012 34940 41064
rect 24032 40944 24084 40996
rect 24676 40987 24728 40996
rect 24676 40953 24685 40987
rect 24685 40953 24719 40987
rect 24719 40953 24728 40987
rect 24676 40944 24728 40953
rect 25412 40944 25464 40996
rect 29000 40944 29052 40996
rect 35808 41080 35860 41132
rect 37740 41080 37792 41132
rect 37832 41080 37884 41132
rect 38568 41080 38620 41132
rect 35900 41012 35952 41064
rect 36084 41012 36136 41064
rect 36176 41012 36228 41064
rect 19156 40876 19208 40928
rect 19248 40876 19300 40928
rect 24584 40876 24636 40928
rect 24768 40876 24820 40928
rect 27068 40876 27120 40928
rect 30564 40876 30616 40928
rect 31300 40876 31352 40928
rect 35348 40944 35400 40996
rect 37832 40944 37884 40996
rect 40040 40944 40092 40996
rect 33232 40876 33284 40928
rect 33508 40919 33560 40928
rect 33508 40885 33517 40919
rect 33517 40885 33551 40919
rect 33551 40885 33560 40919
rect 33508 40876 33560 40885
rect 34152 40919 34204 40928
rect 34152 40885 34161 40919
rect 34161 40885 34195 40919
rect 34195 40885 34204 40919
rect 34152 40876 34204 40885
rect 34796 40876 34848 40928
rect 35808 40919 35860 40928
rect 35808 40885 35817 40919
rect 35817 40885 35851 40919
rect 35851 40885 35860 40919
rect 35808 40876 35860 40885
rect 35900 40919 35952 40928
rect 35900 40885 35909 40919
rect 35909 40885 35943 40919
rect 35943 40885 35952 40919
rect 37280 40919 37332 40928
rect 35900 40876 35952 40885
rect 37280 40885 37289 40919
rect 37289 40885 37323 40919
rect 37323 40885 37332 40919
rect 37280 40876 37332 40885
rect 39672 40919 39724 40928
rect 39672 40885 39681 40919
rect 39681 40885 39715 40919
rect 39715 40885 39724 40919
rect 39672 40876 39724 40885
rect 43168 40876 43220 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 12716 40672 12768 40724
rect 12900 40715 12952 40724
rect 12900 40681 12909 40715
rect 12909 40681 12943 40715
rect 12943 40681 12952 40715
rect 12900 40672 12952 40681
rect 12072 40604 12124 40656
rect 13820 40672 13872 40724
rect 15568 40672 15620 40724
rect 17868 40672 17920 40724
rect 18696 40715 18748 40724
rect 18696 40681 18705 40715
rect 18705 40681 18739 40715
rect 18739 40681 18748 40715
rect 18696 40672 18748 40681
rect 18788 40672 18840 40724
rect 19432 40672 19484 40724
rect 20076 40672 20128 40724
rect 15200 40647 15252 40656
rect 15200 40613 15209 40647
rect 15209 40613 15243 40647
rect 15243 40613 15252 40647
rect 15200 40604 15252 40613
rect 17592 40604 17644 40656
rect 18420 40604 18472 40656
rect 19524 40604 19576 40656
rect 24768 40672 24820 40724
rect 12716 40536 12768 40588
rect 15016 40511 15068 40520
rect 15016 40477 15025 40511
rect 15025 40477 15059 40511
rect 15059 40477 15068 40511
rect 15016 40468 15068 40477
rect 15108 40468 15160 40520
rect 16580 40468 16632 40520
rect 17868 40468 17920 40520
rect 18328 40536 18380 40588
rect 19064 40536 19116 40588
rect 18144 40511 18196 40520
rect 18144 40477 18154 40511
rect 18154 40477 18188 40511
rect 18188 40477 18196 40511
rect 18144 40468 18196 40477
rect 18512 40511 18564 40520
rect 18512 40477 18526 40511
rect 18526 40477 18560 40511
rect 18560 40477 18564 40511
rect 18512 40468 18564 40477
rect 18880 40468 18932 40520
rect 19800 40536 19852 40588
rect 20076 40536 20128 40588
rect 23848 40647 23900 40656
rect 23848 40613 23857 40647
rect 23857 40613 23891 40647
rect 23891 40613 23900 40647
rect 23848 40604 23900 40613
rect 22744 40579 22796 40588
rect 22744 40545 22753 40579
rect 22753 40545 22787 40579
rect 22787 40545 22796 40579
rect 22744 40536 22796 40545
rect 24952 40672 25004 40724
rect 25688 40672 25740 40724
rect 25964 40715 26016 40724
rect 25964 40681 25973 40715
rect 25973 40681 26007 40715
rect 26007 40681 26016 40715
rect 25964 40672 26016 40681
rect 27068 40672 27120 40724
rect 32496 40672 32548 40724
rect 32680 40672 32732 40724
rect 34152 40715 34204 40724
rect 34152 40681 34161 40715
rect 34161 40681 34195 40715
rect 34195 40681 34204 40715
rect 34152 40672 34204 40681
rect 35992 40672 36044 40724
rect 37096 40672 37148 40724
rect 37740 40715 37792 40724
rect 37740 40681 37749 40715
rect 37749 40681 37783 40715
rect 37783 40681 37792 40715
rect 37740 40672 37792 40681
rect 40224 40672 40276 40724
rect 25872 40604 25924 40656
rect 32312 40604 32364 40656
rect 33876 40604 33928 40656
rect 34428 40604 34480 40656
rect 36176 40604 36228 40656
rect 41052 40604 41104 40656
rect 20536 40468 20588 40520
rect 21088 40511 21140 40520
rect 21088 40477 21097 40511
rect 21097 40477 21131 40511
rect 21131 40477 21140 40511
rect 21088 40468 21140 40477
rect 21272 40511 21324 40520
rect 21272 40477 21281 40511
rect 21281 40477 21315 40511
rect 21315 40477 21324 40511
rect 21272 40468 21324 40477
rect 21916 40511 21968 40520
rect 21916 40477 21925 40511
rect 21925 40477 21959 40511
rect 21959 40477 21968 40511
rect 21916 40468 21968 40477
rect 1584 40400 1636 40452
rect 2044 40443 2096 40452
rect 2044 40409 2053 40443
rect 2053 40409 2087 40443
rect 2087 40409 2096 40443
rect 2044 40400 2096 40409
rect 18328 40443 18380 40452
rect 18328 40409 18337 40443
rect 18337 40409 18371 40443
rect 18371 40409 18380 40443
rect 18328 40400 18380 40409
rect 18788 40400 18840 40452
rect 14004 40332 14056 40384
rect 15292 40332 15344 40384
rect 17040 40375 17092 40384
rect 17040 40341 17049 40375
rect 17049 40341 17083 40375
rect 17083 40341 17092 40375
rect 17040 40332 17092 40341
rect 19064 40332 19116 40384
rect 22192 40400 22244 40452
rect 23020 40511 23072 40520
rect 23020 40477 23029 40511
rect 23029 40477 23063 40511
rect 23063 40477 23072 40511
rect 23020 40468 23072 40477
rect 23756 40468 23808 40520
rect 26332 40536 26384 40588
rect 24216 40468 24268 40520
rect 24584 40511 24636 40520
rect 24584 40477 24594 40511
rect 24594 40477 24628 40511
rect 24628 40477 24636 40511
rect 24584 40468 24636 40477
rect 25044 40468 25096 40520
rect 27160 40536 27212 40588
rect 29092 40536 29144 40588
rect 24768 40443 24820 40452
rect 24768 40409 24777 40443
rect 24777 40409 24811 40443
rect 24811 40409 24820 40443
rect 24768 40400 24820 40409
rect 24860 40443 24912 40452
rect 24860 40409 24869 40443
rect 24869 40409 24903 40443
rect 24903 40409 24912 40443
rect 25596 40443 25648 40452
rect 24860 40400 24912 40409
rect 25596 40409 25605 40443
rect 25605 40409 25639 40443
rect 25639 40409 25648 40443
rect 25596 40400 25648 40409
rect 19524 40332 19576 40384
rect 19800 40332 19852 40384
rect 23664 40375 23716 40384
rect 23664 40341 23673 40375
rect 23673 40341 23707 40375
rect 23707 40341 23716 40375
rect 23664 40332 23716 40341
rect 24032 40332 24084 40384
rect 33324 40536 33376 40588
rect 33600 40536 33652 40588
rect 34336 40536 34388 40588
rect 35808 40536 35860 40588
rect 36636 40536 36688 40588
rect 31760 40511 31812 40520
rect 31760 40477 31769 40511
rect 31769 40477 31803 40511
rect 31803 40477 31812 40511
rect 33232 40511 33284 40520
rect 31760 40468 31812 40477
rect 33232 40477 33241 40511
rect 33241 40477 33275 40511
rect 33275 40477 33284 40511
rect 33232 40468 33284 40477
rect 34704 40511 34756 40520
rect 26240 40400 26292 40452
rect 27620 40400 27672 40452
rect 32404 40443 32456 40452
rect 32404 40409 32429 40443
rect 32429 40409 32456 40443
rect 32404 40400 32456 40409
rect 34704 40477 34713 40511
rect 34713 40477 34747 40511
rect 34747 40477 34756 40511
rect 34704 40468 34756 40477
rect 34152 40443 34204 40452
rect 34152 40409 34161 40443
rect 34161 40409 34195 40443
rect 34195 40409 34204 40443
rect 34152 40400 34204 40409
rect 35348 40468 35400 40520
rect 35532 40511 35584 40520
rect 35532 40477 35541 40511
rect 35541 40477 35575 40511
rect 35575 40477 35584 40511
rect 35532 40468 35584 40477
rect 35900 40468 35952 40520
rect 37924 40511 37976 40520
rect 32312 40332 32364 40384
rect 34704 40332 34756 40384
rect 36176 40400 36228 40452
rect 35348 40332 35400 40384
rect 35440 40332 35492 40384
rect 37924 40477 37933 40511
rect 37933 40477 37967 40511
rect 37967 40477 37976 40511
rect 37924 40468 37976 40477
rect 36912 40443 36964 40452
rect 36912 40409 36921 40443
rect 36921 40409 36955 40443
rect 36955 40409 36964 40443
rect 36912 40400 36964 40409
rect 37096 40443 37148 40452
rect 37096 40409 37105 40443
rect 37105 40409 37139 40443
rect 37139 40409 37148 40443
rect 37096 40400 37148 40409
rect 37464 40332 37516 40384
rect 38660 40332 38712 40384
rect 39672 40332 39724 40384
rect 41052 40375 41104 40384
rect 41052 40341 41061 40375
rect 41061 40341 41095 40375
rect 41095 40341 41104 40375
rect 41052 40332 41104 40341
rect 41604 40400 41656 40452
rect 47308 40443 47360 40452
rect 47308 40409 47317 40443
rect 47317 40409 47351 40443
rect 47351 40409 47360 40443
rect 47308 40400 47360 40409
rect 41512 40375 41564 40384
rect 41512 40341 41521 40375
rect 41521 40341 41555 40375
rect 41555 40341 41564 40375
rect 41512 40332 41564 40341
rect 42064 40375 42116 40384
rect 42064 40341 42073 40375
rect 42073 40341 42107 40375
rect 42107 40341 42116 40375
rect 42064 40332 42116 40341
rect 48044 40375 48096 40384
rect 48044 40341 48053 40375
rect 48053 40341 48087 40375
rect 48087 40341 48096 40375
rect 48044 40332 48096 40341
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 1584 40171 1636 40180
rect 1584 40137 1593 40171
rect 1593 40137 1627 40171
rect 1627 40137 1636 40171
rect 1584 40128 1636 40137
rect 13912 40128 13964 40180
rect 14832 40128 14884 40180
rect 15476 40171 15528 40180
rect 15476 40137 15485 40171
rect 15485 40137 15519 40171
rect 15519 40137 15528 40171
rect 15476 40128 15528 40137
rect 17040 40128 17092 40180
rect 20260 40128 20312 40180
rect 23204 40128 23256 40180
rect 23664 40128 23716 40180
rect 24768 40128 24820 40180
rect 25504 40171 25556 40180
rect 25504 40137 25513 40171
rect 25513 40137 25547 40171
rect 25547 40137 25556 40171
rect 25504 40128 25556 40137
rect 26148 40128 26200 40180
rect 27252 40128 27304 40180
rect 35532 40171 35584 40180
rect 35532 40137 35541 40171
rect 35541 40137 35575 40171
rect 35575 40137 35584 40171
rect 35532 40128 35584 40137
rect 35992 40128 36044 40180
rect 36912 40128 36964 40180
rect 11796 40060 11848 40112
rect 12716 40060 12768 40112
rect 17224 40060 17276 40112
rect 12072 40035 12124 40044
rect 12072 40001 12081 40035
rect 12081 40001 12115 40035
rect 12115 40001 12124 40035
rect 12072 39992 12124 40001
rect 12440 39992 12492 40044
rect 14648 39992 14700 40044
rect 17592 40060 17644 40112
rect 19156 40103 19208 40112
rect 19156 40069 19165 40103
rect 19165 40069 19199 40103
rect 19199 40069 19208 40103
rect 19156 40060 19208 40069
rect 19340 40103 19392 40112
rect 19340 40069 19349 40103
rect 19349 40069 19383 40103
rect 19383 40069 19392 40103
rect 19340 40060 19392 40069
rect 20076 40060 20128 40112
rect 20536 40103 20588 40112
rect 20536 40069 20545 40103
rect 20545 40069 20579 40103
rect 20579 40069 20588 40103
rect 20536 40060 20588 40069
rect 23940 40060 23992 40112
rect 14280 39924 14332 39976
rect 17040 39924 17092 39976
rect 17132 39924 17184 39976
rect 17408 39924 17460 39976
rect 18880 39924 18932 39976
rect 19984 39924 20036 39976
rect 20352 40035 20404 40044
rect 20352 40001 20361 40035
rect 20361 40001 20395 40035
rect 20395 40001 20404 40035
rect 20352 39992 20404 40001
rect 21180 40035 21232 40044
rect 20628 39924 20680 39976
rect 14188 39856 14240 39908
rect 15016 39856 15068 39908
rect 18328 39856 18380 39908
rect 21180 40001 21189 40035
rect 21189 40001 21223 40035
rect 21223 40001 21232 40035
rect 21180 39992 21232 40001
rect 22008 40035 22060 40044
rect 22008 40001 22024 40035
rect 22024 40001 22060 40035
rect 22008 39992 22060 40001
rect 23020 40035 23072 40044
rect 23020 40001 23029 40035
rect 23029 40001 23063 40035
rect 23063 40001 23072 40035
rect 23020 39992 23072 40001
rect 23572 39992 23624 40044
rect 25596 40060 25648 40112
rect 25780 40060 25832 40112
rect 25504 39992 25556 40044
rect 25964 40060 26016 40112
rect 26240 40060 26292 40112
rect 27068 40035 27120 40044
rect 27068 40001 27077 40035
rect 27077 40001 27111 40035
rect 27111 40001 27120 40035
rect 27068 39992 27120 40001
rect 22192 39924 22244 39976
rect 24032 39967 24084 39976
rect 24032 39933 24041 39967
rect 24041 39933 24075 39967
rect 24075 39933 24084 39967
rect 24032 39924 24084 39933
rect 25044 39856 25096 39908
rect 15660 39788 15712 39840
rect 16304 39788 16356 39840
rect 17224 39788 17276 39840
rect 18052 39788 18104 39840
rect 18420 39831 18472 39840
rect 18420 39797 18429 39831
rect 18429 39797 18463 39831
rect 18463 39797 18472 39831
rect 18420 39788 18472 39797
rect 19432 39788 19484 39840
rect 20444 39788 20496 39840
rect 20812 39788 20864 39840
rect 21824 39788 21876 39840
rect 22284 39788 22336 39840
rect 24676 39788 24728 39840
rect 26700 39924 26752 39976
rect 27160 39924 27212 39976
rect 27528 39992 27580 40044
rect 32128 40060 32180 40112
rect 33968 40060 34020 40112
rect 30104 40035 30156 40044
rect 30104 40001 30113 40035
rect 30113 40001 30147 40035
rect 30147 40001 30156 40035
rect 30104 39992 30156 40001
rect 30288 40035 30340 40044
rect 30288 40001 30297 40035
rect 30297 40001 30331 40035
rect 30331 40001 30340 40035
rect 30288 39992 30340 40001
rect 30380 39992 30432 40044
rect 30472 39992 30524 40044
rect 32312 39992 32364 40044
rect 33232 39992 33284 40044
rect 33600 40035 33652 40044
rect 33600 40001 33609 40035
rect 33609 40001 33643 40035
rect 33643 40001 33652 40035
rect 33600 39992 33652 40001
rect 33784 39992 33836 40044
rect 34336 39992 34388 40044
rect 30196 39924 30248 39976
rect 32036 39924 32088 39976
rect 26056 39856 26108 39908
rect 29368 39899 29420 39908
rect 25872 39831 25924 39840
rect 25872 39797 25881 39831
rect 25881 39797 25915 39831
rect 25915 39797 25924 39831
rect 25872 39788 25924 39797
rect 26700 39788 26752 39840
rect 28356 39831 28408 39840
rect 28356 39797 28365 39831
rect 28365 39797 28399 39831
rect 28399 39797 28408 39831
rect 28356 39788 28408 39797
rect 29368 39865 29377 39899
rect 29377 39865 29411 39899
rect 29411 39865 29420 39899
rect 29368 39856 29420 39865
rect 30472 39856 30524 39908
rect 33416 39899 33468 39908
rect 33416 39865 33425 39899
rect 33425 39865 33459 39899
rect 33459 39865 33468 39899
rect 33416 39856 33468 39865
rect 34520 39967 34572 39976
rect 34520 39933 34529 39967
rect 34529 39933 34563 39967
rect 34563 39933 34572 39967
rect 35440 40060 35492 40112
rect 35900 39992 35952 40044
rect 34520 39924 34572 39933
rect 35440 39924 35492 39976
rect 35808 39967 35860 39976
rect 35808 39933 35817 39967
rect 35817 39933 35851 39967
rect 35851 39933 35860 39967
rect 35808 39924 35860 39933
rect 36360 39992 36412 40044
rect 36544 40035 36596 40044
rect 36544 40001 36553 40035
rect 36553 40001 36587 40035
rect 36587 40001 36596 40035
rect 36544 39992 36596 40001
rect 37464 40035 37516 40044
rect 37464 40001 37473 40035
rect 37473 40001 37507 40035
rect 37507 40001 37516 40035
rect 37464 39992 37516 40001
rect 41604 40171 41656 40180
rect 41604 40137 41613 40171
rect 41613 40137 41647 40171
rect 41647 40137 41656 40171
rect 41604 40128 41656 40137
rect 38844 40035 38896 40044
rect 36636 39924 36688 39976
rect 37372 39924 37424 39976
rect 37924 39924 37976 39976
rect 38016 39924 38068 39976
rect 38844 40001 38853 40035
rect 38853 40001 38887 40035
rect 38887 40001 38896 40035
rect 38844 39992 38896 40001
rect 39488 40035 39540 40044
rect 39488 40001 39497 40035
rect 39497 40001 39531 40035
rect 39531 40001 39540 40035
rect 39488 39992 39540 40001
rect 40500 40035 40552 40044
rect 40500 40001 40509 40035
rect 40509 40001 40543 40035
rect 40543 40001 40552 40035
rect 40500 39992 40552 40001
rect 41696 39992 41748 40044
rect 40224 39924 40276 39976
rect 30196 39831 30248 39840
rect 30196 39797 30205 39831
rect 30205 39797 30239 39831
rect 30239 39797 30248 39831
rect 30196 39788 30248 39797
rect 31116 39788 31168 39840
rect 32864 39831 32916 39840
rect 32864 39797 32873 39831
rect 32873 39797 32907 39831
rect 32907 39797 32916 39831
rect 32864 39788 32916 39797
rect 34520 39788 34572 39840
rect 35716 39788 35768 39840
rect 36084 39856 36136 39908
rect 39120 39856 39172 39908
rect 40040 39899 40092 39908
rect 40040 39865 40049 39899
rect 40049 39865 40083 39899
rect 40083 39865 40092 39899
rect 40040 39856 40092 39865
rect 41328 39856 41380 39908
rect 37464 39788 37516 39840
rect 39856 39788 39908 39840
rect 40960 39788 41012 39840
rect 42064 39788 42116 39840
rect 43168 39788 43220 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 11152 39627 11204 39636
rect 11152 39593 11161 39627
rect 11161 39593 11195 39627
rect 11195 39593 11204 39627
rect 11152 39584 11204 39593
rect 12808 39627 12860 39636
rect 12808 39593 12817 39627
rect 12817 39593 12851 39627
rect 12851 39593 12860 39627
rect 12808 39584 12860 39593
rect 16948 39584 17000 39636
rect 17040 39584 17092 39636
rect 13820 39448 13872 39500
rect 14464 39448 14516 39500
rect 21180 39584 21232 39636
rect 22376 39584 22428 39636
rect 24492 39584 24544 39636
rect 27068 39584 27120 39636
rect 28816 39584 28868 39636
rect 17960 39448 18012 39500
rect 18328 39448 18380 39500
rect 20352 39448 20404 39500
rect 21824 39491 21876 39500
rect 21824 39457 21833 39491
rect 21833 39457 21867 39491
rect 21867 39457 21876 39491
rect 21824 39448 21876 39457
rect 22652 39448 22704 39500
rect 23388 39448 23440 39500
rect 10876 39312 10928 39364
rect 13636 39312 13688 39364
rect 14372 39312 14424 39364
rect 15752 39380 15804 39432
rect 16120 39380 16172 39432
rect 16396 39423 16448 39432
rect 16396 39389 16405 39423
rect 16405 39389 16439 39423
rect 16439 39389 16448 39423
rect 16396 39380 16448 39389
rect 16948 39380 17000 39432
rect 17776 39423 17828 39432
rect 17776 39389 17785 39423
rect 17785 39389 17819 39423
rect 17819 39389 17828 39423
rect 17776 39380 17828 39389
rect 18052 39423 18104 39432
rect 18052 39389 18061 39423
rect 18061 39389 18095 39423
rect 18095 39389 18104 39423
rect 18052 39380 18104 39389
rect 17316 39312 17368 39364
rect 18880 39380 18932 39432
rect 20628 39423 20680 39432
rect 20628 39389 20637 39423
rect 20637 39389 20671 39423
rect 20671 39389 20680 39423
rect 20628 39380 20680 39389
rect 12256 39287 12308 39296
rect 12256 39253 12265 39287
rect 12265 39253 12299 39287
rect 12299 39253 12308 39287
rect 12256 39244 12308 39253
rect 14556 39244 14608 39296
rect 16212 39287 16264 39296
rect 16212 39253 16221 39287
rect 16221 39253 16255 39287
rect 16255 39253 16264 39287
rect 16212 39244 16264 39253
rect 19340 39287 19392 39296
rect 19340 39253 19349 39287
rect 19349 39253 19383 39287
rect 19383 39253 19392 39287
rect 19340 39244 19392 39253
rect 19432 39244 19484 39296
rect 20536 39312 20588 39364
rect 22100 39423 22152 39432
rect 22100 39389 22109 39423
rect 22109 39389 22143 39423
rect 22143 39389 22152 39423
rect 22100 39380 22152 39389
rect 23940 39516 23992 39568
rect 24860 39516 24912 39568
rect 25504 39516 25556 39568
rect 29828 39584 29880 39636
rect 34336 39584 34388 39636
rect 24584 39448 24636 39500
rect 26056 39448 26108 39500
rect 26148 39448 26200 39500
rect 27160 39448 27212 39500
rect 31392 39516 31444 39568
rect 31760 39516 31812 39568
rect 33968 39516 34020 39568
rect 35900 39584 35952 39636
rect 35992 39584 36044 39636
rect 36360 39584 36412 39636
rect 38660 39584 38712 39636
rect 38844 39584 38896 39636
rect 39028 39584 39080 39636
rect 39120 39584 39172 39636
rect 24216 39380 24268 39432
rect 25504 39423 25556 39432
rect 25504 39389 25513 39423
rect 25513 39389 25547 39423
rect 25547 39389 25556 39423
rect 25504 39380 25556 39389
rect 25596 39423 25648 39432
rect 25596 39389 25605 39423
rect 25605 39389 25639 39423
rect 25639 39389 25648 39423
rect 25596 39380 25648 39389
rect 26424 39380 26476 39432
rect 20812 39312 20864 39364
rect 25228 39312 25280 39364
rect 27344 39380 27396 39432
rect 28080 39380 28132 39432
rect 28356 39380 28408 39432
rect 31944 39448 31996 39500
rect 32680 39448 32732 39500
rect 33048 39448 33100 39500
rect 29000 39380 29052 39432
rect 20720 39244 20772 39296
rect 25044 39244 25096 39296
rect 26148 39244 26200 39296
rect 29092 39312 29144 39364
rect 30564 39380 30616 39432
rect 31576 39423 31628 39432
rect 31208 39312 31260 39364
rect 31576 39389 31585 39423
rect 31585 39389 31619 39423
rect 31619 39389 31628 39423
rect 31576 39380 31628 39389
rect 33692 39380 33744 39432
rect 33968 39423 34020 39432
rect 33968 39389 33977 39423
rect 33977 39389 34011 39423
rect 34011 39389 34020 39423
rect 33968 39380 34020 39389
rect 33140 39312 33192 39364
rect 33416 39312 33468 39364
rect 33600 39312 33652 39364
rect 34336 39380 34388 39432
rect 34980 39448 35032 39500
rect 35440 39516 35492 39568
rect 36728 39516 36780 39568
rect 40960 39516 41012 39568
rect 35348 39380 35400 39432
rect 36268 39448 36320 39500
rect 38384 39448 38436 39500
rect 35532 39380 35584 39432
rect 36360 39380 36412 39432
rect 36544 39423 36596 39432
rect 36544 39389 36553 39423
rect 36553 39389 36587 39423
rect 36587 39389 36596 39423
rect 38108 39423 38160 39432
rect 36544 39380 36596 39389
rect 38108 39389 38117 39423
rect 38117 39389 38151 39423
rect 38151 39389 38160 39423
rect 38108 39380 38160 39389
rect 30472 39244 30524 39296
rect 33508 39244 33560 39296
rect 37004 39312 37056 39364
rect 37648 39312 37700 39364
rect 43536 39448 43588 39500
rect 47124 39448 47176 39500
rect 39856 39423 39908 39432
rect 39856 39389 39865 39423
rect 39865 39389 39899 39423
rect 39899 39389 39908 39423
rect 39856 39380 39908 39389
rect 38660 39312 38712 39364
rect 39120 39355 39172 39364
rect 39120 39321 39129 39355
rect 39129 39321 39163 39355
rect 39163 39321 39172 39355
rect 39120 39312 39172 39321
rect 41512 39380 41564 39432
rect 41604 39355 41656 39364
rect 41604 39321 41613 39355
rect 41613 39321 41647 39355
rect 41647 39321 41656 39355
rect 41604 39312 41656 39321
rect 42064 39312 42116 39364
rect 35348 39287 35400 39296
rect 35348 39253 35357 39287
rect 35357 39253 35391 39287
rect 35391 39253 35400 39287
rect 35348 39244 35400 39253
rect 38752 39244 38804 39296
rect 39856 39244 39908 39296
rect 40592 39287 40644 39296
rect 40592 39253 40601 39287
rect 40601 39253 40635 39287
rect 40635 39253 40644 39287
rect 40592 39244 40644 39253
rect 42708 39287 42760 39296
rect 42708 39253 42717 39287
rect 42717 39253 42751 39287
rect 42751 39253 42760 39287
rect 42708 39244 42760 39253
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 12900 39040 12952 39092
rect 13820 39040 13872 39092
rect 14280 39083 14332 39092
rect 14280 39049 14289 39083
rect 14289 39049 14323 39083
rect 14323 39049 14332 39083
rect 14280 39040 14332 39049
rect 15844 39040 15896 39092
rect 16120 39083 16172 39092
rect 16120 39049 16129 39083
rect 16129 39049 16163 39083
rect 16163 39049 16172 39083
rect 16120 39040 16172 39049
rect 17776 39040 17828 39092
rect 19432 39040 19484 39092
rect 11152 38904 11204 38956
rect 13636 38972 13688 39024
rect 14188 38972 14240 39024
rect 14372 38972 14424 39024
rect 14464 38947 14516 38956
rect 12900 38879 12952 38888
rect 12900 38845 12909 38879
rect 12909 38845 12943 38879
rect 12943 38845 12952 38879
rect 12900 38836 12952 38845
rect 14464 38913 14473 38947
rect 14473 38913 14507 38947
rect 14507 38913 14516 38947
rect 14464 38904 14516 38913
rect 14556 38947 14608 38956
rect 14556 38913 14565 38947
rect 14565 38913 14599 38947
rect 14599 38913 14608 38947
rect 14556 38904 14608 38913
rect 15016 38904 15068 38956
rect 18880 38972 18932 39024
rect 19340 38972 19392 39024
rect 20996 39040 21048 39092
rect 20628 38972 20680 39024
rect 23112 39040 23164 39092
rect 23572 39083 23624 39092
rect 23572 39049 23581 39083
rect 23581 39049 23615 39083
rect 23615 39049 23624 39083
rect 23572 39040 23624 39049
rect 14280 38879 14332 38888
rect 14280 38845 14289 38879
rect 14289 38845 14323 38879
rect 14323 38845 14332 38879
rect 14280 38836 14332 38845
rect 10232 38700 10284 38752
rect 10876 38743 10928 38752
rect 10876 38709 10885 38743
rect 10885 38709 10919 38743
rect 10919 38709 10928 38743
rect 10876 38700 10928 38709
rect 12256 38743 12308 38752
rect 12256 38709 12265 38743
rect 12265 38709 12299 38743
rect 12299 38709 12308 38743
rect 15384 38904 15436 38956
rect 16028 38904 16080 38956
rect 18604 38904 18656 38956
rect 20076 38947 20128 38956
rect 20076 38913 20085 38947
rect 20085 38913 20119 38947
rect 20119 38913 20128 38947
rect 20076 38904 20128 38913
rect 20812 38904 20864 38956
rect 15936 38836 15988 38888
rect 16396 38836 16448 38888
rect 19248 38879 19300 38888
rect 19248 38845 19257 38879
rect 19257 38845 19291 38879
rect 19291 38845 19300 38879
rect 19248 38836 19300 38845
rect 19340 38768 19392 38820
rect 20812 38768 20864 38820
rect 21916 38904 21968 38956
rect 22008 38879 22060 38888
rect 22008 38845 22017 38879
rect 22017 38845 22051 38879
rect 22051 38845 22060 38879
rect 22008 38836 22060 38845
rect 23296 38972 23348 39024
rect 23020 38947 23072 38956
rect 23020 38913 23029 38947
rect 23029 38913 23063 38947
rect 23063 38913 23072 38947
rect 24032 38972 24084 39024
rect 25596 39040 25648 39092
rect 28356 39083 28408 39092
rect 28356 39049 28365 39083
rect 28365 39049 28399 39083
rect 28399 39049 28408 39083
rect 28356 39040 28408 39049
rect 28448 39040 28500 39092
rect 24860 39015 24912 39024
rect 24860 38981 24869 39015
rect 24869 38981 24903 39015
rect 24903 38981 24912 39015
rect 25504 39015 25556 39024
rect 24860 38972 24912 38981
rect 25504 38981 25513 39015
rect 25513 38981 25547 39015
rect 25547 38981 25556 39015
rect 25504 38972 25556 38981
rect 23020 38904 23072 38913
rect 24308 38904 24360 38956
rect 24768 38904 24820 38956
rect 28264 38904 28316 38956
rect 28632 38947 28684 38956
rect 28632 38913 28641 38947
rect 28641 38913 28675 38947
rect 28675 38913 28684 38947
rect 28632 38904 28684 38913
rect 28816 38904 28868 38956
rect 29736 38947 29788 38956
rect 17040 38743 17092 38752
rect 12256 38700 12308 38709
rect 17040 38709 17049 38743
rect 17049 38709 17083 38743
rect 17083 38709 17092 38743
rect 17040 38700 17092 38709
rect 18328 38700 18380 38752
rect 19156 38700 19208 38752
rect 19616 38743 19668 38752
rect 19616 38709 19625 38743
rect 19625 38709 19659 38743
rect 19659 38709 19668 38743
rect 19616 38700 19668 38709
rect 21088 38700 21140 38752
rect 23664 38836 23716 38888
rect 24492 38836 24544 38888
rect 22744 38743 22796 38752
rect 22744 38709 22753 38743
rect 22753 38709 22787 38743
rect 22787 38709 22796 38743
rect 22744 38700 22796 38709
rect 24584 38700 24636 38752
rect 24768 38700 24820 38752
rect 27528 38836 27580 38888
rect 28448 38836 28500 38888
rect 29736 38913 29745 38947
rect 29745 38913 29779 38947
rect 29779 38913 29788 38947
rect 29736 38904 29788 38913
rect 29644 38879 29696 38888
rect 29644 38845 29653 38879
rect 29653 38845 29687 38879
rect 29687 38845 29696 38879
rect 29644 38836 29696 38845
rect 30564 39040 30616 39092
rect 30564 38904 30616 38956
rect 30748 38904 30800 38956
rect 31944 39040 31996 39092
rect 32404 39040 32456 39092
rect 33416 39040 33468 39092
rect 37648 39040 37700 39092
rect 32772 38972 32824 39024
rect 33508 39015 33560 39024
rect 33508 38981 33517 39015
rect 33517 38981 33551 39015
rect 33551 38981 33560 39015
rect 33508 38972 33560 38981
rect 33600 38972 33652 39024
rect 34428 38972 34480 39024
rect 38936 39040 38988 39092
rect 39856 39083 39908 39092
rect 39856 39049 39865 39083
rect 39865 39049 39899 39083
rect 39899 39049 39908 39083
rect 39856 39040 39908 39049
rect 43536 39083 43588 39092
rect 43536 39049 43545 39083
rect 43545 39049 43579 39083
rect 43579 39049 43588 39083
rect 43536 39040 43588 39049
rect 31760 38904 31812 38956
rect 32496 38904 32548 38956
rect 33692 38904 33744 38956
rect 34152 38904 34204 38956
rect 36176 38947 36228 38956
rect 31392 38836 31444 38888
rect 31576 38836 31628 38888
rect 34244 38836 34296 38888
rect 36176 38913 36185 38947
rect 36185 38913 36219 38947
rect 36219 38913 36228 38947
rect 36176 38904 36228 38913
rect 36452 38904 36504 38956
rect 38568 39015 38620 39024
rect 38568 38981 38577 39015
rect 38577 38981 38611 39015
rect 38611 38981 38620 39015
rect 38568 38972 38620 38981
rect 38660 38972 38712 39024
rect 39488 38972 39540 39024
rect 43168 38972 43220 39024
rect 35716 38836 35768 38888
rect 39028 38904 39080 38956
rect 40224 38947 40276 38956
rect 38108 38836 38160 38888
rect 40224 38913 40233 38947
rect 40233 38913 40267 38947
rect 40267 38913 40276 38947
rect 40224 38904 40276 38913
rect 40868 38904 40920 38956
rect 42708 38836 42760 38888
rect 28172 38768 28224 38820
rect 26240 38700 26292 38752
rect 27252 38700 27304 38752
rect 29092 38768 29144 38820
rect 29460 38768 29512 38820
rect 32404 38768 32456 38820
rect 32864 38768 32916 38820
rect 33692 38768 33744 38820
rect 38016 38768 38068 38820
rect 30564 38700 30616 38752
rect 31300 38700 31352 38752
rect 32312 38700 32364 38752
rect 33600 38700 33652 38752
rect 34336 38743 34388 38752
rect 34336 38709 34345 38743
rect 34345 38709 34379 38743
rect 34379 38709 34388 38743
rect 34336 38700 34388 38709
rect 35440 38700 35492 38752
rect 35716 38743 35768 38752
rect 35716 38709 35725 38743
rect 35725 38709 35759 38743
rect 35759 38709 35768 38743
rect 35716 38700 35768 38709
rect 36268 38743 36320 38752
rect 36268 38709 36277 38743
rect 36277 38709 36311 38743
rect 36311 38709 36320 38743
rect 36268 38700 36320 38709
rect 38200 38700 38252 38752
rect 39672 38700 39724 38752
rect 42708 38700 42760 38752
rect 42984 38743 43036 38752
rect 42984 38709 42993 38743
rect 42993 38709 43027 38743
rect 43027 38709 43036 38743
rect 42984 38700 43036 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 11152 38496 11204 38548
rect 14096 38496 14148 38548
rect 14464 38496 14516 38548
rect 16672 38539 16724 38548
rect 13452 38428 13504 38480
rect 15660 38428 15712 38480
rect 15752 38403 15804 38412
rect 15752 38369 15761 38403
rect 15761 38369 15795 38403
rect 15795 38369 15804 38403
rect 15752 38360 15804 38369
rect 16672 38505 16681 38539
rect 16681 38505 16715 38539
rect 16715 38505 16724 38539
rect 16672 38496 16724 38505
rect 17040 38496 17092 38548
rect 19248 38496 19300 38548
rect 20352 38496 20404 38548
rect 20536 38539 20588 38548
rect 20536 38505 20545 38539
rect 20545 38505 20579 38539
rect 20579 38505 20588 38539
rect 20536 38496 20588 38505
rect 21916 38496 21968 38548
rect 22744 38496 22796 38548
rect 22836 38496 22888 38548
rect 23204 38496 23256 38548
rect 23848 38539 23900 38548
rect 23848 38505 23857 38539
rect 23857 38505 23891 38539
rect 23891 38505 23900 38539
rect 23848 38496 23900 38505
rect 25320 38496 25372 38548
rect 25412 38496 25464 38548
rect 27804 38496 27856 38548
rect 27988 38539 28040 38548
rect 27988 38505 27997 38539
rect 27997 38505 28031 38539
rect 28031 38505 28040 38539
rect 27988 38496 28040 38505
rect 29644 38496 29696 38548
rect 30380 38496 30432 38548
rect 32864 38496 32916 38548
rect 16028 38428 16080 38480
rect 18604 38471 18656 38480
rect 18604 38437 18613 38471
rect 18613 38437 18647 38471
rect 18647 38437 18656 38471
rect 18604 38428 18656 38437
rect 19156 38428 19208 38480
rect 21824 38428 21876 38480
rect 23020 38428 23072 38480
rect 16488 38360 16540 38412
rect 12256 38292 12308 38344
rect 12532 38292 12584 38344
rect 15108 38292 15160 38344
rect 15292 38292 15344 38344
rect 16856 38335 16908 38344
rect 1584 38224 1636 38276
rect 12440 38199 12492 38208
rect 12440 38165 12449 38199
rect 12449 38165 12483 38199
rect 12483 38165 12492 38199
rect 13820 38224 13872 38276
rect 14648 38224 14700 38276
rect 15476 38224 15528 38276
rect 16856 38301 16865 38335
rect 16865 38301 16899 38335
rect 16899 38301 16908 38335
rect 16856 38292 16908 38301
rect 17592 38335 17644 38344
rect 17592 38301 17601 38335
rect 17601 38301 17635 38335
rect 17635 38301 17644 38335
rect 17592 38292 17644 38301
rect 18144 38360 18196 38412
rect 18236 38360 18288 38412
rect 18512 38292 18564 38344
rect 19892 38292 19944 38344
rect 20168 38292 20220 38344
rect 20444 38335 20496 38344
rect 20444 38301 20453 38335
rect 20453 38301 20487 38335
rect 20487 38301 20496 38335
rect 20444 38292 20496 38301
rect 20720 38292 20772 38344
rect 21916 38335 21968 38344
rect 21916 38301 21925 38335
rect 21925 38301 21959 38335
rect 21959 38301 21968 38335
rect 21916 38292 21968 38301
rect 22284 38292 22336 38344
rect 16212 38224 16264 38276
rect 18144 38224 18196 38276
rect 18972 38224 19024 38276
rect 22836 38224 22888 38276
rect 23296 38292 23348 38344
rect 23480 38292 23532 38344
rect 26332 38360 26384 38412
rect 27068 38360 27120 38412
rect 27712 38428 27764 38480
rect 28448 38428 28500 38480
rect 29000 38403 29052 38412
rect 29000 38369 29009 38403
rect 29009 38369 29043 38403
rect 29043 38369 29052 38403
rect 29000 38360 29052 38369
rect 33600 38428 33652 38480
rect 33968 38496 34020 38548
rect 42616 38539 42668 38548
rect 42616 38505 42625 38539
rect 42625 38505 42659 38539
rect 42659 38505 42668 38539
rect 42616 38496 42668 38505
rect 36360 38428 36412 38480
rect 12440 38156 12492 38165
rect 13176 38156 13228 38208
rect 16028 38156 16080 38208
rect 16120 38199 16172 38208
rect 16120 38165 16129 38199
rect 16129 38165 16163 38199
rect 16163 38165 16172 38199
rect 17040 38199 17092 38208
rect 16120 38156 16172 38165
rect 17040 38165 17049 38199
rect 17049 38165 17083 38199
rect 17083 38165 17092 38199
rect 17040 38156 17092 38165
rect 17960 38156 18012 38208
rect 21824 38156 21876 38208
rect 23112 38199 23164 38208
rect 23112 38165 23137 38199
rect 23137 38165 23164 38199
rect 23112 38156 23164 38165
rect 23296 38156 23348 38208
rect 24308 38156 24360 38208
rect 24768 38335 24820 38344
rect 24768 38301 24777 38335
rect 24777 38301 24811 38335
rect 24811 38301 24820 38335
rect 24768 38292 24820 38301
rect 24952 38335 25004 38344
rect 24952 38301 24961 38335
rect 24961 38301 24995 38335
rect 24995 38301 25004 38335
rect 24952 38292 25004 38301
rect 25412 38292 25464 38344
rect 26700 38292 26752 38344
rect 27252 38335 27304 38344
rect 27252 38301 27261 38335
rect 27261 38301 27295 38335
rect 27295 38301 27304 38335
rect 27252 38292 27304 38301
rect 27436 38335 27488 38344
rect 27436 38301 27445 38335
rect 27445 38301 27479 38335
rect 27479 38301 27488 38335
rect 27436 38292 27488 38301
rect 27620 38335 27672 38344
rect 27620 38301 27629 38335
rect 27629 38301 27663 38335
rect 27663 38301 27672 38335
rect 27620 38292 27672 38301
rect 27804 38335 27856 38344
rect 27804 38301 27813 38335
rect 27813 38301 27847 38335
rect 27847 38301 27856 38335
rect 27804 38292 27856 38301
rect 28632 38292 28684 38344
rect 29644 38335 29696 38344
rect 29644 38301 29653 38335
rect 29653 38301 29687 38335
rect 29687 38301 29696 38335
rect 29644 38292 29696 38301
rect 29736 38335 29788 38344
rect 29736 38301 29745 38335
rect 29745 38301 29779 38335
rect 29779 38301 29788 38335
rect 31392 38360 31444 38412
rect 29736 38292 29788 38301
rect 30196 38292 30248 38344
rect 28448 38224 28500 38276
rect 33232 38360 33284 38412
rect 35072 38403 35124 38412
rect 32772 38335 32824 38344
rect 32772 38301 32781 38335
rect 32781 38301 32815 38335
rect 32815 38301 32824 38335
rect 33048 38335 33100 38344
rect 32772 38292 32824 38301
rect 33048 38301 33057 38335
rect 33057 38301 33091 38335
rect 33091 38301 33100 38335
rect 33048 38292 33100 38301
rect 33140 38292 33192 38344
rect 33692 38292 33744 38344
rect 35072 38369 35081 38403
rect 35081 38369 35115 38403
rect 35115 38369 35124 38403
rect 35072 38360 35124 38369
rect 35348 38360 35400 38412
rect 35716 38360 35768 38412
rect 37372 38360 37424 38412
rect 38568 38360 38620 38412
rect 42984 38428 43036 38480
rect 25964 38156 26016 38208
rect 26240 38156 26292 38208
rect 29552 38156 29604 38208
rect 29736 38156 29788 38208
rect 32956 38156 33008 38208
rect 33416 38224 33468 38276
rect 34888 38224 34940 38276
rect 35348 38224 35400 38276
rect 36084 38335 36136 38344
rect 36084 38301 36093 38335
rect 36093 38301 36127 38335
rect 36127 38301 36136 38335
rect 36084 38292 36136 38301
rect 36268 38292 36320 38344
rect 38108 38335 38160 38344
rect 38108 38301 38117 38335
rect 38117 38301 38151 38335
rect 38151 38301 38160 38335
rect 38108 38292 38160 38301
rect 38200 38335 38252 38344
rect 38200 38301 38209 38335
rect 38209 38301 38243 38335
rect 38243 38301 38252 38335
rect 38752 38335 38804 38344
rect 38200 38292 38252 38301
rect 38752 38301 38761 38335
rect 38761 38301 38795 38335
rect 38795 38301 38804 38335
rect 38752 38292 38804 38301
rect 38936 38335 38988 38344
rect 38936 38301 38945 38335
rect 38945 38301 38979 38335
rect 38979 38301 38988 38335
rect 38936 38292 38988 38301
rect 40592 38292 40644 38344
rect 34796 38156 34848 38208
rect 34980 38156 35032 38208
rect 35808 38156 35860 38208
rect 37832 38224 37884 38276
rect 42708 38292 42760 38344
rect 43352 38292 43404 38344
rect 42156 38224 42208 38276
rect 39672 38156 39724 38208
rect 39856 38199 39908 38208
rect 39856 38165 39865 38199
rect 39865 38165 39899 38199
rect 39899 38165 39908 38199
rect 39856 38156 39908 38165
rect 43168 38199 43220 38208
rect 43168 38165 43177 38199
rect 43177 38165 43211 38199
rect 43211 38165 43220 38199
rect 43168 38156 43220 38165
rect 48044 38199 48096 38208
rect 48044 38165 48053 38199
rect 48053 38165 48087 38199
rect 48087 38165 48096 38199
rect 48044 38156 48096 38165
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 1584 37995 1636 38004
rect 1584 37961 1593 37995
rect 1593 37961 1627 37995
rect 1627 37961 1636 37995
rect 1584 37952 1636 37961
rect 12440 37952 12492 38004
rect 14188 37952 14240 38004
rect 16856 37995 16908 38004
rect 16856 37961 16858 37995
rect 16858 37961 16892 37995
rect 16892 37961 16908 37995
rect 16856 37952 16908 37961
rect 17224 37952 17276 38004
rect 13268 37884 13320 37936
rect 13452 37927 13504 37936
rect 13452 37893 13461 37927
rect 13461 37893 13495 37927
rect 13495 37893 13504 37927
rect 13452 37884 13504 37893
rect 13544 37884 13596 37936
rect 14556 37927 14608 37936
rect 13912 37859 13964 37868
rect 13912 37825 13921 37859
rect 13921 37825 13955 37859
rect 13955 37825 13964 37859
rect 13912 37816 13964 37825
rect 14556 37893 14565 37927
rect 14565 37893 14599 37927
rect 14599 37893 14608 37927
rect 14556 37884 14608 37893
rect 16488 37884 16540 37936
rect 18144 37952 18196 38004
rect 21456 37952 21508 38004
rect 23204 37952 23256 38004
rect 23848 37952 23900 38004
rect 24400 37952 24452 38004
rect 25688 37952 25740 38004
rect 29920 37952 29972 38004
rect 30104 37995 30156 38004
rect 30104 37961 30113 37995
rect 30113 37961 30147 37995
rect 30147 37961 30156 37995
rect 30104 37952 30156 37961
rect 30288 37952 30340 38004
rect 23296 37884 23348 37936
rect 27160 37927 27212 37936
rect 14280 37859 14332 37868
rect 14280 37825 14289 37859
rect 14289 37825 14323 37859
rect 14323 37825 14332 37859
rect 15200 37859 15252 37868
rect 14280 37816 14332 37825
rect 15200 37825 15209 37859
rect 15209 37825 15243 37859
rect 15243 37825 15252 37859
rect 15200 37816 15252 37825
rect 15476 37859 15528 37868
rect 15476 37825 15485 37859
rect 15485 37825 15519 37859
rect 15519 37825 15528 37859
rect 15476 37816 15528 37825
rect 16672 37859 16724 37868
rect 16672 37825 16681 37859
rect 16681 37825 16715 37859
rect 16715 37825 16724 37859
rect 16672 37816 16724 37825
rect 16948 37859 17000 37868
rect 16948 37825 16957 37859
rect 16957 37825 16991 37859
rect 16991 37825 17000 37859
rect 16948 37816 17000 37825
rect 17868 37859 17920 37868
rect 17868 37825 17877 37859
rect 17877 37825 17911 37859
rect 17911 37825 17920 37859
rect 17868 37816 17920 37825
rect 18972 37859 19024 37868
rect 18972 37825 18981 37859
rect 18981 37825 19015 37859
rect 19015 37825 19024 37859
rect 18972 37816 19024 37825
rect 20352 37859 20404 37868
rect 20352 37825 20361 37859
rect 20361 37825 20395 37859
rect 20395 37825 20404 37859
rect 20352 37816 20404 37825
rect 15292 37791 15344 37800
rect 12900 37680 12952 37732
rect 14924 37680 14976 37732
rect 15292 37757 15301 37791
rect 15301 37757 15335 37791
rect 15335 37757 15344 37791
rect 15292 37748 15344 37757
rect 17684 37748 17736 37800
rect 18696 37791 18748 37800
rect 10324 37612 10376 37664
rect 13176 37612 13228 37664
rect 17224 37680 17276 37732
rect 18696 37757 18705 37791
rect 18705 37757 18739 37791
rect 18739 37757 18748 37791
rect 18696 37748 18748 37757
rect 22468 37816 22520 37868
rect 24032 37816 24084 37868
rect 24216 37859 24268 37868
rect 24216 37825 24225 37859
rect 24225 37825 24259 37859
rect 24259 37825 24268 37859
rect 24216 37816 24268 37825
rect 24492 37859 24544 37868
rect 24492 37825 24501 37859
rect 24501 37825 24535 37859
rect 24535 37825 24544 37859
rect 24492 37816 24544 37825
rect 24676 37859 24728 37868
rect 24676 37825 24685 37859
rect 24685 37825 24719 37859
rect 24719 37825 24728 37859
rect 24676 37816 24728 37825
rect 21732 37748 21784 37800
rect 21824 37748 21876 37800
rect 18144 37680 18196 37732
rect 18236 37723 18288 37732
rect 18236 37689 18245 37723
rect 18245 37689 18279 37723
rect 18279 37689 18288 37723
rect 18236 37680 18288 37689
rect 15752 37612 15804 37664
rect 16028 37655 16080 37664
rect 16028 37621 16037 37655
rect 16037 37621 16071 37655
rect 16071 37621 16080 37655
rect 16028 37612 16080 37621
rect 16120 37612 16172 37664
rect 21640 37680 21692 37732
rect 22192 37748 22244 37800
rect 23112 37748 23164 37800
rect 24400 37791 24452 37800
rect 24400 37757 24409 37791
rect 24409 37757 24443 37791
rect 24443 37757 24452 37791
rect 24584 37791 24636 37800
rect 24400 37748 24452 37757
rect 24584 37757 24593 37791
rect 24593 37757 24627 37791
rect 24627 37757 24636 37791
rect 24584 37748 24636 37757
rect 24860 37816 24912 37868
rect 25964 37859 26016 37868
rect 25964 37825 25973 37859
rect 25973 37825 26007 37859
rect 26007 37825 26016 37859
rect 25964 37816 26016 37825
rect 27160 37893 27169 37927
rect 27169 37893 27203 37927
rect 27203 37893 27212 37927
rect 27160 37884 27212 37893
rect 26424 37816 26476 37868
rect 24860 37680 24912 37732
rect 29000 37884 29052 37936
rect 28356 37859 28408 37868
rect 28356 37825 28365 37859
rect 28365 37825 28399 37859
rect 28399 37825 28408 37859
rect 28356 37816 28408 37825
rect 28632 37816 28684 37868
rect 29552 37816 29604 37868
rect 30288 37859 30340 37868
rect 30288 37825 30297 37859
rect 30297 37825 30331 37859
rect 30331 37825 30340 37859
rect 30288 37816 30340 37825
rect 30564 37816 30616 37868
rect 30748 37816 30800 37868
rect 30932 37859 30984 37868
rect 30932 37825 30941 37859
rect 30941 37825 30975 37859
rect 30975 37825 30984 37859
rect 30932 37816 30984 37825
rect 31300 37816 31352 37868
rect 32036 37816 32088 37868
rect 33048 37952 33100 38004
rect 33140 37952 33192 38004
rect 33508 37952 33560 38004
rect 34888 37995 34940 38004
rect 34888 37961 34897 37995
rect 34897 37961 34931 37995
rect 34931 37961 34940 37995
rect 34888 37952 34940 37961
rect 35716 37952 35768 38004
rect 37464 37952 37516 38004
rect 38384 37952 38436 38004
rect 41052 37952 41104 38004
rect 41696 37995 41748 38004
rect 41696 37961 41705 37995
rect 41705 37961 41739 37995
rect 41739 37961 41748 37995
rect 41696 37952 41748 37961
rect 42984 37952 43036 38004
rect 34336 37884 34388 37936
rect 35532 37884 35584 37936
rect 38108 37884 38160 37936
rect 32588 37859 32640 37868
rect 32588 37825 32597 37859
rect 32597 37825 32631 37859
rect 32631 37825 32640 37859
rect 32588 37816 32640 37825
rect 32772 37859 32824 37868
rect 32772 37825 32781 37859
rect 32781 37825 32815 37859
rect 32815 37825 32824 37859
rect 32772 37816 32824 37825
rect 33508 37816 33560 37868
rect 34520 37816 34572 37868
rect 36176 37859 36228 37868
rect 28448 37748 28500 37800
rect 30012 37748 30064 37800
rect 36176 37825 36185 37859
rect 36185 37825 36219 37859
rect 36219 37825 36228 37859
rect 36176 37816 36228 37825
rect 36268 37816 36320 37868
rect 37464 37859 37516 37868
rect 35992 37748 36044 37800
rect 36544 37748 36596 37800
rect 37464 37825 37473 37859
rect 37473 37825 37507 37859
rect 37507 37825 37516 37859
rect 37464 37816 37516 37825
rect 39120 37816 39172 37868
rect 40132 37816 40184 37868
rect 37556 37748 37608 37800
rect 38476 37791 38528 37800
rect 38476 37757 38485 37791
rect 38485 37757 38519 37791
rect 38519 37757 38528 37791
rect 38476 37748 38528 37757
rect 41144 37748 41196 37800
rect 28356 37680 28408 37732
rect 19892 37655 19944 37664
rect 19892 37621 19901 37655
rect 19901 37621 19935 37655
rect 19935 37621 19944 37655
rect 19892 37612 19944 37621
rect 20628 37655 20680 37664
rect 20628 37621 20637 37655
rect 20637 37621 20671 37655
rect 20671 37621 20680 37655
rect 20628 37612 20680 37621
rect 20812 37655 20864 37664
rect 20812 37621 20821 37655
rect 20821 37621 20855 37655
rect 20855 37621 20864 37655
rect 20812 37612 20864 37621
rect 21824 37655 21876 37664
rect 21824 37621 21833 37655
rect 21833 37621 21867 37655
rect 21867 37621 21876 37655
rect 21824 37612 21876 37621
rect 22008 37612 22060 37664
rect 24124 37612 24176 37664
rect 24400 37612 24452 37664
rect 25780 37612 25832 37664
rect 26056 37612 26108 37664
rect 28448 37612 28500 37664
rect 30196 37680 30248 37732
rect 32680 37680 32732 37732
rect 34060 37680 34112 37732
rect 37372 37680 37424 37732
rect 39212 37723 39264 37732
rect 39212 37689 39221 37723
rect 39221 37689 39255 37723
rect 39255 37689 39264 37723
rect 39212 37680 39264 37689
rect 33600 37655 33652 37664
rect 33600 37621 33609 37655
rect 33609 37621 33643 37655
rect 33643 37621 33652 37655
rect 33600 37612 33652 37621
rect 33692 37612 33744 37664
rect 37832 37612 37884 37664
rect 39028 37612 39080 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 11796 37408 11848 37460
rect 13820 37408 13872 37460
rect 10968 37383 11020 37392
rect 10968 37349 10977 37383
rect 10977 37349 11011 37383
rect 11011 37349 11020 37383
rect 10968 37340 11020 37349
rect 12440 37340 12492 37392
rect 15200 37408 15252 37460
rect 16488 37408 16540 37460
rect 16948 37408 17000 37460
rect 18052 37408 18104 37460
rect 19156 37408 19208 37460
rect 20536 37408 20588 37460
rect 21824 37408 21876 37460
rect 22100 37408 22152 37460
rect 23940 37408 23992 37460
rect 24768 37408 24820 37460
rect 25688 37451 25740 37460
rect 25688 37417 25697 37451
rect 25697 37417 25731 37451
rect 25731 37417 25740 37451
rect 25688 37408 25740 37417
rect 10324 37315 10376 37324
rect 10324 37281 10333 37315
rect 10333 37281 10367 37315
rect 10367 37281 10376 37315
rect 16304 37340 16356 37392
rect 19064 37340 19116 37392
rect 10324 37272 10376 37281
rect 12440 37204 12492 37256
rect 13452 37204 13504 37256
rect 14188 37247 14240 37256
rect 14188 37213 14197 37247
rect 14197 37213 14231 37247
rect 14231 37213 14240 37247
rect 14188 37204 14240 37213
rect 16948 37272 17000 37324
rect 18420 37272 18472 37324
rect 19248 37272 19300 37324
rect 20812 37340 20864 37392
rect 21640 37383 21692 37392
rect 21640 37349 21649 37383
rect 21649 37349 21683 37383
rect 21683 37349 21692 37383
rect 21640 37340 21692 37349
rect 23112 37340 23164 37392
rect 15016 37247 15068 37256
rect 13176 37179 13228 37188
rect 13176 37145 13185 37179
rect 13185 37145 13219 37179
rect 13219 37145 13228 37179
rect 13176 37136 13228 37145
rect 12532 37068 12584 37120
rect 13912 37136 13964 37188
rect 15016 37213 15025 37247
rect 15025 37213 15059 37247
rect 15059 37213 15068 37247
rect 15016 37204 15068 37213
rect 15384 37204 15436 37256
rect 17500 37247 17552 37256
rect 14096 37068 14148 37120
rect 15200 37068 15252 37120
rect 17224 37136 17276 37188
rect 17500 37213 17509 37247
rect 17509 37213 17543 37247
rect 17543 37213 17552 37247
rect 17500 37204 17552 37213
rect 18512 37204 18564 37256
rect 20352 37272 20404 37324
rect 21548 37315 21600 37324
rect 21548 37281 21557 37315
rect 21557 37281 21591 37315
rect 21591 37281 21600 37315
rect 21548 37272 21600 37281
rect 22100 37272 22152 37324
rect 23388 37272 23440 37324
rect 18880 37136 18932 37188
rect 20444 37213 20453 37234
rect 20453 37213 20487 37234
rect 20487 37213 20496 37234
rect 20444 37182 20496 37213
rect 20536 37207 20564 37234
rect 20564 37207 20588 37234
rect 20536 37182 20588 37207
rect 21456 37247 21508 37256
rect 21456 37213 21465 37247
rect 21465 37213 21499 37247
rect 21499 37213 21508 37247
rect 21456 37204 21508 37213
rect 21732 37247 21784 37256
rect 21732 37213 21741 37247
rect 21741 37213 21775 37247
rect 21775 37213 21784 37247
rect 21732 37204 21784 37213
rect 23020 37247 23072 37256
rect 23020 37213 23029 37247
rect 23029 37213 23063 37247
rect 23063 37213 23072 37247
rect 23020 37204 23072 37213
rect 23848 37340 23900 37392
rect 24124 37340 24176 37392
rect 24308 37340 24360 37392
rect 24492 37315 24544 37324
rect 24492 37281 24501 37315
rect 24501 37281 24535 37315
rect 24535 37281 24544 37315
rect 24492 37272 24544 37281
rect 25136 37340 25188 37392
rect 25412 37340 25464 37392
rect 26332 37408 26384 37460
rect 27160 37408 27212 37460
rect 28172 37408 28224 37460
rect 28540 37408 28592 37460
rect 23848 37247 23900 37256
rect 23848 37213 23857 37247
rect 23857 37213 23891 37247
rect 23891 37213 23900 37247
rect 23848 37204 23900 37213
rect 24400 37247 24452 37256
rect 24400 37213 24409 37247
rect 24409 37213 24443 37247
rect 24443 37213 24452 37247
rect 24400 37204 24452 37213
rect 26056 37272 26108 37324
rect 27068 37315 27120 37324
rect 27068 37281 27077 37315
rect 27077 37281 27111 37315
rect 27111 37281 27120 37315
rect 27068 37272 27120 37281
rect 27804 37340 27856 37392
rect 28356 37340 28408 37392
rect 27712 37272 27764 37324
rect 16948 37068 17000 37120
rect 17776 37068 17828 37120
rect 20168 37068 20220 37120
rect 20628 37068 20680 37120
rect 22192 37068 22244 37120
rect 22836 37111 22888 37120
rect 22836 37077 22845 37111
rect 22845 37077 22879 37111
rect 22879 37077 22888 37111
rect 22836 37068 22888 37077
rect 25964 37204 26016 37256
rect 26976 37247 27028 37256
rect 26976 37213 26985 37247
rect 26985 37213 27019 37247
rect 27019 37213 27028 37247
rect 26976 37204 27028 37213
rect 30196 37340 30248 37392
rect 30104 37272 30156 37324
rect 27988 37204 28040 37256
rect 28448 37247 28500 37256
rect 28448 37213 28457 37247
rect 28457 37213 28491 37247
rect 28491 37213 28500 37247
rect 28448 37204 28500 37213
rect 28632 37247 28684 37256
rect 28632 37213 28641 37247
rect 28641 37213 28675 37247
rect 28675 37213 28684 37247
rect 28632 37204 28684 37213
rect 28724 37204 28776 37256
rect 32588 37408 32640 37460
rect 33416 37408 33468 37460
rect 35348 37408 35400 37460
rect 36636 37408 36688 37460
rect 37924 37408 37976 37460
rect 40592 37408 40644 37460
rect 41144 37451 41196 37460
rect 41144 37417 41153 37451
rect 41153 37417 41187 37451
rect 41187 37417 41196 37451
rect 41144 37408 41196 37417
rect 43352 37451 43404 37460
rect 37372 37383 37424 37392
rect 31024 37272 31076 37324
rect 31760 37272 31812 37324
rect 29736 37136 29788 37188
rect 30380 37247 30432 37256
rect 30380 37213 30389 37247
rect 30389 37213 30423 37247
rect 30423 37213 30432 37247
rect 30380 37204 30432 37213
rect 30748 37204 30800 37256
rect 31392 37247 31444 37256
rect 31392 37213 31401 37247
rect 31401 37213 31435 37247
rect 31435 37213 31444 37247
rect 31392 37204 31444 37213
rect 32036 37247 32088 37256
rect 32036 37213 32045 37247
rect 32045 37213 32079 37247
rect 32079 37213 32088 37247
rect 32036 37204 32088 37213
rect 34060 37272 34112 37324
rect 34336 37272 34388 37324
rect 36728 37272 36780 37324
rect 32496 37136 32548 37188
rect 32864 37179 32916 37188
rect 32864 37145 32889 37179
rect 32889 37145 32916 37179
rect 33692 37247 33744 37256
rect 33692 37213 33701 37247
rect 33701 37213 33735 37247
rect 33735 37213 33744 37247
rect 33692 37204 33744 37213
rect 33876 37247 33928 37256
rect 33876 37213 33885 37247
rect 33885 37213 33919 37247
rect 33919 37213 33928 37247
rect 33876 37204 33928 37213
rect 34244 37204 34296 37256
rect 35808 37204 35860 37256
rect 36452 37247 36504 37256
rect 36452 37213 36461 37247
rect 36461 37213 36495 37247
rect 36495 37213 36504 37247
rect 36452 37204 36504 37213
rect 37372 37349 37381 37383
rect 37381 37349 37415 37383
rect 37415 37349 37424 37383
rect 37372 37340 37424 37349
rect 38108 37340 38160 37392
rect 37280 37272 37332 37324
rect 41236 37340 41288 37392
rect 37464 37204 37516 37256
rect 38568 37204 38620 37256
rect 39120 37247 39172 37256
rect 39120 37213 39129 37247
rect 39129 37213 39163 37247
rect 39163 37213 39172 37247
rect 39120 37204 39172 37213
rect 34152 37179 34204 37188
rect 32864 37136 32916 37145
rect 28540 37111 28592 37120
rect 28540 37077 28549 37111
rect 28549 37077 28583 37111
rect 28583 37077 28592 37111
rect 28540 37068 28592 37077
rect 29828 37068 29880 37120
rect 33508 37068 33560 37120
rect 34152 37145 34161 37179
rect 34161 37145 34195 37179
rect 34195 37145 34204 37179
rect 34152 37136 34204 37145
rect 36268 37136 36320 37188
rect 37096 37136 37148 37188
rect 37556 37136 37608 37188
rect 39488 37204 39540 37256
rect 39948 37204 40000 37256
rect 40132 37136 40184 37188
rect 40776 37204 40828 37256
rect 43352 37417 43361 37451
rect 43361 37417 43395 37451
rect 43395 37417 43404 37451
rect 43352 37408 43404 37417
rect 42156 37383 42208 37392
rect 42156 37349 42165 37383
rect 42165 37349 42199 37383
rect 42199 37349 42208 37383
rect 42156 37340 42208 37349
rect 34704 37068 34756 37120
rect 35624 37111 35676 37120
rect 35624 37077 35633 37111
rect 35633 37077 35667 37111
rect 35667 37077 35676 37111
rect 35624 37068 35676 37077
rect 35808 37111 35860 37120
rect 35808 37077 35835 37111
rect 35835 37077 35860 37111
rect 35808 37068 35860 37077
rect 40040 37111 40092 37120
rect 40040 37077 40049 37111
rect 40049 37077 40083 37111
rect 40083 37077 40092 37111
rect 40040 37068 40092 37077
rect 40224 37068 40276 37120
rect 47768 37068 47820 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 10968 36907 11020 36916
rect 10968 36873 10977 36907
rect 10977 36873 11011 36907
rect 11011 36873 11020 36907
rect 10968 36864 11020 36873
rect 12440 36907 12492 36916
rect 12440 36873 12449 36907
rect 12449 36873 12483 36907
rect 12483 36873 12492 36907
rect 13544 36907 13596 36916
rect 12440 36864 12492 36873
rect 13544 36873 13553 36907
rect 13553 36873 13587 36907
rect 13587 36873 13596 36907
rect 13544 36864 13596 36873
rect 14648 36864 14700 36916
rect 11888 36839 11940 36848
rect 11888 36805 11897 36839
rect 11897 36805 11931 36839
rect 11931 36805 11940 36839
rect 11888 36796 11940 36805
rect 13176 36796 13228 36848
rect 13452 36771 13504 36780
rect 13452 36737 13461 36771
rect 13461 36737 13495 36771
rect 13495 36737 13504 36771
rect 13452 36728 13504 36737
rect 13544 36728 13596 36780
rect 13912 36796 13964 36848
rect 16856 36864 16908 36916
rect 20536 36864 20588 36916
rect 20720 36907 20772 36916
rect 20720 36873 20729 36907
rect 20729 36873 20763 36907
rect 20763 36873 20772 36907
rect 20720 36864 20772 36873
rect 15384 36839 15436 36848
rect 14096 36771 14148 36780
rect 14096 36737 14105 36771
rect 14105 36737 14139 36771
rect 14139 36737 14148 36771
rect 14096 36728 14148 36737
rect 15384 36805 15393 36839
rect 15393 36805 15427 36839
rect 15427 36805 15436 36839
rect 15384 36796 15436 36805
rect 15108 36771 15160 36780
rect 15108 36737 15117 36771
rect 15117 36737 15151 36771
rect 15151 36737 15160 36771
rect 15108 36728 15160 36737
rect 17960 36796 18012 36848
rect 18696 36796 18748 36848
rect 20628 36796 20680 36848
rect 18512 36771 18564 36780
rect 18512 36737 18521 36771
rect 18521 36737 18555 36771
rect 18555 36737 18564 36771
rect 18512 36728 18564 36737
rect 18604 36771 18656 36780
rect 18604 36737 18613 36771
rect 18613 36737 18647 36771
rect 18647 36737 18656 36771
rect 18880 36771 18932 36780
rect 18604 36728 18656 36737
rect 18880 36737 18889 36771
rect 18889 36737 18923 36771
rect 18923 36737 18932 36771
rect 18880 36728 18932 36737
rect 19340 36728 19392 36780
rect 19708 36771 19760 36780
rect 19708 36737 19717 36771
rect 19717 36737 19751 36771
rect 19751 36737 19760 36771
rect 19708 36728 19760 36737
rect 19892 36771 19944 36780
rect 19892 36737 19901 36771
rect 19901 36737 19935 36771
rect 19935 36737 19944 36771
rect 19892 36728 19944 36737
rect 20536 36771 20588 36780
rect 18696 36703 18748 36712
rect 12532 36592 12584 36644
rect 15292 36592 15344 36644
rect 18696 36669 18705 36703
rect 18705 36669 18739 36703
rect 18739 36669 18748 36703
rect 18696 36660 18748 36669
rect 20536 36737 20545 36771
rect 20545 36737 20579 36771
rect 20579 36737 20588 36771
rect 20536 36728 20588 36737
rect 20628 36660 20680 36712
rect 22100 36864 22152 36916
rect 22652 36864 22704 36916
rect 23848 36864 23900 36916
rect 24676 36864 24728 36916
rect 26240 36864 26292 36916
rect 28264 36907 28316 36916
rect 28264 36873 28273 36907
rect 28273 36873 28307 36907
rect 28307 36873 28316 36907
rect 28264 36864 28316 36873
rect 28632 36864 28684 36916
rect 33048 36864 33100 36916
rect 37280 36864 37332 36916
rect 38108 36864 38160 36916
rect 40224 36907 40276 36916
rect 19340 36592 19392 36644
rect 19708 36592 19760 36644
rect 20260 36592 20312 36644
rect 20536 36592 20588 36644
rect 22468 36796 22520 36848
rect 23940 36796 23992 36848
rect 24768 36796 24820 36848
rect 25136 36839 25188 36848
rect 25136 36805 25145 36839
rect 25145 36805 25179 36839
rect 25179 36805 25188 36839
rect 25136 36796 25188 36805
rect 25228 36796 25280 36848
rect 25872 36796 25924 36848
rect 29828 36839 29880 36848
rect 29828 36805 29837 36839
rect 29837 36805 29871 36839
rect 29871 36805 29880 36839
rect 29828 36796 29880 36805
rect 31116 36796 31168 36848
rect 32772 36839 32824 36848
rect 23388 36771 23440 36780
rect 23388 36737 23397 36771
rect 23397 36737 23431 36771
rect 23431 36737 23440 36771
rect 23388 36728 23440 36737
rect 24124 36728 24176 36780
rect 24584 36728 24636 36780
rect 27804 36728 27856 36780
rect 28448 36771 28500 36780
rect 28448 36737 28457 36771
rect 28457 36737 28491 36771
rect 28491 36737 28500 36771
rect 28448 36728 28500 36737
rect 28540 36728 28592 36780
rect 28724 36771 28776 36780
rect 28724 36737 28733 36771
rect 28733 36737 28767 36771
rect 28767 36737 28776 36771
rect 28724 36728 28776 36737
rect 29552 36771 29604 36780
rect 22284 36703 22336 36712
rect 22284 36669 22293 36703
rect 22293 36669 22327 36703
rect 22327 36669 22336 36703
rect 22284 36660 22336 36669
rect 22376 36703 22428 36712
rect 22376 36669 22385 36703
rect 22385 36669 22419 36703
rect 22419 36669 22428 36703
rect 22376 36660 22428 36669
rect 22836 36660 22888 36712
rect 23020 36660 23072 36712
rect 23572 36660 23624 36712
rect 27528 36660 27580 36712
rect 29552 36737 29561 36771
rect 29561 36737 29595 36771
rect 29595 36737 29604 36771
rect 29552 36728 29604 36737
rect 30104 36728 30156 36780
rect 30380 36771 30432 36780
rect 30380 36737 30389 36771
rect 30389 36737 30423 36771
rect 30423 36737 30432 36771
rect 30380 36728 30432 36737
rect 30564 36771 30616 36780
rect 30564 36737 30573 36771
rect 30573 36737 30607 36771
rect 30607 36737 30616 36771
rect 30564 36728 30616 36737
rect 25136 36592 25188 36644
rect 26148 36592 26200 36644
rect 15844 36524 15896 36576
rect 16120 36567 16172 36576
rect 16120 36533 16129 36567
rect 16129 36533 16163 36567
rect 16163 36533 16172 36567
rect 16120 36524 16172 36533
rect 16948 36567 17000 36576
rect 16948 36533 16957 36567
rect 16957 36533 16991 36567
rect 16991 36533 17000 36567
rect 16948 36524 17000 36533
rect 20076 36524 20128 36576
rect 25320 36567 25372 36576
rect 25320 36533 25329 36567
rect 25329 36533 25363 36567
rect 25363 36533 25372 36567
rect 25320 36524 25372 36533
rect 25688 36524 25740 36576
rect 25964 36524 26016 36576
rect 28448 36592 28500 36644
rect 31116 36660 31168 36712
rect 31300 36771 31352 36780
rect 31300 36737 31309 36771
rect 31309 36737 31343 36771
rect 31343 36737 31352 36771
rect 32772 36805 32781 36839
rect 32781 36805 32815 36839
rect 32815 36805 32824 36839
rect 32772 36796 32824 36805
rect 33508 36796 33560 36848
rect 32496 36771 32548 36780
rect 31300 36728 31352 36737
rect 32496 36737 32505 36771
rect 32505 36737 32539 36771
rect 32539 36737 32548 36771
rect 32496 36728 32548 36737
rect 31484 36660 31536 36712
rect 32312 36660 32364 36712
rect 29644 36592 29696 36644
rect 28172 36524 28224 36576
rect 29000 36524 29052 36576
rect 30564 36567 30616 36576
rect 30564 36533 30573 36567
rect 30573 36533 30607 36567
rect 30607 36533 30616 36567
rect 30564 36524 30616 36533
rect 32404 36592 32456 36644
rect 32956 36771 33008 36780
rect 32956 36737 32970 36771
rect 32970 36737 33004 36771
rect 33004 36737 33008 36771
rect 32956 36728 33008 36737
rect 33600 36728 33652 36780
rect 35532 36796 35584 36848
rect 34520 36771 34572 36780
rect 34520 36737 34529 36771
rect 34529 36737 34563 36771
rect 34563 36737 34572 36771
rect 34520 36728 34572 36737
rect 34704 36592 34756 36644
rect 31300 36567 31352 36576
rect 31300 36533 31309 36567
rect 31309 36533 31343 36567
rect 31343 36533 31352 36567
rect 31300 36524 31352 36533
rect 31944 36524 31996 36576
rect 32496 36524 32548 36576
rect 33324 36524 33376 36576
rect 33876 36524 33928 36576
rect 34244 36524 34296 36576
rect 34428 36524 34480 36576
rect 35440 36728 35492 36780
rect 35808 36771 35860 36780
rect 35808 36737 35817 36771
rect 35817 36737 35851 36771
rect 35851 36737 35860 36771
rect 35808 36728 35860 36737
rect 35992 36728 36044 36780
rect 38476 36796 38528 36848
rect 40224 36873 40233 36907
rect 40233 36873 40267 36907
rect 40267 36873 40276 36907
rect 40224 36864 40276 36873
rect 42616 36864 42668 36916
rect 43352 36864 43404 36916
rect 38384 36771 38436 36780
rect 36636 36703 36688 36712
rect 36636 36669 36645 36703
rect 36645 36669 36679 36703
rect 36679 36669 36688 36703
rect 38384 36737 38393 36771
rect 38393 36737 38427 36771
rect 38427 36737 38436 36771
rect 38384 36728 38436 36737
rect 38568 36728 38620 36780
rect 39488 36728 39540 36780
rect 40408 36796 40460 36848
rect 40868 36796 40920 36848
rect 41236 36771 41288 36780
rect 41236 36737 41245 36771
rect 41245 36737 41279 36771
rect 41279 36737 41288 36771
rect 41236 36728 41288 36737
rect 44180 36796 44232 36848
rect 47584 36839 47636 36848
rect 47584 36805 47593 36839
rect 47593 36805 47627 36839
rect 47627 36805 47636 36839
rect 47584 36796 47636 36805
rect 47768 36771 47820 36780
rect 36636 36660 36688 36669
rect 39948 36660 40000 36712
rect 37280 36635 37332 36644
rect 37280 36601 37289 36635
rect 37289 36601 37323 36635
rect 37323 36601 37332 36635
rect 37280 36592 37332 36601
rect 38660 36592 38712 36644
rect 40316 36592 40368 36644
rect 35348 36524 35400 36576
rect 38200 36567 38252 36576
rect 38200 36533 38209 36567
rect 38209 36533 38243 36567
rect 38243 36533 38252 36567
rect 38200 36524 38252 36533
rect 39120 36524 39172 36576
rect 39856 36567 39908 36576
rect 39856 36533 39865 36567
rect 39865 36533 39899 36567
rect 39899 36533 39908 36567
rect 47768 36737 47777 36771
rect 47777 36737 47811 36771
rect 47811 36737 47820 36771
rect 47768 36728 47820 36737
rect 47952 36771 48004 36780
rect 47952 36737 47961 36771
rect 47961 36737 47995 36771
rect 47995 36737 48004 36771
rect 47952 36728 48004 36737
rect 47216 36592 47268 36644
rect 47768 36592 47820 36644
rect 39856 36524 39908 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 11888 36363 11940 36372
rect 11888 36329 11897 36363
rect 11897 36329 11931 36363
rect 11931 36329 11940 36363
rect 11888 36320 11940 36329
rect 15936 36363 15988 36372
rect 15936 36329 15945 36363
rect 15945 36329 15979 36363
rect 15979 36329 15988 36363
rect 15936 36320 15988 36329
rect 18236 36363 18288 36372
rect 18236 36329 18245 36363
rect 18245 36329 18279 36363
rect 18279 36329 18288 36363
rect 18236 36320 18288 36329
rect 18512 36320 18564 36372
rect 19340 36363 19392 36372
rect 19340 36329 19349 36363
rect 19349 36329 19383 36363
rect 19383 36329 19392 36363
rect 19340 36320 19392 36329
rect 20444 36320 20496 36372
rect 22744 36320 22796 36372
rect 25412 36320 25464 36372
rect 26792 36320 26844 36372
rect 27528 36363 27580 36372
rect 27528 36329 27537 36363
rect 27537 36329 27571 36363
rect 27571 36329 27580 36363
rect 27528 36320 27580 36329
rect 27620 36320 27672 36372
rect 30380 36320 30432 36372
rect 30840 36320 30892 36372
rect 31392 36320 31444 36372
rect 32772 36320 32824 36372
rect 34612 36320 34664 36372
rect 35624 36363 35676 36372
rect 35624 36329 35633 36363
rect 35633 36329 35667 36363
rect 35667 36329 35676 36363
rect 35624 36320 35676 36329
rect 38384 36320 38436 36372
rect 21732 36252 21784 36304
rect 15568 36227 15620 36236
rect 15568 36193 15577 36227
rect 15577 36193 15611 36227
rect 15611 36193 15620 36227
rect 15568 36184 15620 36193
rect 17224 36227 17276 36236
rect 17224 36193 17233 36227
rect 17233 36193 17267 36227
rect 17267 36193 17276 36227
rect 17224 36184 17276 36193
rect 17776 36184 17828 36236
rect 12992 36159 13044 36168
rect 12992 36125 13001 36159
rect 13001 36125 13035 36159
rect 13035 36125 13044 36159
rect 15660 36159 15712 36168
rect 12992 36116 13044 36125
rect 11888 36048 11940 36100
rect 14096 36048 14148 36100
rect 1492 36023 1544 36032
rect 1492 35989 1501 36023
rect 1501 35989 1535 36023
rect 1535 35989 1544 36023
rect 1492 35980 1544 35989
rect 13728 35980 13780 36032
rect 15660 36125 15669 36159
rect 15669 36125 15703 36159
rect 15703 36125 15712 36159
rect 15660 36116 15712 36125
rect 16856 36116 16908 36168
rect 17500 36116 17552 36168
rect 17684 36159 17736 36168
rect 17684 36125 17693 36159
rect 17693 36125 17727 36159
rect 17727 36125 17736 36159
rect 19984 36184 20036 36236
rect 21456 36184 21508 36236
rect 17684 36116 17736 36125
rect 19432 36159 19484 36168
rect 16028 36048 16080 36100
rect 16580 36048 16632 36100
rect 19432 36125 19441 36159
rect 19441 36125 19475 36159
rect 19475 36125 19484 36159
rect 19432 36116 19484 36125
rect 20444 36159 20496 36168
rect 20444 36125 20453 36159
rect 20453 36125 20487 36159
rect 20487 36125 20496 36159
rect 20444 36116 20496 36125
rect 20628 36159 20680 36168
rect 20628 36125 20637 36159
rect 20637 36125 20671 36159
rect 20671 36125 20680 36159
rect 20628 36116 20680 36125
rect 22836 36227 22888 36236
rect 22836 36193 22845 36227
rect 22845 36193 22879 36227
rect 22879 36193 22888 36227
rect 22836 36184 22888 36193
rect 22744 36159 22796 36168
rect 18328 36048 18380 36100
rect 18696 36048 18748 36100
rect 22744 36125 22753 36159
rect 22753 36125 22787 36159
rect 22787 36125 22796 36159
rect 22744 36116 22796 36125
rect 25228 36116 25280 36168
rect 28632 36252 28684 36304
rect 28908 36252 28960 36304
rect 28448 36184 28500 36236
rect 31300 36252 31352 36304
rect 26148 36116 26200 36168
rect 27712 36159 27764 36168
rect 27712 36125 27721 36159
rect 27721 36125 27755 36159
rect 27755 36125 27764 36159
rect 27712 36116 27764 36125
rect 27988 36116 28040 36168
rect 28172 36116 28224 36168
rect 25320 36091 25372 36100
rect 16672 35980 16724 36032
rect 17960 35980 18012 36032
rect 18512 35980 18564 36032
rect 19156 35980 19208 36032
rect 21456 36023 21508 36032
rect 21456 35989 21465 36023
rect 21465 35989 21499 36023
rect 21499 35989 21508 36023
rect 21456 35980 21508 35989
rect 25320 36057 25329 36091
rect 25329 36057 25363 36091
rect 25363 36057 25372 36091
rect 25320 36048 25372 36057
rect 22468 35980 22520 36032
rect 22744 35980 22796 36032
rect 23480 35980 23532 36032
rect 23664 35980 23716 36032
rect 24308 35980 24360 36032
rect 24768 35980 24820 36032
rect 25412 35980 25464 36032
rect 25780 35980 25832 36032
rect 26056 35980 26108 36032
rect 28724 36116 28776 36168
rect 31852 36184 31904 36236
rect 34704 36184 34756 36236
rect 34796 36227 34848 36236
rect 34796 36193 34805 36227
rect 34805 36193 34839 36227
rect 34839 36193 34848 36227
rect 34796 36184 34848 36193
rect 30564 36159 30616 36168
rect 30564 36125 30573 36159
rect 30573 36125 30607 36159
rect 30607 36125 30616 36159
rect 30564 36116 30616 36125
rect 31484 36116 31536 36168
rect 31944 36159 31996 36168
rect 31944 36125 31953 36159
rect 31953 36125 31987 36159
rect 31987 36125 31996 36159
rect 31944 36116 31996 36125
rect 33048 36159 33100 36168
rect 33048 36125 33057 36159
rect 33057 36125 33091 36159
rect 33091 36125 33100 36159
rect 33048 36116 33100 36125
rect 33692 36159 33744 36168
rect 33692 36125 33701 36159
rect 33701 36125 33735 36159
rect 33735 36125 33744 36159
rect 33692 36116 33744 36125
rect 33876 36159 33928 36168
rect 33876 36125 33885 36159
rect 33885 36125 33919 36159
rect 33919 36125 33928 36159
rect 33876 36116 33928 36125
rect 38660 36252 38712 36304
rect 36268 36159 36320 36168
rect 36268 36125 36277 36159
rect 36277 36125 36311 36159
rect 36311 36125 36320 36159
rect 36268 36116 36320 36125
rect 36636 36116 36688 36168
rect 37004 36159 37056 36168
rect 37004 36125 37013 36159
rect 37013 36125 37047 36159
rect 37047 36125 37056 36159
rect 37004 36116 37056 36125
rect 37464 36116 37516 36168
rect 37740 36116 37792 36168
rect 38200 36159 38252 36168
rect 31300 36048 31352 36100
rect 35808 36048 35860 36100
rect 31760 35980 31812 36032
rect 32220 35980 32272 36032
rect 36452 36048 36504 36100
rect 38200 36125 38209 36159
rect 38209 36125 38243 36159
rect 38243 36125 38252 36159
rect 38200 36116 38252 36125
rect 40040 36252 40092 36304
rect 40408 36320 40460 36372
rect 41880 36320 41932 36372
rect 42616 36320 42668 36372
rect 47216 36363 47268 36372
rect 47216 36329 47225 36363
rect 47225 36329 47259 36363
rect 47259 36329 47268 36363
rect 47216 36320 47268 36329
rect 39212 36116 39264 36168
rect 39856 36116 39908 36168
rect 40132 36116 40184 36168
rect 40868 36116 40920 36168
rect 41236 36137 41288 36146
rect 41236 36103 41245 36137
rect 41245 36103 41279 36137
rect 41279 36103 41288 36137
rect 41236 36094 41288 36103
rect 39856 36023 39908 36032
rect 39856 35989 39865 36023
rect 39865 35989 39899 36023
rect 39899 35989 39908 36023
rect 39856 35980 39908 35989
rect 40316 35980 40368 36032
rect 47860 36091 47912 36100
rect 47860 36057 47869 36091
rect 47869 36057 47903 36091
rect 47903 36057 47912 36091
rect 47860 36048 47912 36057
rect 48044 36091 48096 36100
rect 48044 36057 48053 36091
rect 48053 36057 48087 36091
rect 48087 36057 48096 36091
rect 48044 36048 48096 36057
rect 42984 36023 43036 36032
rect 42984 35989 42993 36023
rect 42993 35989 43027 36023
rect 43027 35989 43036 36023
rect 42984 35980 43036 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 10232 35776 10284 35828
rect 12716 35819 12768 35828
rect 12716 35785 12725 35819
rect 12725 35785 12759 35819
rect 12759 35785 12768 35819
rect 12716 35776 12768 35785
rect 13268 35819 13320 35828
rect 13268 35785 13277 35819
rect 13277 35785 13311 35819
rect 13311 35785 13320 35819
rect 13268 35776 13320 35785
rect 12992 35708 13044 35760
rect 17500 35776 17552 35828
rect 18236 35708 18288 35760
rect 19800 35776 19852 35828
rect 21916 35776 21968 35828
rect 24032 35819 24084 35828
rect 24032 35785 24041 35819
rect 24041 35785 24075 35819
rect 24075 35785 24084 35819
rect 24032 35776 24084 35785
rect 24676 35776 24728 35828
rect 25412 35776 25464 35828
rect 25504 35776 25556 35828
rect 30012 35776 30064 35828
rect 30656 35776 30708 35828
rect 31300 35776 31352 35828
rect 33140 35776 33192 35828
rect 33416 35776 33468 35828
rect 33692 35776 33744 35828
rect 35532 35819 35584 35828
rect 35532 35785 35541 35819
rect 35541 35785 35575 35819
rect 35575 35785 35584 35819
rect 35532 35776 35584 35785
rect 36268 35776 36320 35828
rect 38200 35776 38252 35828
rect 38844 35776 38896 35828
rect 48044 35819 48096 35828
rect 24216 35708 24268 35760
rect 14280 35683 14332 35692
rect 14280 35649 14289 35683
rect 14289 35649 14323 35683
rect 14323 35649 14332 35683
rect 14280 35640 14332 35649
rect 15384 35683 15436 35692
rect 13820 35572 13872 35624
rect 15384 35649 15393 35683
rect 15393 35649 15427 35683
rect 15427 35649 15436 35683
rect 15384 35640 15436 35649
rect 16580 35640 16632 35692
rect 15476 35615 15528 35624
rect 15476 35581 15485 35615
rect 15485 35581 15519 35615
rect 15519 35581 15528 35615
rect 15476 35572 15528 35581
rect 16856 35683 16908 35692
rect 16856 35649 16865 35683
rect 16865 35649 16899 35683
rect 16899 35649 16908 35683
rect 16856 35640 16908 35649
rect 17224 35640 17276 35692
rect 18512 35640 18564 35692
rect 18972 35640 19024 35692
rect 19064 35683 19116 35692
rect 19064 35649 19073 35683
rect 19073 35649 19107 35683
rect 19107 35649 19116 35683
rect 19064 35640 19116 35649
rect 19432 35640 19484 35692
rect 19892 35683 19944 35692
rect 19892 35649 19901 35683
rect 19901 35649 19935 35683
rect 19935 35649 19944 35683
rect 19892 35640 19944 35649
rect 19984 35640 20036 35692
rect 20812 35683 20864 35692
rect 20812 35649 20821 35683
rect 20821 35649 20855 35683
rect 20855 35649 20864 35683
rect 20812 35640 20864 35649
rect 21456 35640 21508 35692
rect 22376 35640 22428 35692
rect 22560 35683 22612 35692
rect 22560 35649 22569 35683
rect 22569 35649 22603 35683
rect 22603 35649 22612 35683
rect 22560 35640 22612 35649
rect 25964 35708 26016 35760
rect 24676 35683 24728 35692
rect 24676 35649 24685 35683
rect 24685 35649 24719 35683
rect 24719 35649 24728 35683
rect 24676 35640 24728 35649
rect 17500 35572 17552 35624
rect 18420 35572 18472 35624
rect 18880 35615 18932 35624
rect 18880 35581 18889 35615
rect 18889 35581 18923 35615
rect 18923 35581 18932 35615
rect 18880 35572 18932 35581
rect 24952 35640 25004 35692
rect 13728 35504 13780 35556
rect 17960 35504 18012 35556
rect 9128 35436 9180 35488
rect 11888 35436 11940 35488
rect 14096 35436 14148 35488
rect 14464 35479 14516 35488
rect 14464 35445 14473 35479
rect 14473 35445 14507 35479
rect 14507 35445 14516 35479
rect 14464 35436 14516 35445
rect 23756 35504 23808 35556
rect 24400 35504 24452 35556
rect 25872 35683 25924 35692
rect 25872 35649 25882 35683
rect 25882 35649 25916 35683
rect 25916 35649 25924 35683
rect 26792 35708 26844 35760
rect 27160 35708 27212 35760
rect 30288 35708 30340 35760
rect 34060 35751 34112 35760
rect 34060 35717 34069 35751
rect 34069 35717 34103 35751
rect 34103 35717 34112 35751
rect 34060 35708 34112 35717
rect 25872 35640 25924 35649
rect 27620 35640 27672 35692
rect 29092 35640 29144 35692
rect 30104 35640 30156 35692
rect 26056 35615 26108 35624
rect 26056 35581 26065 35615
rect 26065 35581 26099 35615
rect 26099 35581 26108 35615
rect 26056 35572 26108 35581
rect 18328 35436 18380 35488
rect 22376 35436 22428 35488
rect 22744 35436 22796 35488
rect 23572 35436 23624 35488
rect 25136 35436 25188 35488
rect 27712 35572 27764 35624
rect 26976 35504 27028 35556
rect 29460 35572 29512 35624
rect 29828 35572 29880 35624
rect 30288 35572 30340 35624
rect 30840 35640 30892 35692
rect 31484 35640 31536 35692
rect 32220 35683 32272 35692
rect 32220 35649 32229 35683
rect 32229 35649 32263 35683
rect 32263 35649 32272 35683
rect 32220 35640 32272 35649
rect 32404 35683 32456 35692
rect 32404 35649 32413 35683
rect 32413 35649 32447 35683
rect 32447 35649 32456 35683
rect 32404 35640 32456 35649
rect 33508 35640 33560 35692
rect 34244 35640 34296 35692
rect 34428 35640 34480 35692
rect 30748 35615 30800 35624
rect 30748 35581 30757 35615
rect 30757 35581 30791 35615
rect 30791 35581 30800 35615
rect 30748 35572 30800 35581
rect 28816 35504 28868 35556
rect 27068 35479 27120 35488
rect 27068 35445 27077 35479
rect 27077 35445 27111 35479
rect 27111 35445 27120 35479
rect 27068 35436 27120 35445
rect 27252 35436 27304 35488
rect 29552 35479 29604 35488
rect 29552 35445 29561 35479
rect 29561 35445 29595 35479
rect 29595 35445 29604 35479
rect 29552 35436 29604 35445
rect 33600 35572 33652 35624
rect 36452 35640 36504 35692
rect 36544 35640 36596 35692
rect 37004 35640 37056 35692
rect 37464 35683 37516 35692
rect 37464 35649 37473 35683
rect 37473 35649 37507 35683
rect 37507 35649 37516 35683
rect 38292 35751 38344 35760
rect 48044 35785 48053 35819
rect 48053 35785 48087 35819
rect 48087 35785 48096 35819
rect 48044 35776 48096 35785
rect 38292 35717 38317 35751
rect 38317 35717 38344 35751
rect 38292 35708 38344 35717
rect 37464 35640 37516 35649
rect 38844 35640 38896 35692
rect 39028 35683 39080 35692
rect 39028 35649 39037 35683
rect 39037 35649 39071 35683
rect 39071 35649 39080 35683
rect 39028 35640 39080 35649
rect 40040 35640 40092 35692
rect 40316 35683 40368 35692
rect 40316 35649 40325 35683
rect 40325 35649 40359 35683
rect 40359 35649 40368 35683
rect 40316 35640 40368 35649
rect 39212 35547 39264 35556
rect 39212 35513 39221 35547
rect 39221 35513 39255 35547
rect 39255 35513 39264 35547
rect 39212 35504 39264 35513
rect 34796 35479 34848 35488
rect 34796 35445 34805 35479
rect 34805 35445 34839 35479
rect 34839 35445 34848 35479
rect 34796 35436 34848 35445
rect 39028 35436 39080 35488
rect 40132 35479 40184 35488
rect 40132 35445 40141 35479
rect 40141 35445 40175 35479
rect 40175 35445 40184 35479
rect 40132 35436 40184 35445
rect 41420 35479 41472 35488
rect 41420 35445 41429 35479
rect 41429 35445 41463 35479
rect 41463 35445 41472 35479
rect 41420 35436 41472 35445
rect 41512 35436 41564 35488
rect 42156 35436 42208 35488
rect 42984 35436 43036 35488
rect 43260 35436 43312 35488
rect 43536 35479 43588 35488
rect 43536 35445 43545 35479
rect 43545 35445 43579 35479
rect 43579 35445 43588 35479
rect 43536 35436 43588 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 10876 35232 10928 35284
rect 1952 34960 2004 35012
rect 12624 35096 12676 35148
rect 14096 35164 14148 35216
rect 15568 35232 15620 35284
rect 18236 35232 18288 35284
rect 18328 35275 18380 35284
rect 18328 35241 18337 35275
rect 18337 35241 18371 35275
rect 18371 35241 18380 35275
rect 18328 35232 18380 35241
rect 18880 35232 18932 35284
rect 19432 35232 19484 35284
rect 19892 35232 19944 35284
rect 20812 35232 20864 35284
rect 22284 35232 22336 35284
rect 24768 35232 24820 35284
rect 26976 35232 27028 35284
rect 28172 35232 28224 35284
rect 28264 35232 28316 35284
rect 11520 35028 11572 35080
rect 11980 35071 12032 35080
rect 11980 35037 11989 35071
rect 11989 35037 12023 35071
rect 12023 35037 12032 35071
rect 11980 35028 12032 35037
rect 12440 35028 12492 35080
rect 12808 35071 12860 35080
rect 12808 35037 12817 35071
rect 12817 35037 12851 35071
rect 12851 35037 12860 35071
rect 12808 35028 12860 35037
rect 13268 35003 13320 35012
rect 13268 34969 13277 35003
rect 13277 34969 13311 35003
rect 13311 34969 13320 35003
rect 13268 34960 13320 34969
rect 13544 35071 13596 35080
rect 13544 35037 13553 35071
rect 13553 35037 13587 35071
rect 13587 35037 13596 35071
rect 15844 35096 15896 35148
rect 13544 35028 13596 35037
rect 12716 34892 12768 34944
rect 15568 35071 15620 35080
rect 15568 35037 15577 35071
rect 15577 35037 15611 35071
rect 15611 35037 15620 35071
rect 15568 35028 15620 35037
rect 17040 35096 17092 35148
rect 16672 35028 16724 35080
rect 17132 35028 17184 35080
rect 18144 35028 18196 35080
rect 19984 35096 20036 35148
rect 22560 35164 22612 35216
rect 21088 35096 21140 35148
rect 21456 35096 21508 35148
rect 22744 35139 22796 35148
rect 22744 35105 22753 35139
rect 22753 35105 22787 35139
rect 22787 35105 22796 35139
rect 22744 35096 22796 35105
rect 23020 35139 23072 35148
rect 23020 35105 23029 35139
rect 23029 35105 23063 35139
rect 23063 35105 23072 35139
rect 23020 35096 23072 35105
rect 18512 35071 18564 35080
rect 18512 35037 18521 35071
rect 18521 35037 18555 35071
rect 18555 35037 18564 35071
rect 18512 35028 18564 35037
rect 19800 35071 19852 35080
rect 19800 35037 19809 35071
rect 19809 35037 19843 35071
rect 19843 35037 19852 35071
rect 19800 35028 19852 35037
rect 20720 35071 20772 35080
rect 20720 35037 20729 35071
rect 20729 35037 20763 35071
rect 20763 35037 20772 35071
rect 20720 35028 20772 35037
rect 21548 35071 21600 35080
rect 21548 35037 21557 35071
rect 21557 35037 21591 35071
rect 21591 35037 21600 35071
rect 21548 35028 21600 35037
rect 21640 35071 21692 35080
rect 21640 35037 21649 35071
rect 21649 35037 21683 35071
rect 21683 35037 21692 35071
rect 21640 35028 21692 35037
rect 19432 34960 19484 35012
rect 20076 34960 20128 35012
rect 22560 35071 22612 35080
rect 22560 35037 22569 35071
rect 22569 35037 22603 35071
rect 22603 35037 22612 35071
rect 22560 35028 22612 35037
rect 23112 35071 23164 35080
rect 23112 35037 23121 35071
rect 23121 35037 23155 35071
rect 23155 35037 23164 35071
rect 23112 35028 23164 35037
rect 24492 35071 24544 35080
rect 24492 35037 24501 35071
rect 24501 35037 24535 35071
rect 24535 35037 24544 35071
rect 24492 35028 24544 35037
rect 24952 35028 25004 35080
rect 25136 35096 25188 35148
rect 27712 35164 27764 35216
rect 30288 35232 30340 35284
rect 30840 35232 30892 35284
rect 31300 35232 31352 35284
rect 32036 35232 32088 35284
rect 33232 35275 33284 35284
rect 33232 35241 33241 35275
rect 33241 35241 33275 35275
rect 33275 35241 33284 35275
rect 33232 35232 33284 35241
rect 33508 35232 33560 35284
rect 26148 35071 26200 35080
rect 14556 34935 14608 34944
rect 14556 34901 14565 34935
rect 14565 34901 14599 34935
rect 14599 34901 14608 34935
rect 14556 34892 14608 34901
rect 15384 34892 15436 34944
rect 15936 34892 15988 34944
rect 18052 34892 18104 34944
rect 18788 34892 18840 34944
rect 19340 34892 19392 34944
rect 24860 34960 24912 35012
rect 25872 34960 25924 35012
rect 26148 35037 26157 35071
rect 26157 35037 26191 35071
rect 26191 35037 26200 35071
rect 26148 35028 26200 35037
rect 26240 35028 26292 35080
rect 26792 34960 26844 35012
rect 27068 35028 27120 35080
rect 27252 35071 27304 35080
rect 27252 35037 27261 35071
rect 27261 35037 27295 35071
rect 27295 35037 27304 35071
rect 27252 35028 27304 35037
rect 26056 34892 26108 34944
rect 27252 34892 27304 34944
rect 27344 34892 27396 34944
rect 27620 34960 27672 35012
rect 28264 35028 28316 35080
rect 31576 35164 31628 35216
rect 33600 35164 33652 35216
rect 36544 35207 36596 35216
rect 30840 35096 30892 35148
rect 29920 35028 29972 35080
rect 30564 35071 30616 35080
rect 30564 35037 30568 35071
rect 30568 35037 30602 35071
rect 30602 35037 30616 35071
rect 30564 35028 30616 35037
rect 31944 35096 31996 35148
rect 34152 35096 34204 35148
rect 34704 35139 34756 35148
rect 34704 35105 34713 35139
rect 34713 35105 34747 35139
rect 34747 35105 34756 35139
rect 34704 35096 34756 35105
rect 32036 35028 32088 35080
rect 33416 35071 33468 35080
rect 33416 35037 33425 35071
rect 33425 35037 33459 35071
rect 33459 35037 33468 35071
rect 33416 35028 33468 35037
rect 33784 35071 33836 35080
rect 30472 34960 30524 35012
rect 28264 34935 28316 34944
rect 28264 34901 28273 34935
rect 28273 34901 28307 34935
rect 28307 34901 28316 34935
rect 28264 34892 28316 34901
rect 28908 34892 28960 34944
rect 30748 35003 30800 35012
rect 30748 34969 30757 35003
rect 30757 34969 30791 35003
rect 30791 34969 30800 35003
rect 30748 34960 30800 34969
rect 31944 34960 31996 35012
rect 32128 34960 32180 35012
rect 32404 35003 32456 35012
rect 32404 34969 32413 35003
rect 32413 34969 32447 35003
rect 32447 34969 32456 35003
rect 32404 34960 32456 34969
rect 33784 35037 33793 35071
rect 33793 35037 33827 35071
rect 33827 35037 33836 35071
rect 33784 35028 33836 35037
rect 34888 35028 34940 35080
rect 36544 35173 36553 35207
rect 36553 35173 36587 35207
rect 36587 35173 36596 35207
rect 36544 35164 36596 35173
rect 38108 35164 38160 35216
rect 38568 35164 38620 35216
rect 36268 35139 36320 35148
rect 36268 35105 36277 35139
rect 36277 35105 36311 35139
rect 36311 35105 36320 35139
rect 36268 35096 36320 35105
rect 37372 35028 37424 35080
rect 37924 35071 37976 35080
rect 37924 35037 37933 35071
rect 37933 35037 37967 35071
rect 37967 35037 37976 35071
rect 37924 35028 37976 35037
rect 38200 35028 38252 35080
rect 41512 35275 41564 35284
rect 41512 35241 41521 35275
rect 41521 35241 41555 35275
rect 41555 35241 41564 35275
rect 41512 35232 41564 35241
rect 38844 35164 38896 35216
rect 43536 35232 43588 35284
rect 40132 35139 40184 35148
rect 40132 35105 40141 35139
rect 40141 35105 40175 35139
rect 40175 35105 40184 35139
rect 40132 35096 40184 35105
rect 39764 35028 39816 35080
rect 40868 35028 40920 35080
rect 39120 34960 39172 35012
rect 39948 34960 40000 35012
rect 41420 35028 41472 35080
rect 41972 35028 42024 35080
rect 41512 34960 41564 35012
rect 41880 34960 41932 35012
rect 31760 34892 31812 34944
rect 34520 34892 34572 34944
rect 37004 34935 37056 34944
rect 37004 34901 37013 34935
rect 37013 34901 37047 34935
rect 37047 34901 37056 34935
rect 37004 34892 37056 34901
rect 38108 34892 38160 34944
rect 39304 34935 39356 34944
rect 39304 34901 39313 34935
rect 39313 34901 39347 34935
rect 39347 34901 39356 34935
rect 39304 34892 39356 34901
rect 39764 34892 39816 34944
rect 41696 34892 41748 34944
rect 43076 34935 43128 34944
rect 43076 34901 43085 34935
rect 43085 34901 43119 34935
rect 43119 34901 43128 34935
rect 43076 34892 43128 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 1952 34731 2004 34740
rect 1952 34697 1961 34731
rect 1961 34697 1995 34731
rect 1995 34697 2004 34731
rect 1952 34688 2004 34697
rect 9128 34731 9180 34740
rect 9128 34697 9137 34731
rect 9137 34697 9171 34731
rect 9171 34697 9180 34731
rect 9128 34688 9180 34697
rect 10232 34731 10284 34740
rect 10232 34697 10241 34731
rect 10241 34697 10275 34731
rect 10275 34697 10284 34731
rect 10232 34688 10284 34697
rect 11980 34688 12032 34740
rect 12072 34688 12124 34740
rect 12808 34688 12860 34740
rect 13268 34688 13320 34740
rect 14556 34688 14608 34740
rect 15660 34688 15712 34740
rect 16856 34688 16908 34740
rect 19340 34688 19392 34740
rect 19984 34688 20036 34740
rect 21640 34688 21692 34740
rect 23112 34731 23164 34740
rect 23112 34697 23121 34731
rect 23121 34697 23155 34731
rect 23155 34697 23164 34731
rect 23112 34688 23164 34697
rect 24676 34688 24728 34740
rect 25044 34688 25096 34740
rect 26148 34688 26200 34740
rect 1584 34552 1636 34604
rect 12624 34620 12676 34672
rect 10324 34484 10376 34536
rect 12440 34595 12492 34604
rect 12440 34561 12449 34595
rect 12449 34561 12483 34595
rect 12483 34561 12492 34595
rect 12716 34595 12768 34604
rect 12440 34552 12492 34561
rect 12716 34561 12725 34595
rect 12725 34561 12759 34595
rect 12759 34561 12768 34595
rect 12716 34552 12768 34561
rect 13820 34595 13872 34604
rect 13820 34561 13829 34595
rect 13829 34561 13863 34595
rect 13863 34561 13872 34595
rect 13820 34552 13872 34561
rect 10232 34416 10284 34468
rect 14280 34484 14332 34536
rect 14464 34552 14516 34604
rect 14740 34595 14792 34604
rect 14740 34561 14749 34595
rect 14749 34561 14783 34595
rect 14783 34561 14792 34595
rect 14740 34552 14792 34561
rect 16580 34620 16632 34672
rect 15292 34484 15344 34536
rect 15844 34552 15896 34604
rect 17960 34620 18012 34672
rect 18788 34663 18840 34672
rect 18788 34629 18797 34663
rect 18797 34629 18831 34663
rect 18831 34629 18840 34663
rect 18788 34620 18840 34629
rect 15384 34459 15436 34468
rect 15384 34425 15393 34459
rect 15393 34425 15427 34459
rect 15427 34425 15436 34459
rect 15384 34416 15436 34425
rect 16672 34484 16724 34536
rect 16764 34527 16816 34536
rect 16764 34493 16773 34527
rect 16773 34493 16807 34527
rect 16807 34493 16816 34527
rect 21272 34620 21324 34672
rect 23480 34663 23532 34672
rect 23480 34629 23489 34663
rect 23489 34629 23523 34663
rect 23523 34629 23532 34663
rect 23480 34620 23532 34629
rect 19248 34595 19300 34604
rect 19248 34561 19257 34595
rect 19257 34561 19291 34595
rect 19291 34561 19300 34595
rect 19248 34552 19300 34561
rect 19340 34595 19392 34604
rect 19340 34561 19349 34595
rect 19349 34561 19383 34595
rect 19383 34561 19392 34595
rect 19340 34552 19392 34561
rect 16764 34484 16816 34493
rect 19432 34484 19484 34536
rect 21088 34552 21140 34604
rect 22376 34552 22428 34604
rect 20720 34484 20772 34536
rect 22192 34527 22244 34536
rect 22192 34493 22201 34527
rect 22201 34493 22235 34527
rect 22235 34493 22244 34527
rect 22192 34484 22244 34493
rect 17316 34416 17368 34468
rect 23664 34595 23716 34604
rect 23664 34561 23672 34595
rect 23672 34561 23706 34595
rect 23706 34561 23716 34595
rect 23664 34552 23716 34561
rect 24032 34552 24084 34604
rect 24216 34595 24268 34604
rect 24216 34561 24225 34595
rect 24225 34561 24259 34595
rect 24259 34561 24268 34595
rect 24216 34552 24268 34561
rect 24768 34552 24820 34604
rect 25228 34595 25280 34604
rect 23480 34484 23532 34536
rect 25228 34561 25237 34595
rect 25237 34561 25271 34595
rect 25271 34561 25280 34595
rect 25228 34552 25280 34561
rect 25780 34595 25832 34604
rect 25780 34561 25789 34595
rect 25789 34561 25823 34595
rect 25823 34561 25832 34595
rect 25780 34552 25832 34561
rect 26056 34595 26108 34604
rect 26056 34561 26065 34595
rect 26065 34561 26099 34595
rect 26099 34561 26108 34595
rect 26056 34552 26108 34561
rect 26240 34552 26292 34604
rect 27160 34595 27212 34604
rect 27160 34561 27169 34595
rect 27169 34561 27203 34595
rect 27203 34561 27212 34595
rect 27160 34552 27212 34561
rect 30748 34688 30800 34740
rect 31484 34731 31536 34740
rect 31484 34697 31493 34731
rect 31493 34697 31527 34731
rect 31527 34697 31536 34731
rect 31484 34688 31536 34697
rect 31576 34688 31628 34740
rect 32220 34731 32272 34740
rect 32220 34697 32229 34731
rect 32229 34697 32263 34731
rect 32263 34697 32272 34731
rect 32220 34688 32272 34697
rect 33416 34731 33468 34740
rect 33416 34697 33425 34731
rect 33425 34697 33459 34731
rect 33459 34697 33468 34731
rect 33416 34688 33468 34697
rect 34152 34731 34204 34740
rect 34152 34697 34161 34731
rect 34161 34697 34195 34731
rect 34195 34697 34204 34731
rect 34152 34688 34204 34697
rect 36268 34688 36320 34740
rect 38292 34688 38344 34740
rect 38660 34688 38712 34740
rect 39028 34688 39080 34740
rect 39948 34688 40000 34740
rect 41236 34688 41288 34740
rect 27620 34620 27672 34672
rect 28264 34620 28316 34672
rect 25412 34484 25464 34536
rect 25688 34484 25740 34536
rect 27068 34527 27120 34536
rect 27068 34493 27077 34527
rect 27077 34493 27111 34527
rect 27111 34493 27120 34527
rect 27068 34484 27120 34493
rect 27252 34527 27304 34536
rect 27252 34493 27261 34527
rect 27261 34493 27295 34527
rect 27295 34493 27304 34527
rect 28172 34552 28224 34604
rect 28724 34552 28776 34604
rect 28908 34595 28960 34604
rect 28908 34561 28917 34595
rect 28917 34561 28951 34595
rect 28951 34561 28960 34595
rect 28908 34552 28960 34561
rect 27252 34484 27304 34493
rect 27620 34484 27672 34536
rect 28816 34527 28868 34536
rect 28816 34493 28825 34527
rect 28825 34493 28859 34527
rect 28859 34493 28868 34527
rect 28816 34484 28868 34493
rect 31300 34620 31352 34672
rect 29920 34595 29972 34604
rect 29920 34561 29929 34595
rect 29929 34561 29963 34595
rect 29963 34561 29972 34595
rect 30748 34595 30800 34604
rect 29920 34552 29972 34561
rect 30748 34561 30757 34595
rect 30757 34561 30791 34595
rect 30791 34561 30800 34595
rect 30748 34552 30800 34561
rect 31760 34552 31812 34604
rect 33324 34595 33376 34604
rect 33324 34561 33333 34595
rect 33333 34561 33367 34595
rect 33367 34561 33376 34595
rect 33324 34552 33376 34561
rect 33600 34595 33652 34604
rect 33600 34561 33609 34595
rect 33609 34561 33643 34595
rect 33643 34561 33652 34595
rect 33600 34552 33652 34561
rect 35900 34620 35952 34672
rect 30840 34527 30892 34536
rect 30840 34493 30849 34527
rect 30849 34493 30883 34527
rect 30883 34493 30892 34527
rect 30840 34484 30892 34493
rect 28356 34416 28408 34468
rect 28724 34459 28776 34468
rect 28724 34425 28733 34459
rect 28733 34425 28767 34459
rect 28767 34425 28776 34459
rect 28724 34416 28776 34425
rect 30104 34416 30156 34468
rect 33968 34484 34020 34536
rect 34244 34484 34296 34536
rect 35532 34595 35584 34604
rect 35532 34561 35541 34595
rect 35541 34561 35575 34595
rect 35575 34561 35584 34595
rect 36728 34620 36780 34672
rect 35532 34552 35584 34561
rect 36452 34552 36504 34604
rect 37556 34595 37608 34604
rect 35440 34484 35492 34536
rect 36268 34484 36320 34536
rect 37556 34561 37565 34595
rect 37565 34561 37599 34595
rect 37599 34561 37608 34595
rect 37556 34552 37608 34561
rect 38108 34552 38160 34604
rect 39120 34595 39172 34604
rect 39120 34561 39129 34595
rect 39129 34561 39163 34595
rect 39163 34561 39172 34595
rect 39120 34552 39172 34561
rect 39304 34595 39356 34604
rect 39304 34561 39313 34595
rect 39313 34561 39347 34595
rect 39347 34561 39356 34595
rect 39304 34552 39356 34561
rect 40408 34595 40460 34604
rect 40408 34561 40417 34595
rect 40417 34561 40451 34595
rect 40451 34561 40460 34595
rect 40408 34552 40460 34561
rect 40592 34595 40644 34604
rect 40592 34561 40601 34595
rect 40601 34561 40635 34595
rect 40635 34561 40644 34595
rect 40592 34552 40644 34561
rect 42064 34484 42116 34536
rect 33692 34416 33744 34468
rect 9772 34391 9824 34400
rect 9772 34357 9781 34391
rect 9781 34357 9815 34391
rect 9815 34357 9824 34391
rect 9772 34348 9824 34357
rect 11520 34348 11572 34400
rect 14832 34348 14884 34400
rect 17960 34348 18012 34400
rect 22008 34348 22060 34400
rect 25044 34391 25096 34400
rect 25044 34357 25053 34391
rect 25053 34357 25087 34391
rect 25087 34357 25096 34391
rect 25044 34348 25096 34357
rect 28448 34391 28500 34400
rect 28448 34357 28457 34391
rect 28457 34357 28491 34391
rect 28491 34357 28500 34391
rect 28448 34348 28500 34357
rect 33968 34348 34020 34400
rect 35716 34416 35768 34468
rect 39856 34348 39908 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 10232 34144 10284 34196
rect 14740 34144 14792 34196
rect 15568 34144 15620 34196
rect 1584 34119 1636 34128
rect 1584 34085 1593 34119
rect 1593 34085 1627 34119
rect 1627 34085 1636 34119
rect 1584 34076 1636 34085
rect 16856 34144 16908 34196
rect 17960 34187 18012 34196
rect 17960 34153 17969 34187
rect 17969 34153 18003 34187
rect 18003 34153 18012 34187
rect 17960 34144 18012 34153
rect 21640 34187 21692 34196
rect 21640 34153 21649 34187
rect 21649 34153 21683 34187
rect 21683 34153 21692 34187
rect 21640 34144 21692 34153
rect 22560 34144 22612 34196
rect 25136 34187 25188 34196
rect 25136 34153 25145 34187
rect 25145 34153 25179 34187
rect 25179 34153 25188 34187
rect 25136 34144 25188 34153
rect 25228 34144 25280 34196
rect 25504 34144 25556 34196
rect 25872 34187 25924 34196
rect 25872 34153 25881 34187
rect 25881 34153 25915 34187
rect 25915 34153 25924 34187
rect 25872 34144 25924 34153
rect 27620 34187 27672 34196
rect 27620 34153 27629 34187
rect 27629 34153 27663 34187
rect 27663 34153 27672 34187
rect 27620 34144 27672 34153
rect 29276 34144 29328 34196
rect 29552 34144 29604 34196
rect 31392 34144 31444 34196
rect 32404 34187 32456 34196
rect 32404 34153 32413 34187
rect 32413 34153 32447 34187
rect 32447 34153 32456 34187
rect 32404 34144 32456 34153
rect 11520 34051 11572 34060
rect 11520 34017 11529 34051
rect 11529 34017 11563 34051
rect 11563 34017 11572 34051
rect 11520 34008 11572 34017
rect 11980 34051 12032 34060
rect 11980 34017 11989 34051
rect 11989 34017 12023 34051
rect 12023 34017 12032 34051
rect 11980 34008 12032 34017
rect 13268 34051 13320 34060
rect 13268 34017 13277 34051
rect 13277 34017 13311 34051
rect 13311 34017 13320 34051
rect 13268 34008 13320 34017
rect 13820 34008 13872 34060
rect 10876 33983 10928 33992
rect 10876 33949 10885 33983
rect 10885 33949 10919 33983
rect 10919 33949 10928 33983
rect 10876 33940 10928 33949
rect 11612 33940 11664 33992
rect 12072 33940 12124 33992
rect 12900 33940 12952 33992
rect 14280 33983 14332 33992
rect 14280 33949 14289 33983
rect 14289 33949 14323 33983
rect 14323 33949 14332 33983
rect 14280 33940 14332 33949
rect 14832 33940 14884 33992
rect 15016 33940 15068 33992
rect 16672 34076 16724 34128
rect 19064 34076 19116 34128
rect 15476 33940 15528 33992
rect 16580 33940 16632 33992
rect 19248 34008 19300 34060
rect 20444 34008 20496 34060
rect 22928 34051 22980 34060
rect 22928 34017 22937 34051
rect 22937 34017 22971 34051
rect 22971 34017 22980 34051
rect 22928 34008 22980 34017
rect 24216 34076 24268 34128
rect 27988 34076 28040 34128
rect 27528 34008 27580 34060
rect 18420 33940 18472 33992
rect 19340 33940 19392 33992
rect 21456 33983 21508 33992
rect 21456 33949 21465 33983
rect 21465 33949 21499 33983
rect 21499 33949 21508 33983
rect 21456 33940 21508 33949
rect 21548 33983 21600 33992
rect 21548 33949 21557 33983
rect 21557 33949 21591 33983
rect 21591 33949 21600 33983
rect 22836 33983 22888 33992
rect 21548 33940 21600 33949
rect 22836 33949 22845 33983
rect 22845 33949 22879 33983
rect 22879 33949 22888 33983
rect 22836 33940 22888 33949
rect 24768 33983 24820 33992
rect 24768 33949 24777 33983
rect 24777 33949 24811 33983
rect 24811 33949 24820 33983
rect 24768 33940 24820 33949
rect 26792 33983 26844 33992
rect 26792 33949 26801 33983
rect 26801 33949 26835 33983
rect 26835 33949 26844 33983
rect 26792 33940 26844 33949
rect 26976 33983 27028 33992
rect 26976 33949 26985 33983
rect 26985 33949 27019 33983
rect 27019 33949 27028 33983
rect 26976 33940 27028 33949
rect 28264 33940 28316 33992
rect 28448 33983 28500 33992
rect 28448 33949 28457 33983
rect 28457 33949 28491 33983
rect 28491 33949 28500 33983
rect 28448 33940 28500 33949
rect 30840 34076 30892 34128
rect 32312 34008 32364 34060
rect 30932 33940 30984 33992
rect 31300 33983 31352 33992
rect 31300 33949 31309 33983
rect 31309 33949 31343 33983
rect 31343 33949 31352 33983
rect 31300 33940 31352 33949
rect 18696 33872 18748 33924
rect 20996 33872 21048 33924
rect 25412 33872 25464 33924
rect 27712 33872 27764 33924
rect 9772 33847 9824 33856
rect 9772 33813 9781 33847
rect 9781 33813 9815 33847
rect 9815 33813 9824 33847
rect 9772 33804 9824 33813
rect 12624 33804 12676 33856
rect 14464 33804 14516 33856
rect 18512 33804 18564 33856
rect 18972 33804 19024 33856
rect 20536 33847 20588 33856
rect 20536 33813 20545 33847
rect 20545 33813 20579 33847
rect 20579 33813 20588 33847
rect 20536 33804 20588 33813
rect 26976 33847 27028 33856
rect 26976 33813 26985 33847
rect 26985 33813 27019 33847
rect 27019 33813 27028 33847
rect 26976 33804 27028 33813
rect 27620 33847 27672 33856
rect 27620 33813 27629 33847
rect 27629 33813 27663 33847
rect 27663 33813 27672 33847
rect 27620 33804 27672 33813
rect 28540 33847 28592 33856
rect 28540 33813 28549 33847
rect 28549 33813 28583 33847
rect 28583 33813 28592 33847
rect 28540 33804 28592 33813
rect 30288 33915 30340 33924
rect 30288 33881 30323 33915
rect 30323 33881 30340 33915
rect 30288 33872 30340 33881
rect 31392 33872 31444 33924
rect 31576 33804 31628 33856
rect 33140 34008 33192 34060
rect 33784 34144 33836 34196
rect 34428 34144 34480 34196
rect 35440 34144 35492 34196
rect 36268 34144 36320 34196
rect 39672 34144 39724 34196
rect 42064 34187 42116 34196
rect 42064 34153 42073 34187
rect 42073 34153 42107 34187
rect 42107 34153 42116 34187
rect 42064 34144 42116 34153
rect 37556 34076 37608 34128
rect 35348 34008 35400 34060
rect 35532 34051 35584 34060
rect 35532 34017 35541 34051
rect 35541 34017 35575 34051
rect 35575 34017 35584 34051
rect 35532 34008 35584 34017
rect 38200 34051 38252 34060
rect 38200 34017 38209 34051
rect 38209 34017 38243 34051
rect 38243 34017 38252 34051
rect 38200 34008 38252 34017
rect 40316 34076 40368 34128
rect 40776 34076 40828 34128
rect 42524 34119 42576 34128
rect 42524 34085 42533 34119
rect 42533 34085 42567 34119
rect 42567 34085 42576 34119
rect 42524 34076 42576 34085
rect 38660 34051 38712 34060
rect 38660 34017 38694 34051
rect 38694 34017 38712 34051
rect 38660 34008 38712 34017
rect 33324 33940 33376 33992
rect 33692 33940 33744 33992
rect 33968 33940 34020 33992
rect 35808 33983 35860 33992
rect 33048 33872 33100 33924
rect 35808 33949 35817 33983
rect 35817 33949 35851 33983
rect 35851 33949 35860 33983
rect 35808 33940 35860 33949
rect 36176 33940 36228 33992
rect 36452 33983 36504 33992
rect 36452 33949 36461 33983
rect 36461 33949 36495 33983
rect 36495 33949 36504 33983
rect 36452 33940 36504 33949
rect 37372 33983 37424 33992
rect 37372 33949 37381 33983
rect 37381 33949 37415 33983
rect 37415 33949 37424 33983
rect 37372 33940 37424 33949
rect 38108 33940 38160 33992
rect 40592 34008 40644 34060
rect 48136 34051 48188 34060
rect 48136 34017 48145 34051
rect 48145 34017 48179 34051
rect 48179 34017 48188 34051
rect 48136 34008 48188 34017
rect 33784 33804 33836 33856
rect 33968 33847 34020 33856
rect 33968 33813 33977 33847
rect 33977 33813 34011 33847
rect 34011 33813 34020 33847
rect 33968 33804 34020 33813
rect 35900 33872 35952 33924
rect 40776 33940 40828 33992
rect 47860 33983 47912 33992
rect 36084 33804 36136 33856
rect 37832 33804 37884 33856
rect 40684 33804 40736 33856
rect 47860 33949 47869 33983
rect 47869 33949 47903 33983
rect 47903 33949 47912 33983
rect 47860 33940 47912 33949
rect 43168 33847 43220 33856
rect 43168 33813 43177 33847
rect 43177 33813 43211 33847
rect 43211 33813 43220 33847
rect 43168 33804 43220 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 2044 33600 2096 33652
rect 10876 33600 10928 33652
rect 13268 33600 13320 33652
rect 15384 33600 15436 33652
rect 11152 33532 11204 33584
rect 11704 33575 11756 33584
rect 11704 33541 11713 33575
rect 11713 33541 11747 33575
rect 11747 33541 11756 33575
rect 11704 33532 11756 33541
rect 12716 33575 12768 33584
rect 12716 33541 12725 33575
rect 12725 33541 12759 33575
rect 12759 33541 12768 33575
rect 12716 33532 12768 33541
rect 12900 33575 12952 33584
rect 12900 33541 12909 33575
rect 12909 33541 12943 33575
rect 12943 33541 12952 33575
rect 12900 33532 12952 33541
rect 13452 33532 13504 33584
rect 11520 33507 11572 33516
rect 11520 33473 11529 33507
rect 11529 33473 11563 33507
rect 11563 33473 11572 33507
rect 11520 33464 11572 33473
rect 12808 33464 12860 33516
rect 13820 33507 13872 33516
rect 13820 33473 13829 33507
rect 13829 33473 13863 33507
rect 13863 33473 13872 33507
rect 13820 33464 13872 33473
rect 14464 33464 14516 33516
rect 15016 33507 15068 33516
rect 15016 33473 15025 33507
rect 15025 33473 15059 33507
rect 15059 33473 15068 33507
rect 15016 33464 15068 33473
rect 15292 33464 15344 33516
rect 18144 33600 18196 33652
rect 19248 33643 19300 33652
rect 19248 33609 19257 33643
rect 19257 33609 19291 33643
rect 19291 33609 19300 33643
rect 19248 33600 19300 33609
rect 15660 33507 15712 33516
rect 15660 33473 15669 33507
rect 15669 33473 15703 33507
rect 15703 33473 15712 33507
rect 15660 33464 15712 33473
rect 14096 33396 14148 33448
rect 18696 33532 18748 33584
rect 20076 33532 20128 33584
rect 18052 33464 18104 33516
rect 18144 33507 18196 33516
rect 18144 33473 18153 33507
rect 18153 33473 18187 33507
rect 18187 33473 18196 33507
rect 18144 33464 18196 33473
rect 18328 33464 18380 33516
rect 18512 33464 18564 33516
rect 24124 33600 24176 33652
rect 24768 33600 24820 33652
rect 21088 33532 21140 33584
rect 22284 33532 22336 33584
rect 22468 33532 22520 33584
rect 20536 33464 20588 33516
rect 22836 33507 22888 33516
rect 18420 33396 18472 33448
rect 16580 33328 16632 33380
rect 16764 33328 16816 33380
rect 18696 33396 18748 33448
rect 18880 33328 18932 33380
rect 19248 33396 19300 33448
rect 20168 33439 20220 33448
rect 20168 33405 20177 33439
rect 20177 33405 20211 33439
rect 20211 33405 20220 33439
rect 22836 33473 22845 33507
rect 22845 33473 22879 33507
rect 22879 33473 22888 33507
rect 22836 33464 22888 33473
rect 23112 33464 23164 33516
rect 23480 33464 23532 33516
rect 20168 33396 20220 33405
rect 23296 33396 23348 33448
rect 24768 33464 24820 33516
rect 25044 33464 25096 33516
rect 25228 33464 25280 33516
rect 27620 33600 27672 33652
rect 27896 33600 27948 33652
rect 25780 33507 25832 33516
rect 25780 33473 25789 33507
rect 25789 33473 25823 33507
rect 25823 33473 25832 33507
rect 25780 33464 25832 33473
rect 27344 33507 27396 33516
rect 27344 33473 27353 33507
rect 27353 33473 27387 33507
rect 27387 33473 27396 33507
rect 27344 33464 27396 33473
rect 27436 33507 27488 33516
rect 27436 33473 27445 33507
rect 27445 33473 27479 33507
rect 27479 33473 27488 33507
rect 27712 33507 27764 33516
rect 27436 33464 27488 33473
rect 27712 33473 27721 33507
rect 27721 33473 27755 33507
rect 27755 33473 27764 33507
rect 27712 33464 27764 33473
rect 28356 33600 28408 33652
rect 29920 33600 29972 33652
rect 30840 33600 30892 33652
rect 31484 33600 31536 33652
rect 31944 33532 31996 33584
rect 33600 33600 33652 33652
rect 36176 33643 36228 33652
rect 36176 33609 36185 33643
rect 36185 33609 36219 33643
rect 36219 33609 36228 33643
rect 36176 33600 36228 33609
rect 36268 33600 36320 33652
rect 34520 33532 34572 33584
rect 29184 33464 29236 33516
rect 30380 33507 30432 33516
rect 30380 33473 30389 33507
rect 30389 33473 30423 33507
rect 30423 33473 30432 33507
rect 30380 33464 30432 33473
rect 31300 33464 31352 33516
rect 31392 33507 31444 33516
rect 31392 33473 31401 33507
rect 31401 33473 31435 33507
rect 31435 33473 31444 33507
rect 31392 33464 31444 33473
rect 26976 33396 27028 33448
rect 30472 33439 30524 33448
rect 30472 33405 30481 33439
rect 30481 33405 30515 33439
rect 30515 33405 30524 33439
rect 30472 33396 30524 33405
rect 30564 33396 30616 33448
rect 32128 33396 32180 33448
rect 32404 33507 32456 33516
rect 32404 33473 32413 33507
rect 32413 33473 32447 33507
rect 32447 33473 32456 33507
rect 32588 33507 32640 33516
rect 32404 33464 32456 33473
rect 32588 33473 32597 33507
rect 32597 33473 32631 33507
rect 32631 33473 32640 33507
rect 32588 33464 32640 33473
rect 35532 33532 35584 33584
rect 36452 33532 36504 33584
rect 37556 33600 37608 33652
rect 38660 33643 38712 33652
rect 38660 33609 38669 33643
rect 38669 33609 38703 33643
rect 38703 33609 38712 33643
rect 38660 33600 38712 33609
rect 36176 33464 36228 33516
rect 38384 33532 38436 33584
rect 40408 33532 40460 33584
rect 32956 33396 33008 33448
rect 34520 33439 34572 33448
rect 34520 33405 34529 33439
rect 34529 33405 34563 33439
rect 34563 33405 34572 33439
rect 34520 33396 34572 33405
rect 21272 33328 21324 33380
rect 24216 33328 24268 33380
rect 24768 33328 24820 33380
rect 25136 33371 25188 33380
rect 25136 33337 25145 33371
rect 25145 33337 25179 33371
rect 25179 33337 25188 33371
rect 25136 33328 25188 33337
rect 34336 33328 34388 33380
rect 35624 33396 35676 33448
rect 36176 33328 36228 33380
rect 37740 33464 37792 33516
rect 38108 33464 38160 33516
rect 39120 33507 39172 33516
rect 39120 33473 39129 33507
rect 39129 33473 39163 33507
rect 39163 33473 39172 33507
rect 39120 33464 39172 33473
rect 39304 33507 39356 33516
rect 39304 33473 39313 33507
rect 39313 33473 39347 33507
rect 39347 33473 39356 33507
rect 39304 33464 39356 33473
rect 39580 33507 39632 33516
rect 39580 33473 39589 33507
rect 39589 33473 39623 33507
rect 39623 33473 39632 33507
rect 39580 33464 39632 33473
rect 40132 33464 40184 33516
rect 41052 33600 41104 33652
rect 48136 33643 48188 33652
rect 48136 33609 48145 33643
rect 48145 33609 48179 33643
rect 48179 33609 48188 33643
rect 48136 33600 48188 33609
rect 40684 33507 40736 33516
rect 40684 33473 40693 33507
rect 40693 33473 40727 33507
rect 40727 33473 40736 33507
rect 40684 33464 40736 33473
rect 38016 33396 38068 33448
rect 40040 33396 40092 33448
rect 39856 33328 39908 33380
rect 40868 33507 40920 33516
rect 40868 33473 40877 33507
rect 40877 33473 40911 33507
rect 40911 33473 40920 33507
rect 43076 33532 43128 33584
rect 40868 33464 40920 33473
rect 41052 33507 41104 33516
rect 41052 33473 41061 33507
rect 41061 33473 41095 33507
rect 41095 33473 41104 33507
rect 41052 33464 41104 33473
rect 47860 33464 47912 33516
rect 41420 33328 41472 33380
rect 12716 33260 12768 33312
rect 15568 33260 15620 33312
rect 18144 33260 18196 33312
rect 25688 33303 25740 33312
rect 25688 33269 25697 33303
rect 25697 33269 25731 33303
rect 25731 33269 25740 33303
rect 25688 33260 25740 33269
rect 27160 33260 27212 33312
rect 29920 33260 29972 33312
rect 31484 33260 31536 33312
rect 32220 33260 32272 33312
rect 33232 33260 33284 33312
rect 34428 33260 34480 33312
rect 40408 33303 40460 33312
rect 40408 33269 40417 33303
rect 40417 33269 40451 33303
rect 40451 33269 40460 33303
rect 40408 33260 40460 33269
rect 40776 33260 40828 33312
rect 40868 33260 40920 33312
rect 43168 33260 43220 33312
rect 44180 33260 44232 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 11612 33099 11664 33108
rect 11612 33065 11621 33099
rect 11621 33065 11655 33099
rect 11655 33065 11664 33099
rect 11612 33056 11664 33065
rect 12440 33056 12492 33108
rect 17132 33056 17184 33108
rect 17868 33056 17920 33108
rect 20168 33099 20220 33108
rect 20168 33065 20177 33099
rect 20177 33065 20211 33099
rect 20211 33065 20220 33099
rect 20168 33056 20220 33065
rect 20720 33099 20772 33108
rect 20720 33065 20729 33099
rect 20729 33065 20763 33099
rect 20763 33065 20772 33099
rect 20720 33056 20772 33065
rect 22192 33056 22244 33108
rect 22836 33099 22888 33108
rect 22836 33065 22845 33099
rect 22845 33065 22879 33099
rect 22879 33065 22888 33099
rect 22836 33056 22888 33065
rect 22928 33056 22980 33108
rect 23388 33099 23440 33108
rect 23388 33065 23397 33099
rect 23397 33065 23431 33099
rect 23431 33065 23440 33099
rect 23388 33056 23440 33065
rect 25780 33056 25832 33108
rect 27528 33056 27580 33108
rect 28448 33056 28500 33108
rect 29644 33056 29696 33108
rect 30472 33056 30524 33108
rect 18880 32988 18932 33040
rect 23296 32988 23348 33040
rect 11980 32920 12032 32972
rect 11520 32895 11572 32904
rect 11520 32861 11529 32895
rect 11529 32861 11563 32895
rect 11563 32861 11572 32895
rect 11520 32852 11572 32861
rect 11704 32895 11756 32904
rect 11704 32861 11713 32895
rect 11713 32861 11747 32895
rect 11747 32861 11756 32895
rect 11704 32852 11756 32861
rect 12808 32895 12860 32904
rect 12808 32861 12817 32895
rect 12817 32861 12851 32895
rect 12851 32861 12860 32895
rect 12808 32852 12860 32861
rect 12992 32852 13044 32904
rect 13820 32852 13872 32904
rect 13452 32784 13504 32836
rect 13176 32716 13228 32768
rect 15292 32852 15344 32904
rect 15752 32920 15804 32972
rect 19340 32920 19392 32972
rect 25688 32963 25740 32972
rect 25688 32929 25697 32963
rect 25697 32929 25731 32963
rect 25731 32929 25740 32963
rect 25688 32920 25740 32929
rect 26792 32988 26844 33040
rect 31116 32988 31168 33040
rect 32128 32920 32180 32972
rect 15568 32895 15620 32904
rect 15568 32861 15577 32895
rect 15577 32861 15611 32895
rect 15611 32861 15620 32895
rect 15568 32852 15620 32861
rect 15936 32895 15988 32904
rect 15936 32861 15945 32895
rect 15945 32861 15979 32895
rect 15979 32861 15988 32895
rect 15936 32852 15988 32861
rect 16672 32852 16724 32904
rect 17040 32895 17092 32904
rect 17040 32861 17049 32895
rect 17049 32861 17083 32895
rect 17083 32861 17092 32895
rect 17040 32852 17092 32861
rect 17316 32895 17368 32904
rect 17316 32861 17325 32895
rect 17325 32861 17359 32895
rect 17359 32861 17368 32895
rect 17316 32852 17368 32861
rect 17500 32895 17552 32904
rect 17500 32861 17509 32895
rect 17509 32861 17543 32895
rect 17543 32861 17552 32895
rect 17500 32852 17552 32861
rect 17960 32895 18012 32904
rect 17960 32861 17969 32895
rect 17969 32861 18003 32895
rect 18003 32861 18012 32895
rect 17960 32852 18012 32861
rect 18144 32895 18196 32904
rect 18144 32861 18153 32895
rect 18153 32861 18187 32895
rect 18187 32861 18196 32895
rect 18144 32852 18196 32861
rect 19984 32895 20036 32904
rect 19984 32861 19993 32895
rect 19993 32861 20027 32895
rect 20027 32861 20036 32895
rect 19984 32852 20036 32861
rect 20444 32852 20496 32904
rect 20996 32852 21048 32904
rect 21732 32895 21784 32904
rect 21732 32861 21747 32895
rect 21747 32861 21781 32895
rect 21781 32861 21784 32895
rect 21916 32895 21968 32904
rect 21732 32852 21784 32861
rect 21916 32861 21925 32895
rect 21925 32861 21959 32895
rect 21959 32861 21968 32895
rect 21916 32852 21968 32861
rect 22376 32895 22428 32904
rect 22376 32861 22385 32895
rect 22385 32861 22419 32895
rect 22419 32861 22428 32895
rect 22376 32852 22428 32861
rect 22652 32895 22704 32904
rect 22652 32861 22661 32895
rect 22661 32861 22695 32895
rect 22695 32861 22704 32895
rect 22652 32852 22704 32861
rect 23112 32852 23164 32904
rect 23480 32895 23532 32904
rect 23480 32861 23489 32895
rect 23489 32861 23523 32895
rect 23523 32861 23532 32895
rect 23480 32852 23532 32861
rect 24768 32895 24820 32904
rect 24768 32861 24777 32895
rect 24777 32861 24811 32895
rect 24811 32861 24820 32895
rect 24768 32852 24820 32861
rect 24860 32852 24912 32904
rect 25504 32852 25556 32904
rect 25964 32852 26016 32904
rect 26700 32895 26752 32904
rect 26700 32861 26709 32895
rect 26709 32861 26743 32895
rect 26743 32861 26752 32895
rect 26700 32852 26752 32861
rect 21824 32784 21876 32836
rect 26608 32784 26660 32836
rect 27068 32852 27120 32904
rect 28356 32895 28408 32904
rect 28356 32861 28365 32895
rect 28365 32861 28399 32895
rect 28399 32861 28408 32895
rect 28356 32852 28408 32861
rect 27896 32784 27948 32836
rect 14740 32716 14792 32768
rect 18052 32759 18104 32768
rect 18052 32725 18061 32759
rect 18061 32725 18095 32759
rect 18095 32725 18104 32759
rect 18052 32716 18104 32725
rect 18788 32716 18840 32768
rect 22284 32716 22336 32768
rect 27620 32716 27672 32768
rect 27804 32716 27856 32768
rect 29552 32852 29604 32904
rect 30288 32852 30340 32904
rect 30564 32895 30616 32904
rect 30564 32861 30573 32895
rect 30573 32861 30607 32895
rect 30607 32861 30616 32895
rect 33140 33056 33192 33108
rect 34060 33056 34112 33108
rect 36084 33056 36136 33108
rect 37372 33056 37424 33108
rect 37924 33056 37976 33108
rect 40040 33056 40092 33108
rect 40868 33099 40920 33108
rect 40868 33065 40877 33099
rect 40877 33065 40911 33099
rect 40911 33065 40920 33099
rect 40868 33056 40920 33065
rect 32680 32988 32732 33040
rect 30564 32852 30616 32861
rect 32772 32895 32824 32904
rect 32404 32784 32456 32836
rect 32772 32861 32781 32895
rect 32781 32861 32815 32895
rect 32815 32861 32824 32895
rect 32772 32852 32824 32861
rect 32864 32895 32916 32904
rect 32864 32861 32873 32895
rect 32873 32861 32907 32895
rect 32907 32861 32916 32895
rect 32864 32852 32916 32861
rect 28816 32716 28868 32768
rect 29644 32759 29696 32768
rect 29644 32725 29653 32759
rect 29653 32725 29687 32759
rect 29687 32725 29696 32759
rect 29644 32716 29696 32725
rect 30840 32716 30892 32768
rect 33416 32784 33468 32836
rect 33784 32988 33836 33040
rect 39856 32988 39908 33040
rect 41420 33031 41472 33040
rect 41420 32997 41429 33031
rect 41429 32997 41463 33031
rect 41463 32997 41472 33031
rect 41420 32988 41472 32997
rect 42524 33031 42576 33040
rect 42524 32997 42533 33031
rect 42533 32997 42567 33031
rect 42567 32997 42576 33031
rect 42524 32988 42576 32997
rect 34796 32852 34848 32904
rect 34980 32895 35032 32904
rect 34980 32861 34989 32895
rect 34989 32861 35023 32895
rect 35023 32861 35032 32895
rect 34980 32852 35032 32861
rect 35716 32852 35768 32904
rect 37648 32895 37700 32904
rect 37648 32861 37657 32895
rect 37657 32861 37691 32895
rect 37691 32861 37700 32895
rect 37648 32852 37700 32861
rect 38108 32895 38160 32904
rect 38108 32861 38117 32895
rect 38117 32861 38151 32895
rect 38151 32861 38160 32895
rect 38108 32852 38160 32861
rect 38384 32852 38436 32904
rect 39948 32852 40000 32904
rect 40684 32920 40736 32972
rect 40316 32895 40368 32904
rect 40316 32861 40325 32895
rect 40325 32861 40359 32895
rect 40359 32861 40368 32895
rect 40316 32852 40368 32861
rect 40408 32895 40460 32904
rect 40408 32861 40417 32895
rect 40417 32861 40451 32895
rect 40451 32861 40460 32895
rect 40408 32852 40460 32861
rect 37740 32784 37792 32836
rect 34704 32716 34756 32768
rect 38660 32716 38712 32768
rect 39672 32716 39724 32768
rect 41512 32716 41564 32768
rect 41972 32759 42024 32768
rect 41972 32725 41981 32759
rect 41981 32725 42015 32759
rect 42015 32725 42024 32759
rect 41972 32716 42024 32725
rect 47860 32716 47912 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 10692 32512 10744 32564
rect 14188 32512 14240 32564
rect 16672 32555 16724 32564
rect 1584 32376 1636 32428
rect 12624 32419 12676 32428
rect 12624 32385 12633 32419
rect 12633 32385 12667 32419
rect 12667 32385 12676 32419
rect 12624 32376 12676 32385
rect 12716 32419 12768 32428
rect 12716 32385 12725 32419
rect 12725 32385 12759 32419
rect 12759 32385 12768 32419
rect 13820 32444 13872 32496
rect 12716 32376 12768 32385
rect 13176 32376 13228 32428
rect 13268 32308 13320 32360
rect 14188 32308 14240 32360
rect 15292 32487 15344 32496
rect 15292 32453 15301 32487
rect 15301 32453 15335 32487
rect 15335 32453 15344 32487
rect 15292 32444 15344 32453
rect 16672 32521 16681 32555
rect 16681 32521 16715 32555
rect 16715 32521 16724 32555
rect 16672 32512 16724 32521
rect 17408 32512 17460 32564
rect 19432 32512 19484 32564
rect 22652 32512 22704 32564
rect 25964 32555 26016 32564
rect 16856 32419 16908 32428
rect 16856 32385 16865 32419
rect 16865 32385 16899 32419
rect 16899 32385 16908 32419
rect 16856 32376 16908 32385
rect 17316 32376 17368 32428
rect 17868 32444 17920 32496
rect 21824 32444 21876 32496
rect 22008 32444 22060 32496
rect 18328 32376 18380 32428
rect 14740 32308 14792 32360
rect 17500 32308 17552 32360
rect 18236 32308 18288 32360
rect 19340 32376 19392 32428
rect 19984 32376 20036 32428
rect 20996 32376 21048 32428
rect 21456 32376 21508 32428
rect 22100 32376 22152 32428
rect 22284 32376 22336 32428
rect 23572 32444 23624 32496
rect 25964 32521 25973 32555
rect 25973 32521 26007 32555
rect 26007 32521 26016 32555
rect 25964 32512 26016 32521
rect 27804 32512 27856 32564
rect 24952 32444 25004 32496
rect 23388 32419 23440 32428
rect 23388 32385 23397 32419
rect 23397 32385 23431 32419
rect 23431 32385 23440 32419
rect 23388 32376 23440 32385
rect 22468 32308 22520 32360
rect 23296 32308 23348 32360
rect 12808 32283 12860 32292
rect 12808 32249 12817 32283
rect 12817 32249 12851 32283
rect 12851 32249 12860 32283
rect 12808 32240 12860 32249
rect 16672 32240 16724 32292
rect 17960 32240 18012 32292
rect 20444 32240 20496 32292
rect 1952 32215 2004 32224
rect 1952 32181 1961 32215
rect 1961 32181 1995 32215
rect 1995 32181 2004 32215
rect 1952 32172 2004 32181
rect 8944 32172 8996 32224
rect 11980 32215 12032 32224
rect 11980 32181 11989 32215
rect 11989 32181 12023 32215
rect 12023 32181 12032 32215
rect 11980 32172 12032 32181
rect 13544 32215 13596 32224
rect 13544 32181 13553 32215
rect 13553 32181 13587 32215
rect 13587 32181 13596 32215
rect 13544 32172 13596 32181
rect 14832 32172 14884 32224
rect 15200 32172 15252 32224
rect 17040 32172 17092 32224
rect 17592 32172 17644 32224
rect 20720 32172 20772 32224
rect 20812 32172 20864 32224
rect 22284 32240 22336 32292
rect 23480 32240 23532 32292
rect 24676 32240 24728 32292
rect 25504 32419 25556 32428
rect 25504 32385 25513 32419
rect 25513 32385 25547 32419
rect 25547 32385 25556 32419
rect 25504 32376 25556 32385
rect 26792 32376 26844 32428
rect 27528 32444 27580 32496
rect 27988 32444 28040 32496
rect 28540 32512 28592 32564
rect 29552 32555 29604 32564
rect 29552 32521 29561 32555
rect 29561 32521 29595 32555
rect 29595 32521 29604 32555
rect 29552 32512 29604 32521
rect 31484 32555 31536 32564
rect 31484 32521 31493 32555
rect 31493 32521 31527 32555
rect 31527 32521 31536 32555
rect 31484 32512 31536 32521
rect 32772 32512 32824 32564
rect 32956 32512 33008 32564
rect 33968 32555 34020 32564
rect 33968 32521 33977 32555
rect 33977 32521 34011 32555
rect 34011 32521 34020 32555
rect 33968 32512 34020 32521
rect 35348 32512 35400 32564
rect 35900 32512 35952 32564
rect 37648 32512 37700 32564
rect 39856 32512 39908 32564
rect 30748 32487 30800 32496
rect 27160 32419 27212 32428
rect 27160 32385 27169 32419
rect 27169 32385 27203 32419
rect 27203 32385 27212 32419
rect 27160 32376 27212 32385
rect 27620 32376 27672 32428
rect 28816 32419 28868 32428
rect 27804 32351 27856 32360
rect 27804 32317 27813 32351
rect 27813 32317 27847 32351
rect 27847 32317 27856 32351
rect 27804 32308 27856 32317
rect 28264 32308 28316 32360
rect 28816 32385 28825 32419
rect 28825 32385 28859 32419
rect 28859 32385 28868 32419
rect 28816 32376 28868 32385
rect 29736 32419 29788 32428
rect 29736 32385 29745 32419
rect 29745 32385 29779 32419
rect 29779 32385 29788 32419
rect 29736 32376 29788 32385
rect 29920 32419 29972 32428
rect 29920 32385 29929 32419
rect 29929 32385 29963 32419
rect 29963 32385 29972 32419
rect 29920 32376 29972 32385
rect 30748 32453 30757 32487
rect 30757 32453 30791 32487
rect 30791 32453 30800 32487
rect 30748 32444 30800 32453
rect 30840 32444 30892 32496
rect 31576 32444 31628 32496
rect 32128 32444 32180 32496
rect 33416 32444 33468 32496
rect 30656 32419 30708 32428
rect 29368 32308 29420 32360
rect 29644 32308 29696 32360
rect 30656 32385 30665 32419
rect 30665 32385 30699 32419
rect 30699 32385 30708 32419
rect 30656 32376 30708 32385
rect 34704 32444 34756 32496
rect 33784 32419 33836 32428
rect 33784 32385 33793 32419
rect 33793 32385 33827 32419
rect 33827 32385 33836 32419
rect 33784 32376 33836 32385
rect 34060 32419 34112 32428
rect 34060 32385 34069 32419
rect 34069 32385 34103 32419
rect 34103 32385 34112 32419
rect 34060 32376 34112 32385
rect 34796 32419 34848 32428
rect 34796 32385 34805 32419
rect 34805 32385 34839 32419
rect 34839 32385 34848 32419
rect 34796 32376 34848 32385
rect 35440 32376 35492 32428
rect 35716 32419 35768 32428
rect 35716 32385 35725 32419
rect 35725 32385 35759 32419
rect 35759 32385 35768 32419
rect 35716 32376 35768 32385
rect 38660 32444 38712 32496
rect 39672 32444 39724 32496
rect 37464 32419 37516 32428
rect 32404 32308 32456 32360
rect 32680 32308 32732 32360
rect 33324 32308 33376 32360
rect 34980 32308 35032 32360
rect 35900 32351 35952 32360
rect 35900 32317 35909 32351
rect 35909 32317 35943 32351
rect 35943 32317 35952 32351
rect 35900 32308 35952 32317
rect 25228 32240 25280 32292
rect 25596 32240 25648 32292
rect 28356 32240 28408 32292
rect 28632 32240 28684 32292
rect 30932 32283 30984 32292
rect 22192 32172 22244 32224
rect 27896 32172 27948 32224
rect 29000 32172 29052 32224
rect 29736 32172 29788 32224
rect 30012 32172 30064 32224
rect 30932 32249 30941 32283
rect 30941 32249 30975 32283
rect 30975 32249 30984 32283
rect 30932 32240 30984 32249
rect 30840 32172 30892 32224
rect 33968 32172 34020 32224
rect 34520 32172 34572 32224
rect 35808 32240 35860 32292
rect 37464 32385 37473 32419
rect 37473 32385 37507 32419
rect 37507 32385 37516 32419
rect 37464 32376 37516 32385
rect 37740 32376 37792 32428
rect 38108 32376 38160 32428
rect 38752 32376 38804 32428
rect 43260 32376 43312 32428
rect 47676 32376 47728 32428
rect 38384 32308 38436 32360
rect 39580 32308 39632 32360
rect 40960 32308 41012 32360
rect 38568 32240 38620 32292
rect 36544 32172 36596 32224
rect 40408 32172 40460 32224
rect 41972 32172 42024 32224
rect 48044 32215 48096 32224
rect 48044 32181 48053 32215
rect 48053 32181 48087 32215
rect 48087 32181 48096 32215
rect 48044 32172 48096 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 1584 32011 1636 32020
rect 1584 31977 1593 32011
rect 1593 31977 1627 32011
rect 1627 31977 1636 32011
rect 1584 31968 1636 31977
rect 10692 32011 10744 32020
rect 10692 31977 10701 32011
rect 10701 31977 10735 32011
rect 10735 31977 10744 32011
rect 10692 31968 10744 31977
rect 11796 32011 11848 32020
rect 11796 31977 11805 32011
rect 11805 31977 11839 32011
rect 11839 31977 11848 32011
rect 11796 31968 11848 31977
rect 12808 31968 12860 32020
rect 1952 31900 2004 31952
rect 15200 31900 15252 31952
rect 13728 31832 13780 31884
rect 15660 31968 15712 32020
rect 16580 32011 16632 32020
rect 16580 31977 16589 32011
rect 16589 31977 16623 32011
rect 16623 31977 16632 32011
rect 16580 31968 16632 31977
rect 19340 31968 19392 32020
rect 18880 31900 18932 31952
rect 20812 31943 20864 31952
rect 12348 31807 12400 31816
rect 12348 31773 12357 31807
rect 12357 31773 12391 31807
rect 12391 31773 12400 31807
rect 12348 31764 12400 31773
rect 12532 31764 12584 31816
rect 13544 31764 13596 31816
rect 13636 31764 13688 31816
rect 13820 31764 13872 31816
rect 14188 31807 14240 31816
rect 14188 31773 14197 31807
rect 14197 31773 14231 31807
rect 14231 31773 14240 31807
rect 14188 31764 14240 31773
rect 14832 31764 14884 31816
rect 13728 31628 13780 31680
rect 17132 31807 17184 31816
rect 17132 31773 17141 31807
rect 17141 31773 17175 31807
rect 17175 31773 17184 31807
rect 17132 31764 17184 31773
rect 17408 31807 17460 31816
rect 17408 31773 17417 31807
rect 17417 31773 17451 31807
rect 17451 31773 17460 31807
rect 17408 31764 17460 31773
rect 17868 31764 17920 31816
rect 15016 31739 15068 31748
rect 15016 31705 15043 31739
rect 15043 31705 15068 31739
rect 15016 31696 15068 31705
rect 15384 31696 15436 31748
rect 17500 31696 17552 31748
rect 18328 31807 18380 31816
rect 18328 31773 18337 31807
rect 18337 31773 18371 31807
rect 18371 31773 18380 31807
rect 18328 31764 18380 31773
rect 18788 31764 18840 31816
rect 19432 31807 19484 31816
rect 19432 31773 19441 31807
rect 19441 31773 19475 31807
rect 19475 31773 19484 31807
rect 19432 31764 19484 31773
rect 20812 31909 20821 31943
rect 20821 31909 20855 31943
rect 20855 31909 20864 31943
rect 20812 31900 20864 31909
rect 22284 31900 22336 31952
rect 20720 31875 20772 31884
rect 20720 31841 20729 31875
rect 20729 31841 20763 31875
rect 20763 31841 20772 31875
rect 20720 31832 20772 31841
rect 22376 31832 22428 31884
rect 22652 31900 22704 31952
rect 25504 31968 25556 32020
rect 25596 32011 25648 32020
rect 25596 31977 25605 32011
rect 25605 31977 25639 32011
rect 25639 31977 25648 32011
rect 25596 31968 25648 31977
rect 28080 31968 28132 32020
rect 28356 31968 28408 32020
rect 29000 32011 29052 32020
rect 21088 31807 21140 31816
rect 21088 31773 21097 31807
rect 21097 31773 21131 31807
rect 21131 31773 21140 31807
rect 21088 31764 21140 31773
rect 21732 31764 21784 31816
rect 23112 31832 23164 31884
rect 21916 31696 21968 31748
rect 26700 31900 26752 31952
rect 27804 31900 27856 31952
rect 29000 31977 29009 32011
rect 29009 31977 29043 32011
rect 29043 31977 29052 32011
rect 29000 31968 29052 31977
rect 29920 31968 29972 32020
rect 30656 31968 30708 32020
rect 30840 31968 30892 32020
rect 32588 31968 32640 32020
rect 34060 31968 34112 32020
rect 34796 32011 34848 32020
rect 34796 31977 34805 32011
rect 34805 31977 34839 32011
rect 34839 31977 34848 32011
rect 34796 31968 34848 31977
rect 38384 31968 38436 32020
rect 40408 32011 40460 32020
rect 40408 31977 40417 32011
rect 40417 31977 40451 32011
rect 40451 31977 40460 32011
rect 40408 31968 40460 31977
rect 40684 31968 40736 32020
rect 47676 32011 47728 32020
rect 47676 31977 47685 32011
rect 47685 31977 47719 32011
rect 47719 31977 47728 32011
rect 47676 31968 47728 31977
rect 23572 31875 23624 31884
rect 23572 31841 23581 31875
rect 23581 31841 23615 31875
rect 23615 31841 23624 31875
rect 23572 31832 23624 31841
rect 25688 31832 25740 31884
rect 28264 31832 28316 31884
rect 28356 31832 28408 31884
rect 29644 31875 29696 31884
rect 23480 31764 23532 31816
rect 24952 31764 25004 31816
rect 25780 31807 25832 31816
rect 25780 31773 25789 31807
rect 25789 31773 25823 31807
rect 25823 31773 25832 31807
rect 25780 31764 25832 31773
rect 26608 31764 26660 31816
rect 27068 31764 27120 31816
rect 27620 31807 27672 31816
rect 24308 31696 24360 31748
rect 24676 31739 24728 31748
rect 24676 31705 24685 31739
rect 24685 31705 24719 31739
rect 24719 31705 24728 31739
rect 24676 31696 24728 31705
rect 26792 31739 26844 31748
rect 26792 31705 26801 31739
rect 26801 31705 26835 31739
rect 26835 31705 26844 31739
rect 26792 31696 26844 31705
rect 27620 31773 27629 31807
rect 27629 31773 27663 31807
rect 27663 31773 27672 31807
rect 27620 31764 27672 31773
rect 27896 31807 27948 31816
rect 27896 31773 27905 31807
rect 27905 31773 27939 31807
rect 27939 31773 27948 31807
rect 27896 31764 27948 31773
rect 28540 31807 28592 31816
rect 28540 31773 28549 31807
rect 28549 31773 28583 31807
rect 28583 31773 28592 31807
rect 28540 31764 28592 31773
rect 29368 31764 29420 31816
rect 29644 31841 29653 31875
rect 29653 31841 29687 31875
rect 29687 31841 29696 31875
rect 29644 31832 29696 31841
rect 30012 31832 30064 31884
rect 30748 31900 30800 31952
rect 32220 31875 32272 31884
rect 32220 31841 32229 31875
rect 32229 31841 32263 31875
rect 32263 31841 32272 31875
rect 32220 31832 32272 31841
rect 29000 31696 29052 31748
rect 30472 31764 30524 31816
rect 30748 31807 30800 31816
rect 30748 31773 30757 31807
rect 30757 31773 30791 31807
rect 30791 31773 30800 31807
rect 30748 31764 30800 31773
rect 32128 31807 32180 31816
rect 32128 31773 32137 31807
rect 32137 31773 32171 31807
rect 32171 31773 32180 31807
rect 32128 31764 32180 31773
rect 33968 31832 34020 31884
rect 34704 31832 34756 31884
rect 30196 31696 30248 31748
rect 17408 31628 17460 31680
rect 17592 31628 17644 31680
rect 17960 31628 18012 31680
rect 22100 31628 22152 31680
rect 27712 31671 27764 31680
rect 27712 31637 27721 31671
rect 27721 31637 27755 31671
rect 27755 31637 27764 31671
rect 27712 31628 27764 31637
rect 30656 31628 30708 31680
rect 31300 31671 31352 31680
rect 31300 31637 31309 31671
rect 31309 31637 31343 31671
rect 31343 31637 31352 31671
rect 31300 31628 31352 31637
rect 32220 31696 32272 31748
rect 32956 31628 33008 31680
rect 34520 31764 34572 31816
rect 35440 31900 35492 31952
rect 35900 31900 35952 31952
rect 35716 31832 35768 31884
rect 36544 31875 36596 31884
rect 36544 31841 36553 31875
rect 36553 31841 36587 31875
rect 36587 31841 36596 31875
rect 36544 31832 36596 31841
rect 35900 31764 35952 31816
rect 36728 31807 36780 31816
rect 36728 31773 36737 31807
rect 36737 31773 36771 31807
rect 36771 31773 36780 31807
rect 36728 31764 36780 31773
rect 37832 31832 37884 31884
rect 38476 31832 38528 31884
rect 38660 31875 38712 31884
rect 38660 31841 38669 31875
rect 38669 31841 38703 31875
rect 38703 31841 38712 31875
rect 38660 31832 38712 31841
rect 37464 31807 37516 31816
rect 37464 31773 37473 31807
rect 37473 31773 37507 31807
rect 37507 31773 37516 31807
rect 37464 31764 37516 31773
rect 35348 31696 35400 31748
rect 33324 31628 33376 31680
rect 37648 31696 37700 31748
rect 38844 31764 38896 31816
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 12348 31399 12400 31408
rect 12348 31365 12357 31399
rect 12357 31365 12391 31399
rect 12391 31365 12400 31399
rect 12348 31356 12400 31365
rect 13820 31424 13872 31476
rect 15016 31424 15068 31476
rect 15200 31424 15252 31476
rect 16488 31424 16540 31476
rect 17868 31467 17920 31476
rect 17868 31433 17877 31467
rect 17877 31433 17911 31467
rect 17911 31433 17920 31467
rect 17868 31424 17920 31433
rect 12532 31331 12584 31340
rect 12532 31297 12541 31331
rect 12541 31297 12575 31331
rect 12575 31297 12584 31331
rect 12532 31288 12584 31297
rect 13452 31331 13504 31340
rect 13452 31297 13461 31331
rect 13461 31297 13495 31331
rect 13495 31297 13504 31331
rect 13452 31288 13504 31297
rect 13728 31331 13780 31340
rect 13728 31297 13737 31331
rect 13737 31297 13771 31331
rect 13771 31297 13780 31331
rect 13728 31288 13780 31297
rect 14832 31331 14884 31340
rect 14832 31297 14841 31331
rect 14841 31297 14875 31331
rect 14875 31297 14884 31331
rect 14832 31288 14884 31297
rect 15016 31331 15068 31340
rect 15016 31297 15025 31331
rect 15025 31297 15059 31331
rect 15059 31297 15068 31331
rect 15016 31288 15068 31297
rect 15844 31356 15896 31408
rect 14188 31220 14240 31272
rect 15200 31220 15252 31272
rect 17316 31288 17368 31340
rect 17500 31331 17552 31340
rect 17500 31297 17509 31331
rect 17509 31297 17543 31331
rect 17543 31297 17552 31331
rect 17500 31288 17552 31297
rect 18052 31288 18104 31340
rect 19248 31356 19300 31408
rect 19984 31424 20036 31476
rect 21088 31467 21140 31476
rect 21088 31433 21097 31467
rect 21097 31433 21131 31467
rect 21131 31433 21140 31467
rect 21088 31424 21140 31433
rect 23296 31424 23348 31476
rect 24216 31467 24268 31476
rect 24216 31433 24225 31467
rect 24225 31433 24259 31467
rect 24259 31433 24268 31467
rect 24216 31424 24268 31433
rect 24860 31424 24912 31476
rect 24952 31424 25004 31476
rect 26240 31424 26292 31476
rect 27252 31424 27304 31476
rect 27528 31424 27580 31476
rect 27620 31467 27672 31476
rect 27620 31433 27635 31467
rect 27635 31433 27669 31467
rect 27669 31433 27672 31467
rect 27620 31424 27672 31433
rect 27988 31424 28040 31476
rect 29000 31467 29052 31476
rect 29000 31433 29009 31467
rect 29009 31433 29043 31467
rect 29043 31433 29052 31467
rect 29000 31424 29052 31433
rect 29460 31467 29512 31476
rect 29460 31433 29469 31467
rect 29469 31433 29503 31467
rect 29503 31433 29512 31467
rect 29460 31424 29512 31433
rect 30472 31424 30524 31476
rect 32864 31424 32916 31476
rect 34520 31424 34572 31476
rect 35532 31467 35584 31476
rect 35532 31433 35541 31467
rect 35541 31433 35575 31467
rect 35575 31433 35584 31467
rect 35532 31424 35584 31433
rect 37648 31467 37700 31476
rect 37648 31433 37657 31467
rect 37657 31433 37691 31467
rect 37691 31433 37700 31467
rect 37648 31424 37700 31433
rect 38844 31467 38896 31476
rect 38844 31433 38853 31467
rect 38853 31433 38887 31467
rect 38887 31433 38896 31467
rect 38844 31424 38896 31433
rect 39948 31424 40000 31476
rect 18972 31331 19024 31340
rect 18972 31297 18981 31331
rect 18981 31297 19015 31331
rect 19015 31297 19024 31331
rect 18972 31288 19024 31297
rect 19892 31331 19944 31340
rect 19892 31297 19901 31331
rect 19901 31297 19935 31331
rect 19935 31297 19944 31331
rect 19892 31288 19944 31297
rect 21456 31356 21508 31408
rect 22100 31356 22152 31408
rect 22560 31356 22612 31408
rect 20996 31288 21048 31340
rect 22008 31288 22060 31340
rect 22284 31288 22336 31340
rect 25780 31356 25832 31408
rect 26056 31356 26108 31408
rect 26240 31288 26292 31340
rect 27068 31288 27120 31340
rect 27896 31288 27948 31340
rect 29092 31356 29144 31408
rect 28264 31331 28316 31340
rect 28264 31297 28273 31331
rect 28273 31297 28307 31331
rect 28307 31297 28316 31331
rect 28264 31288 28316 31297
rect 28356 31288 28408 31340
rect 29460 31288 29512 31340
rect 30012 31288 30064 31340
rect 31484 31356 31536 31408
rect 33784 31356 33836 31408
rect 30656 31288 30708 31340
rect 31024 31331 31076 31340
rect 31024 31297 31033 31331
rect 31033 31297 31067 31331
rect 31067 31297 31076 31331
rect 31024 31288 31076 31297
rect 31392 31288 31444 31340
rect 32128 31288 32180 31340
rect 32680 31331 32732 31340
rect 20076 31152 20128 31204
rect 28172 31220 28224 31272
rect 28540 31220 28592 31272
rect 31484 31220 31536 31272
rect 32680 31297 32689 31331
rect 32689 31297 32723 31331
rect 32723 31297 32732 31331
rect 32680 31288 32732 31297
rect 32772 31331 32824 31340
rect 32772 31297 32807 31331
rect 32807 31297 32824 31331
rect 32772 31288 32824 31297
rect 33140 31288 33192 31340
rect 33416 31331 33468 31340
rect 33416 31297 33425 31331
rect 33425 31297 33459 31331
rect 33459 31297 33468 31331
rect 33416 31288 33468 31297
rect 35348 31356 35400 31408
rect 38568 31356 38620 31408
rect 33324 31152 33376 31204
rect 12992 31084 13044 31136
rect 16396 31084 16448 31136
rect 16488 31084 16540 31136
rect 19800 31084 19852 31136
rect 19984 31084 20036 31136
rect 20444 31084 20496 31136
rect 22008 31127 22060 31136
rect 22008 31093 22017 31127
rect 22017 31093 22051 31127
rect 22051 31093 22060 31127
rect 22008 31084 22060 31093
rect 25504 31084 25556 31136
rect 27068 31127 27120 31136
rect 27068 31093 27077 31127
rect 27077 31093 27111 31127
rect 27111 31093 27120 31127
rect 27068 31084 27120 31093
rect 29644 31127 29696 31136
rect 29644 31093 29653 31127
rect 29653 31093 29687 31127
rect 29687 31093 29696 31127
rect 29644 31084 29696 31093
rect 31484 31084 31536 31136
rect 37648 31288 37700 31340
rect 37832 31288 37884 31340
rect 34152 31220 34204 31272
rect 35440 31220 35492 31272
rect 36084 31127 36136 31136
rect 36084 31093 36093 31127
rect 36093 31093 36127 31127
rect 36127 31093 36136 31127
rect 36084 31084 36136 31093
rect 36452 31084 36504 31136
rect 37280 31127 37332 31136
rect 37280 31093 37289 31127
rect 37289 31093 37323 31127
rect 37323 31093 37332 31127
rect 37280 31084 37332 31093
rect 38660 31084 38712 31136
rect 38752 31084 38804 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 13728 30880 13780 30932
rect 15200 30923 15252 30932
rect 15200 30889 15209 30923
rect 15209 30889 15243 30923
rect 15243 30889 15252 30923
rect 15200 30880 15252 30889
rect 16856 30880 16908 30932
rect 17408 30923 17460 30932
rect 17408 30889 17417 30923
rect 17417 30889 17451 30923
rect 17451 30889 17460 30923
rect 17408 30880 17460 30889
rect 18696 30923 18748 30932
rect 18696 30889 18705 30923
rect 18705 30889 18739 30923
rect 18739 30889 18748 30923
rect 18696 30880 18748 30889
rect 19984 30923 20036 30932
rect 19984 30889 19993 30923
rect 19993 30889 20027 30923
rect 20027 30889 20036 30923
rect 19984 30880 20036 30889
rect 20076 30880 20128 30932
rect 20996 30880 21048 30932
rect 21456 30880 21508 30932
rect 22376 30923 22428 30932
rect 22376 30889 22385 30923
rect 22385 30889 22419 30923
rect 22419 30889 22428 30923
rect 22376 30880 22428 30889
rect 27712 30880 27764 30932
rect 30012 30880 30064 30932
rect 30748 30923 30800 30932
rect 30748 30889 30757 30923
rect 30757 30889 30791 30923
rect 30791 30889 30800 30923
rect 30748 30880 30800 30889
rect 33140 30880 33192 30932
rect 37096 30923 37148 30932
rect 37096 30889 37105 30923
rect 37105 30889 37139 30923
rect 37139 30889 37148 30923
rect 37096 30880 37148 30889
rect 38016 30880 38068 30932
rect 38752 30923 38804 30932
rect 38752 30889 38761 30923
rect 38761 30889 38795 30923
rect 38795 30889 38804 30923
rect 38752 30880 38804 30889
rect 15568 30812 15620 30864
rect 17316 30812 17368 30864
rect 19800 30812 19852 30864
rect 20444 30812 20496 30864
rect 20536 30812 20588 30864
rect 14832 30744 14884 30796
rect 12348 30719 12400 30728
rect 12348 30685 12357 30719
rect 12357 30685 12391 30719
rect 12391 30685 12400 30719
rect 12348 30676 12400 30685
rect 12532 30719 12584 30728
rect 12532 30685 12541 30719
rect 12541 30685 12575 30719
rect 12575 30685 12584 30719
rect 12532 30676 12584 30685
rect 12992 30719 13044 30728
rect 12992 30685 13001 30719
rect 13001 30685 13035 30719
rect 13035 30685 13044 30719
rect 12992 30676 13044 30685
rect 13268 30676 13320 30728
rect 13820 30608 13872 30660
rect 15292 30608 15344 30660
rect 16856 30676 16908 30728
rect 17500 30744 17552 30796
rect 21180 30744 21232 30796
rect 27252 30812 27304 30864
rect 18052 30676 18104 30728
rect 19432 30676 19484 30728
rect 15844 30608 15896 30660
rect 16028 30608 16080 30660
rect 17316 30608 17368 30660
rect 20352 30608 20404 30660
rect 21272 30676 21324 30728
rect 24308 30744 24360 30796
rect 20628 30651 20680 30660
rect 20076 30540 20128 30592
rect 20628 30617 20653 30651
rect 20653 30617 20680 30651
rect 20628 30608 20680 30617
rect 22100 30608 22152 30660
rect 24124 30676 24176 30728
rect 24492 30676 24544 30728
rect 32680 30744 32732 30796
rect 33232 30744 33284 30796
rect 25964 30676 26016 30728
rect 26792 30719 26844 30728
rect 26792 30685 26801 30719
rect 26801 30685 26835 30719
rect 26835 30685 26844 30719
rect 26792 30676 26844 30685
rect 29460 30676 29512 30728
rect 27528 30608 27580 30660
rect 27896 30651 27948 30660
rect 27896 30617 27905 30651
rect 27905 30617 27939 30651
rect 27939 30617 27948 30651
rect 27896 30608 27948 30617
rect 29276 30608 29328 30660
rect 30656 30676 30708 30728
rect 31392 30676 31444 30728
rect 20996 30540 21048 30592
rect 21732 30540 21784 30592
rect 23756 30583 23808 30592
rect 23756 30549 23765 30583
rect 23765 30549 23799 30583
rect 23799 30549 23808 30583
rect 23756 30540 23808 30549
rect 24032 30540 24084 30592
rect 24768 30540 24820 30592
rect 24860 30540 24912 30592
rect 26240 30540 26292 30592
rect 26516 30540 26568 30592
rect 26976 30540 27028 30592
rect 29000 30583 29052 30592
rect 29000 30549 29009 30583
rect 29009 30549 29043 30583
rect 29043 30549 29052 30583
rect 29000 30540 29052 30549
rect 29184 30540 29236 30592
rect 29552 30540 29604 30592
rect 30104 30540 30156 30592
rect 31024 30608 31076 30660
rect 32220 30676 32272 30728
rect 32956 30719 33008 30728
rect 32956 30685 32965 30719
rect 32965 30685 32999 30719
rect 32999 30685 33008 30719
rect 33508 30719 33560 30728
rect 32956 30676 33008 30685
rect 33508 30685 33517 30719
rect 33517 30685 33551 30719
rect 33551 30685 33560 30719
rect 33508 30676 33560 30685
rect 32036 30608 32088 30660
rect 32496 30608 32548 30660
rect 34704 30608 34756 30660
rect 36452 30676 36504 30728
rect 33232 30540 33284 30592
rect 34060 30540 34112 30592
rect 37096 30608 37148 30660
rect 35900 30540 35952 30592
rect 35992 30583 36044 30592
rect 35992 30549 36001 30583
rect 36001 30549 36035 30583
rect 36035 30549 36044 30583
rect 35992 30540 36044 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 12348 30336 12400 30388
rect 12532 30379 12584 30388
rect 12532 30345 12541 30379
rect 12541 30345 12575 30379
rect 12575 30345 12584 30379
rect 12532 30336 12584 30345
rect 15384 30379 15436 30388
rect 15384 30345 15393 30379
rect 15393 30345 15427 30379
rect 15427 30345 15436 30379
rect 15384 30336 15436 30345
rect 15844 30336 15896 30388
rect 17316 30336 17368 30388
rect 18052 30336 18104 30388
rect 19432 30336 19484 30388
rect 20536 30336 20588 30388
rect 22284 30379 22336 30388
rect 1584 30200 1636 30252
rect 13176 30243 13228 30252
rect 13176 30209 13185 30243
rect 13185 30209 13219 30243
rect 13219 30209 13228 30243
rect 13176 30200 13228 30209
rect 15292 30243 15344 30252
rect 15292 30209 15301 30243
rect 15301 30209 15335 30243
rect 15335 30209 15344 30243
rect 15292 30200 15344 30209
rect 15568 30243 15620 30252
rect 15568 30209 15577 30243
rect 15577 30209 15611 30243
rect 15611 30209 15620 30243
rect 15568 30200 15620 30209
rect 16304 30200 16356 30252
rect 16672 30243 16724 30252
rect 16672 30209 16681 30243
rect 16681 30209 16715 30243
rect 16715 30209 16724 30243
rect 16672 30200 16724 30209
rect 16580 30132 16632 30184
rect 16948 30243 17000 30252
rect 16948 30209 16957 30243
rect 16957 30209 16991 30243
rect 16991 30209 17000 30243
rect 16948 30200 17000 30209
rect 21180 30268 21232 30320
rect 22284 30345 22293 30379
rect 22293 30345 22327 30379
rect 22327 30345 22336 30379
rect 22284 30336 22336 30345
rect 24768 30336 24820 30388
rect 27436 30268 27488 30320
rect 29092 30336 29144 30388
rect 19248 30200 19300 30252
rect 19524 30243 19576 30252
rect 19524 30209 19533 30243
rect 19533 30209 19567 30243
rect 19567 30209 19576 30243
rect 19524 30200 19576 30209
rect 19340 30132 19392 30184
rect 17776 29996 17828 30048
rect 17960 30039 18012 30048
rect 17960 30005 17969 30039
rect 17969 30005 18003 30039
rect 18003 30005 18012 30039
rect 17960 29996 18012 30005
rect 19432 30064 19484 30116
rect 20628 30200 20680 30252
rect 20076 30132 20128 30184
rect 20996 30243 21048 30252
rect 20996 30209 21005 30243
rect 21005 30209 21039 30243
rect 21039 30209 21048 30243
rect 20996 30200 21048 30209
rect 21272 30243 21324 30252
rect 21272 30209 21281 30243
rect 21281 30209 21315 30243
rect 21315 30209 21324 30243
rect 23020 30243 23072 30252
rect 21272 30200 21324 30209
rect 23020 30209 23029 30243
rect 23029 30209 23063 30243
rect 23063 30209 23072 30243
rect 23020 30200 23072 30209
rect 24032 30243 24084 30252
rect 24032 30209 24041 30243
rect 24041 30209 24075 30243
rect 24075 30209 24084 30243
rect 24032 30200 24084 30209
rect 23940 30175 23992 30184
rect 23940 30141 23949 30175
rect 23949 30141 23983 30175
rect 23983 30141 23992 30175
rect 25136 30243 25188 30252
rect 24400 30175 24452 30184
rect 23940 30132 23992 30141
rect 24400 30141 24409 30175
rect 24409 30141 24443 30175
rect 24443 30141 24452 30175
rect 24400 30132 24452 30141
rect 25136 30209 25145 30243
rect 25145 30209 25179 30243
rect 25179 30209 25188 30243
rect 25136 30200 25188 30209
rect 25780 30243 25832 30252
rect 25780 30209 25789 30243
rect 25789 30209 25823 30243
rect 25823 30209 25832 30243
rect 25780 30200 25832 30209
rect 26884 30200 26936 30252
rect 26792 30064 26844 30116
rect 28356 30243 28408 30252
rect 28356 30209 28365 30243
rect 28365 30209 28399 30243
rect 28399 30209 28408 30243
rect 28540 30243 28592 30252
rect 28356 30200 28408 30209
rect 28540 30209 28549 30243
rect 28549 30209 28583 30243
rect 28583 30209 28592 30243
rect 28540 30200 28592 30209
rect 28816 30268 28868 30320
rect 29092 30243 29144 30252
rect 29092 30209 29101 30243
rect 29101 30209 29135 30243
rect 29135 30209 29144 30243
rect 29092 30200 29144 30209
rect 29644 30200 29696 30252
rect 29920 30200 29972 30252
rect 29552 30175 29604 30184
rect 29552 30141 29561 30175
rect 29561 30141 29595 30175
rect 29595 30141 29604 30175
rect 29552 30132 29604 30141
rect 30196 30132 30248 30184
rect 31392 30243 31444 30252
rect 31392 30209 31401 30243
rect 31401 30209 31435 30243
rect 31435 30209 31444 30243
rect 31392 30200 31444 30209
rect 32772 30336 32824 30388
rect 35716 30336 35768 30388
rect 37096 30336 37148 30388
rect 38660 30336 38712 30388
rect 39396 30336 39448 30388
rect 32956 30268 33008 30320
rect 32220 30243 32272 30252
rect 31484 30132 31536 30184
rect 32220 30209 32229 30243
rect 32229 30209 32263 30243
rect 32263 30209 32272 30243
rect 32220 30200 32272 30209
rect 32496 30243 32548 30252
rect 32496 30209 32505 30243
rect 32505 30209 32539 30243
rect 32539 30209 32548 30243
rect 32496 30200 32548 30209
rect 33140 30200 33192 30252
rect 33600 30243 33652 30252
rect 33600 30209 33609 30243
rect 33609 30209 33643 30243
rect 33643 30209 33652 30243
rect 33600 30200 33652 30209
rect 34060 30243 34112 30252
rect 34060 30209 34069 30243
rect 34069 30209 34103 30243
rect 34103 30209 34112 30243
rect 34060 30200 34112 30209
rect 34152 30132 34204 30184
rect 34704 30200 34756 30252
rect 35256 30200 35308 30252
rect 36544 30200 36596 30252
rect 34796 30175 34848 30184
rect 34796 30141 34805 30175
rect 34805 30141 34839 30175
rect 34839 30141 34848 30175
rect 34796 30132 34848 30141
rect 37280 30200 37332 30252
rect 39488 30132 39540 30184
rect 20628 29996 20680 30048
rect 25228 29996 25280 30048
rect 26240 29996 26292 30048
rect 27068 29996 27120 30048
rect 27620 30039 27672 30048
rect 27620 30005 27629 30039
rect 27629 30005 27663 30039
rect 27663 30005 27672 30039
rect 27620 29996 27672 30005
rect 27804 29996 27856 30048
rect 28816 29996 28868 30048
rect 29552 29996 29604 30048
rect 29828 29996 29880 30048
rect 31484 29996 31536 30048
rect 33324 29996 33376 30048
rect 33692 29996 33744 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 1584 29835 1636 29844
rect 1584 29801 1593 29835
rect 1593 29801 1627 29835
rect 1627 29801 1636 29835
rect 1584 29792 1636 29801
rect 15384 29792 15436 29844
rect 16028 29835 16080 29844
rect 16028 29801 16037 29835
rect 16037 29801 16071 29835
rect 16071 29801 16080 29835
rect 16028 29792 16080 29801
rect 16948 29835 17000 29844
rect 15292 29724 15344 29776
rect 16948 29801 16957 29835
rect 16957 29801 16991 29835
rect 16991 29801 17000 29835
rect 16948 29792 17000 29801
rect 17776 29835 17828 29844
rect 17776 29801 17785 29835
rect 17785 29801 17819 29835
rect 17819 29801 17828 29835
rect 17776 29792 17828 29801
rect 16304 29724 16356 29776
rect 18972 29792 19024 29844
rect 20076 29792 20128 29844
rect 21180 29835 21232 29844
rect 21180 29801 21189 29835
rect 21189 29801 21223 29835
rect 21223 29801 21232 29835
rect 21180 29792 21232 29801
rect 22836 29835 22888 29844
rect 22836 29801 22845 29835
rect 22845 29801 22879 29835
rect 22879 29801 22888 29835
rect 22836 29792 22888 29801
rect 25136 29792 25188 29844
rect 19340 29724 19392 29776
rect 16488 29656 16540 29708
rect 25872 29724 25924 29776
rect 26792 29792 26844 29844
rect 27896 29792 27948 29844
rect 28908 29835 28960 29844
rect 28908 29801 28917 29835
rect 28917 29801 28951 29835
rect 28951 29801 28960 29835
rect 28908 29792 28960 29801
rect 29736 29792 29788 29844
rect 30472 29835 30524 29844
rect 30472 29801 30481 29835
rect 30481 29801 30515 29835
rect 30515 29801 30524 29835
rect 30472 29792 30524 29801
rect 30564 29792 30616 29844
rect 33508 29792 33560 29844
rect 34244 29792 34296 29844
rect 20536 29656 20588 29708
rect 16856 29631 16908 29640
rect 16856 29597 16865 29631
rect 16865 29597 16899 29631
rect 16899 29597 16908 29631
rect 16856 29588 16908 29597
rect 17040 29631 17092 29640
rect 17040 29597 17049 29631
rect 17049 29597 17083 29631
rect 17083 29597 17092 29631
rect 17040 29588 17092 29597
rect 18604 29588 18656 29640
rect 19340 29631 19392 29640
rect 19340 29597 19349 29631
rect 19349 29597 19383 29631
rect 19383 29597 19392 29631
rect 19340 29588 19392 29597
rect 19524 29588 19576 29640
rect 20076 29588 20128 29640
rect 20168 29588 20220 29640
rect 20628 29631 20680 29640
rect 20628 29597 20637 29631
rect 20637 29597 20671 29631
rect 20671 29597 20680 29631
rect 20628 29588 20680 29597
rect 20996 29588 21048 29640
rect 22284 29656 22336 29708
rect 22744 29656 22796 29708
rect 22836 29656 22888 29708
rect 23296 29656 23348 29708
rect 25228 29699 25280 29708
rect 22008 29631 22060 29640
rect 16580 29520 16632 29572
rect 17684 29520 17736 29572
rect 19156 29520 19208 29572
rect 22008 29597 22017 29631
rect 22017 29597 22051 29631
rect 22051 29597 22060 29631
rect 22008 29588 22060 29597
rect 25228 29665 25237 29699
rect 25237 29665 25271 29699
rect 25271 29665 25280 29699
rect 25228 29656 25280 29665
rect 26424 29656 26476 29708
rect 27528 29656 27580 29708
rect 27620 29656 27672 29708
rect 22376 29520 22428 29572
rect 23756 29631 23808 29640
rect 23756 29597 23765 29631
rect 23765 29597 23799 29631
rect 23799 29597 23808 29631
rect 23756 29588 23808 29597
rect 25044 29588 25096 29640
rect 25780 29588 25832 29640
rect 25964 29588 26016 29640
rect 26884 29588 26936 29640
rect 27160 29588 27212 29640
rect 28356 29631 28408 29640
rect 28356 29597 28365 29631
rect 28365 29597 28399 29631
rect 28399 29597 28408 29631
rect 28356 29588 28408 29597
rect 29368 29588 29420 29640
rect 29552 29631 29604 29640
rect 29552 29597 29561 29631
rect 29561 29597 29595 29631
rect 29595 29597 29604 29631
rect 29552 29588 29604 29597
rect 29828 29631 29880 29640
rect 29828 29597 29837 29631
rect 29837 29597 29871 29631
rect 29871 29597 29880 29631
rect 29828 29588 29880 29597
rect 31392 29724 31444 29776
rect 31484 29631 31536 29640
rect 31484 29597 31493 29631
rect 31493 29597 31527 29631
rect 31527 29597 31536 29631
rect 31484 29588 31536 29597
rect 24492 29520 24544 29572
rect 15476 29495 15528 29504
rect 15476 29461 15485 29495
rect 15485 29461 15519 29495
rect 15519 29461 15528 29495
rect 15476 29452 15528 29461
rect 18420 29452 18472 29504
rect 19432 29495 19484 29504
rect 19432 29461 19441 29495
rect 19441 29461 19475 29495
rect 19475 29461 19484 29495
rect 19432 29452 19484 29461
rect 20260 29495 20312 29504
rect 20260 29461 20269 29495
rect 20269 29461 20303 29495
rect 20303 29461 20312 29495
rect 20260 29452 20312 29461
rect 21916 29495 21968 29504
rect 21916 29461 21925 29495
rect 21925 29461 21959 29495
rect 21959 29461 21968 29495
rect 21916 29452 21968 29461
rect 22560 29452 22612 29504
rect 23664 29495 23716 29504
rect 23664 29461 23666 29495
rect 23666 29461 23700 29495
rect 23700 29461 23716 29495
rect 23664 29452 23716 29461
rect 24860 29452 24912 29504
rect 25688 29452 25740 29504
rect 33140 29699 33192 29708
rect 33140 29665 33149 29699
rect 33149 29665 33183 29699
rect 33183 29665 33192 29699
rect 33140 29656 33192 29665
rect 33324 29724 33376 29776
rect 35992 29792 36044 29844
rect 37464 29792 37516 29844
rect 35348 29767 35400 29776
rect 35348 29733 35357 29767
rect 35357 29733 35391 29767
rect 35391 29733 35400 29767
rect 35348 29724 35400 29733
rect 34244 29656 34296 29708
rect 35900 29699 35952 29708
rect 35900 29665 35909 29699
rect 35909 29665 35943 29699
rect 35943 29665 35952 29699
rect 48136 29699 48188 29708
rect 35900 29656 35952 29665
rect 32496 29631 32548 29640
rect 32496 29597 32505 29631
rect 32505 29597 32539 29631
rect 32539 29597 32548 29631
rect 32496 29588 32548 29597
rect 32680 29631 32732 29640
rect 32680 29597 32689 29631
rect 32689 29597 32723 29631
rect 32723 29597 32732 29631
rect 32680 29588 32732 29597
rect 33600 29631 33652 29640
rect 33600 29597 33609 29631
rect 33609 29597 33643 29631
rect 33643 29597 33652 29631
rect 33600 29588 33652 29597
rect 33692 29588 33744 29640
rect 35808 29631 35860 29640
rect 35808 29597 35817 29631
rect 35817 29597 35851 29631
rect 35851 29597 35860 29631
rect 35808 29588 35860 29597
rect 48136 29665 48145 29699
rect 48145 29665 48179 29699
rect 48179 29665 48188 29699
rect 48136 29656 48188 29665
rect 34612 29520 34664 29572
rect 46388 29588 46440 29640
rect 28264 29452 28316 29504
rect 29644 29452 29696 29504
rect 30932 29452 30984 29504
rect 32036 29495 32088 29504
rect 32036 29461 32045 29495
rect 32045 29461 32079 29495
rect 32079 29461 32088 29495
rect 32036 29452 32088 29461
rect 33416 29495 33468 29504
rect 33416 29461 33425 29495
rect 33425 29461 33459 29495
rect 33459 29461 33468 29495
rect 33416 29452 33468 29461
rect 33692 29452 33744 29504
rect 36544 29495 36596 29504
rect 36544 29461 36553 29495
rect 36553 29461 36587 29495
rect 36587 29461 36596 29495
rect 36544 29452 36596 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 16856 29248 16908 29300
rect 17040 29291 17092 29300
rect 17040 29257 17049 29291
rect 17049 29257 17083 29291
rect 17083 29257 17092 29291
rect 17040 29248 17092 29257
rect 17684 29291 17736 29300
rect 17684 29257 17693 29291
rect 17693 29257 17727 29291
rect 17727 29257 17736 29291
rect 17684 29248 17736 29257
rect 18880 29291 18932 29300
rect 18880 29257 18889 29291
rect 18889 29257 18923 29291
rect 18923 29257 18932 29291
rect 18880 29248 18932 29257
rect 19340 29248 19392 29300
rect 20996 29291 21048 29300
rect 20996 29257 21005 29291
rect 21005 29257 21039 29291
rect 21039 29257 21048 29291
rect 20996 29248 21048 29257
rect 22560 29291 22612 29300
rect 22560 29257 22569 29291
rect 22569 29257 22603 29291
rect 22603 29257 22612 29291
rect 22560 29248 22612 29257
rect 23296 29291 23348 29300
rect 23296 29257 23305 29291
rect 23305 29257 23339 29291
rect 23339 29257 23348 29291
rect 23296 29248 23348 29257
rect 23940 29248 23992 29300
rect 24768 29248 24820 29300
rect 27620 29248 27672 29300
rect 28264 29291 28316 29300
rect 28264 29257 28273 29291
rect 28273 29257 28307 29291
rect 28307 29257 28316 29291
rect 28264 29248 28316 29257
rect 28724 29248 28776 29300
rect 30472 29291 30524 29300
rect 30472 29257 30481 29291
rect 30481 29257 30515 29291
rect 30515 29257 30524 29291
rect 30472 29248 30524 29257
rect 30932 29291 30984 29300
rect 30932 29257 30941 29291
rect 30941 29257 30975 29291
rect 30975 29257 30984 29291
rect 30932 29248 30984 29257
rect 33140 29248 33192 29300
rect 34796 29248 34848 29300
rect 35808 29291 35860 29300
rect 35808 29257 35817 29291
rect 35817 29257 35851 29291
rect 35851 29257 35860 29291
rect 35808 29248 35860 29257
rect 48136 29291 48188 29300
rect 48136 29257 48145 29291
rect 48145 29257 48179 29291
rect 48179 29257 48188 29291
rect 48136 29248 48188 29257
rect 18420 29180 18472 29232
rect 20628 29223 20680 29232
rect 14832 29019 14884 29028
rect 14832 28985 14841 29019
rect 14841 28985 14875 29019
rect 14875 28985 14884 29019
rect 16120 29155 16172 29164
rect 16120 29121 16129 29155
rect 16129 29121 16163 29155
rect 16163 29121 16172 29155
rect 16120 29112 16172 29121
rect 17224 29112 17276 29164
rect 17592 29155 17644 29164
rect 17592 29121 17601 29155
rect 17601 29121 17635 29155
rect 17635 29121 17644 29155
rect 17592 29112 17644 29121
rect 17960 29155 18012 29164
rect 17960 29121 17969 29155
rect 17969 29121 18003 29155
rect 18003 29121 18012 29155
rect 17960 29112 18012 29121
rect 18788 29155 18840 29164
rect 18788 29121 18797 29155
rect 18797 29121 18831 29155
rect 18831 29121 18840 29155
rect 18788 29112 18840 29121
rect 19064 29155 19116 29164
rect 19064 29121 19073 29155
rect 19073 29121 19107 29155
rect 19107 29121 19116 29155
rect 19064 29112 19116 29121
rect 19156 29112 19208 29164
rect 19524 29112 19576 29164
rect 20628 29189 20637 29223
rect 20637 29189 20671 29223
rect 20671 29189 20680 29223
rect 20628 29180 20680 29189
rect 21088 29180 21140 29232
rect 19800 29112 19852 29164
rect 22008 29112 22060 29164
rect 23020 29155 23072 29164
rect 18236 29044 18288 29096
rect 14832 28976 14884 28985
rect 15476 28976 15528 29028
rect 16948 28976 17000 29028
rect 17776 28976 17828 29028
rect 20076 29044 20128 29096
rect 22100 29044 22152 29096
rect 23020 29121 23029 29155
rect 23029 29121 23063 29155
rect 23063 29121 23072 29155
rect 23020 29112 23072 29121
rect 23664 29112 23716 29164
rect 24492 29155 24544 29164
rect 24492 29121 24501 29155
rect 24501 29121 24535 29155
rect 24535 29121 24544 29155
rect 24492 29112 24544 29121
rect 24676 29112 24728 29164
rect 25136 29112 25188 29164
rect 29736 29180 29788 29232
rect 32496 29180 32548 29232
rect 33968 29180 34020 29232
rect 25688 29155 25740 29164
rect 25688 29121 25697 29155
rect 25697 29121 25731 29155
rect 25731 29121 25740 29155
rect 26976 29155 27028 29164
rect 25688 29112 25740 29121
rect 26976 29121 26985 29155
rect 26985 29121 27019 29155
rect 27019 29121 27028 29155
rect 26976 29112 27028 29121
rect 27988 29112 28040 29164
rect 28172 29155 28224 29164
rect 28172 29121 28181 29155
rect 28181 29121 28215 29155
rect 28215 29121 28224 29155
rect 29368 29155 29420 29164
rect 28172 29112 28224 29121
rect 29368 29121 29377 29155
rect 29377 29121 29411 29155
rect 29411 29121 29420 29155
rect 29368 29112 29420 29121
rect 29920 29112 29972 29164
rect 30104 29155 30156 29164
rect 30104 29121 30113 29155
rect 30113 29121 30147 29155
rect 30147 29121 30156 29155
rect 30104 29112 30156 29121
rect 30196 29155 30248 29164
rect 30196 29121 30205 29155
rect 30205 29121 30239 29155
rect 30239 29121 30248 29155
rect 30196 29112 30248 29121
rect 32680 29112 32732 29164
rect 26332 29044 26384 29096
rect 19984 28951 20036 28960
rect 19984 28917 19993 28951
rect 19993 28917 20027 28951
rect 20027 28917 20036 28951
rect 27896 29019 27948 29028
rect 27896 28985 27905 29019
rect 27905 28985 27939 29019
rect 27939 28985 27948 29019
rect 27896 28976 27948 28985
rect 19984 28908 20036 28917
rect 20536 28908 20588 28960
rect 22376 28951 22428 28960
rect 22376 28917 22385 28951
rect 22385 28917 22419 28951
rect 22419 28917 22428 28951
rect 22376 28908 22428 28917
rect 22928 28908 22980 28960
rect 24860 28908 24912 28960
rect 25688 28908 25740 28960
rect 26516 28908 26568 28960
rect 36544 29112 36596 29164
rect 33416 29044 33468 29096
rect 34336 28976 34388 29028
rect 34520 29087 34572 29096
rect 34520 29053 34529 29087
rect 34529 29053 34563 29087
rect 34563 29053 34572 29087
rect 34520 29044 34572 29053
rect 37280 29044 37332 29096
rect 31944 28908 31996 28960
rect 34796 28908 34848 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 15384 28704 15436 28756
rect 18328 28704 18380 28756
rect 18880 28704 18932 28756
rect 19064 28704 19116 28756
rect 20444 28704 20496 28756
rect 23480 28704 23532 28756
rect 24216 28704 24268 28756
rect 25044 28747 25096 28756
rect 25044 28713 25053 28747
rect 25053 28713 25087 28747
rect 25087 28713 25096 28747
rect 25044 28704 25096 28713
rect 26332 28747 26384 28756
rect 26332 28713 26341 28747
rect 26341 28713 26375 28747
rect 26375 28713 26384 28747
rect 26332 28704 26384 28713
rect 17776 28636 17828 28688
rect 20352 28636 20404 28688
rect 22928 28636 22980 28688
rect 28172 28704 28224 28756
rect 29644 28747 29696 28756
rect 29644 28713 29653 28747
rect 29653 28713 29687 28747
rect 29687 28713 29696 28747
rect 29644 28704 29696 28713
rect 30196 28704 30248 28756
rect 20536 28611 20588 28620
rect 20536 28577 20545 28611
rect 20545 28577 20579 28611
rect 20579 28577 20588 28611
rect 20536 28568 20588 28577
rect 21088 28611 21140 28620
rect 21088 28577 21097 28611
rect 21097 28577 21131 28611
rect 21131 28577 21140 28611
rect 21088 28568 21140 28577
rect 22744 28568 22796 28620
rect 24584 28611 24636 28620
rect 24584 28577 24593 28611
rect 24593 28577 24627 28611
rect 24627 28577 24636 28611
rect 24584 28568 24636 28577
rect 27896 28611 27948 28620
rect 27896 28577 27905 28611
rect 27905 28577 27939 28611
rect 27939 28577 27948 28611
rect 27896 28568 27948 28577
rect 28264 28568 28316 28620
rect 29368 28568 29420 28620
rect 16672 28500 16724 28552
rect 17592 28543 17644 28552
rect 17592 28509 17601 28543
rect 17601 28509 17635 28543
rect 17635 28509 17644 28543
rect 17592 28500 17644 28509
rect 17684 28543 17736 28552
rect 17684 28509 17693 28543
rect 17693 28509 17727 28543
rect 17727 28509 17736 28543
rect 17684 28500 17736 28509
rect 17960 28500 18012 28552
rect 19340 28543 19392 28552
rect 19340 28509 19349 28543
rect 19349 28509 19383 28543
rect 19383 28509 19392 28543
rect 19340 28500 19392 28509
rect 20260 28500 20312 28552
rect 20628 28500 20680 28552
rect 21916 28500 21968 28552
rect 23112 28500 23164 28552
rect 24860 28500 24912 28552
rect 22100 28432 22152 28484
rect 23020 28432 23072 28484
rect 15752 28407 15804 28416
rect 15752 28373 15761 28407
rect 15761 28373 15795 28407
rect 15795 28373 15804 28407
rect 15752 28364 15804 28373
rect 16120 28364 16172 28416
rect 17960 28364 18012 28416
rect 26332 28543 26384 28552
rect 26332 28509 26341 28543
rect 26341 28509 26375 28543
rect 26375 28509 26384 28543
rect 26332 28500 26384 28509
rect 27160 28500 27212 28552
rect 27988 28543 28040 28552
rect 27988 28509 27997 28543
rect 27997 28509 28031 28543
rect 28031 28509 28040 28543
rect 27988 28500 28040 28509
rect 30380 28568 30432 28620
rect 32036 28636 32088 28688
rect 34520 28704 34572 28756
rect 29736 28543 29788 28552
rect 29736 28509 29745 28543
rect 29745 28509 29779 28543
rect 29779 28509 29788 28543
rect 29736 28500 29788 28509
rect 30196 28500 30248 28552
rect 31852 28543 31904 28552
rect 26792 28475 26844 28484
rect 26792 28441 26801 28475
rect 26801 28441 26835 28475
rect 26835 28441 26844 28475
rect 26792 28432 26844 28441
rect 27068 28432 27120 28484
rect 31852 28509 31861 28543
rect 31861 28509 31895 28543
rect 31895 28509 31904 28543
rect 31852 28500 31904 28509
rect 34612 28636 34664 28688
rect 35440 28636 35492 28688
rect 34796 28611 34848 28620
rect 32496 28500 32548 28552
rect 33416 28500 33468 28552
rect 32312 28432 32364 28484
rect 26884 28364 26936 28416
rect 28816 28407 28868 28416
rect 28816 28373 28825 28407
rect 28825 28373 28859 28407
rect 28859 28373 28868 28407
rect 28816 28364 28868 28373
rect 29460 28364 29512 28416
rect 31024 28364 31076 28416
rect 34796 28577 34805 28611
rect 34805 28577 34839 28611
rect 34839 28577 34848 28611
rect 34796 28568 34848 28577
rect 34060 28500 34112 28552
rect 35348 28500 35400 28552
rect 45284 28364 45336 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 18420 28203 18472 28212
rect 18420 28169 18429 28203
rect 18429 28169 18463 28203
rect 18463 28169 18472 28203
rect 18420 28160 18472 28169
rect 20628 28160 20680 28212
rect 18328 28135 18380 28144
rect 18328 28101 18337 28135
rect 18337 28101 18371 28135
rect 18371 28101 18380 28135
rect 18328 28092 18380 28101
rect 18788 28092 18840 28144
rect 27068 28160 27120 28212
rect 27896 28160 27948 28212
rect 29736 28160 29788 28212
rect 29920 28160 29972 28212
rect 31852 28160 31904 28212
rect 32220 28203 32272 28212
rect 32220 28169 32229 28203
rect 32229 28169 32263 28203
rect 32263 28169 32272 28203
rect 32220 28160 32272 28169
rect 32496 28160 32548 28212
rect 18236 28067 18288 28076
rect 1492 27931 1544 27940
rect 1492 27897 1501 27931
rect 1501 27897 1535 27931
rect 1535 27897 1544 27931
rect 1492 27888 1544 27897
rect 18236 28033 18245 28067
rect 18245 28033 18279 28067
rect 18279 28033 18288 28067
rect 18236 28024 18288 28033
rect 15292 27956 15344 28008
rect 19708 28067 19760 28076
rect 19708 28033 19717 28067
rect 19717 28033 19751 28067
rect 19751 28033 19760 28067
rect 19708 28024 19760 28033
rect 19892 28024 19944 28076
rect 22284 28067 22336 28076
rect 22284 28033 22293 28067
rect 22293 28033 22327 28067
rect 22327 28033 22336 28067
rect 22284 28024 22336 28033
rect 23480 28092 23532 28144
rect 26056 28135 26108 28144
rect 26056 28101 26065 28135
rect 26065 28101 26099 28135
rect 26099 28101 26108 28135
rect 26056 28092 26108 28101
rect 24768 28024 24820 28076
rect 25964 28067 26016 28076
rect 25964 28033 25973 28067
rect 25973 28033 26007 28067
rect 26007 28033 26016 28067
rect 25964 28024 26016 28033
rect 26516 28024 26568 28076
rect 31944 28092 31996 28144
rect 32128 28092 32180 28144
rect 34612 28160 34664 28212
rect 34520 28135 34572 28144
rect 34520 28101 34529 28135
rect 34529 28101 34563 28135
rect 34563 28101 34572 28135
rect 37556 28160 37608 28212
rect 34520 28092 34572 28101
rect 28816 28024 28868 28076
rect 30196 28067 30248 28076
rect 30196 28033 30205 28067
rect 30205 28033 30239 28067
rect 30239 28033 30248 28067
rect 30196 28024 30248 28033
rect 30380 28067 30432 28076
rect 30380 28033 30389 28067
rect 30389 28033 30423 28067
rect 30423 28033 30432 28067
rect 30380 28024 30432 28033
rect 30840 28067 30892 28076
rect 30840 28033 30849 28067
rect 30849 28033 30883 28067
rect 30883 28033 30892 28067
rect 30840 28024 30892 28033
rect 31024 28067 31076 28076
rect 31024 28033 31033 28067
rect 31033 28033 31067 28067
rect 31067 28033 31076 28067
rect 31024 28024 31076 28033
rect 32864 28067 32916 28076
rect 32864 28033 32873 28067
rect 32873 28033 32907 28067
rect 32907 28033 32916 28067
rect 32864 28024 32916 28033
rect 33508 28024 33560 28076
rect 34060 28067 34112 28076
rect 34060 28033 34069 28067
rect 34069 28033 34103 28067
rect 34103 28033 34112 28067
rect 34060 28024 34112 28033
rect 23480 27999 23532 28008
rect 23480 27965 23489 27999
rect 23489 27965 23523 27999
rect 23523 27965 23532 27999
rect 23480 27956 23532 27965
rect 25228 27956 25280 28008
rect 27712 27999 27764 28008
rect 27712 27965 27721 27999
rect 27721 27965 27755 27999
rect 27755 27965 27764 27999
rect 27712 27956 27764 27965
rect 17960 27888 18012 27940
rect 19248 27888 19300 27940
rect 19432 27931 19484 27940
rect 19432 27897 19441 27931
rect 19441 27897 19475 27931
rect 19475 27897 19484 27931
rect 19432 27888 19484 27897
rect 24860 27888 24912 27940
rect 25504 27888 25556 27940
rect 26792 27888 26844 27940
rect 18604 27820 18656 27872
rect 19340 27820 19392 27872
rect 23572 27820 23624 27872
rect 24952 27863 25004 27872
rect 24952 27829 24961 27863
rect 24961 27829 24995 27863
rect 24995 27829 25004 27863
rect 24952 27820 25004 27829
rect 28816 27820 28868 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 19432 27616 19484 27668
rect 20076 27616 20128 27668
rect 22100 27616 22152 27668
rect 26056 27616 26108 27668
rect 27160 27616 27212 27668
rect 27988 27616 28040 27668
rect 30840 27616 30892 27668
rect 32864 27616 32916 27668
rect 18604 27591 18656 27600
rect 18604 27557 18613 27591
rect 18613 27557 18647 27591
rect 18647 27557 18656 27591
rect 18604 27548 18656 27557
rect 20996 27591 21048 27600
rect 20996 27557 21005 27591
rect 21005 27557 21039 27591
rect 21039 27557 21048 27591
rect 20996 27548 21048 27557
rect 22192 27548 22244 27600
rect 24952 27548 25004 27600
rect 33508 27591 33560 27600
rect 33508 27557 33517 27591
rect 33517 27557 33551 27591
rect 33551 27557 33560 27591
rect 33508 27548 33560 27557
rect 33600 27548 33652 27600
rect 46388 27548 46440 27600
rect 19708 27455 19760 27464
rect 19708 27421 19717 27455
rect 19717 27421 19751 27455
rect 19751 27421 19760 27455
rect 19708 27412 19760 27421
rect 19892 27455 19944 27464
rect 19892 27421 19901 27455
rect 19901 27421 19935 27455
rect 19935 27421 19944 27455
rect 19892 27412 19944 27421
rect 21548 27455 21600 27464
rect 21548 27421 21557 27455
rect 21557 27421 21591 27455
rect 21591 27421 21600 27455
rect 21548 27412 21600 27421
rect 22284 27412 22336 27464
rect 34796 27480 34848 27532
rect 48136 27523 48188 27532
rect 48136 27489 48145 27523
rect 48145 27489 48179 27523
rect 48179 27489 48188 27523
rect 48136 27480 48188 27489
rect 20168 27344 20220 27396
rect 22928 27412 22980 27464
rect 23572 27455 23624 27464
rect 23572 27421 23581 27455
rect 23581 27421 23615 27455
rect 23615 27421 23624 27455
rect 23572 27412 23624 27421
rect 24768 27412 24820 27464
rect 25136 27455 25188 27464
rect 25136 27421 25145 27455
rect 25145 27421 25179 27455
rect 25179 27421 25188 27455
rect 25136 27412 25188 27421
rect 26240 27412 26292 27464
rect 23020 27344 23072 27396
rect 26516 27344 26568 27396
rect 27160 27412 27212 27464
rect 20536 27319 20588 27328
rect 20536 27285 20545 27319
rect 20545 27285 20579 27319
rect 20579 27285 20588 27319
rect 20536 27276 20588 27285
rect 24952 27319 25004 27328
rect 24952 27285 24961 27319
rect 24961 27285 24995 27319
rect 24995 27285 25004 27319
rect 24952 27276 25004 27285
rect 25964 27276 26016 27328
rect 27160 27319 27212 27328
rect 27160 27285 27169 27319
rect 27169 27285 27203 27319
rect 27203 27285 27212 27319
rect 27160 27276 27212 27285
rect 27344 27276 27396 27328
rect 27436 27276 27488 27328
rect 29000 27412 29052 27464
rect 30840 27412 30892 27464
rect 31116 27412 31168 27464
rect 32128 27455 32180 27464
rect 32128 27421 32137 27455
rect 32137 27421 32171 27455
rect 32171 27421 32180 27455
rect 32128 27412 32180 27421
rect 30656 27344 30708 27396
rect 31024 27387 31076 27396
rect 31024 27353 31033 27387
rect 31033 27353 31067 27387
rect 31067 27353 31076 27387
rect 31024 27344 31076 27353
rect 32036 27344 32088 27396
rect 32496 27412 32548 27464
rect 34060 27412 34112 27464
rect 36544 27412 36596 27464
rect 32312 27276 32364 27328
rect 33968 27319 34020 27328
rect 33968 27285 33977 27319
rect 33977 27285 34011 27319
rect 34011 27285 34020 27319
rect 33968 27276 34020 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 18604 27072 18656 27124
rect 19984 27072 20036 27124
rect 19616 27004 19668 27056
rect 20352 27047 20404 27056
rect 20352 27013 20361 27047
rect 20361 27013 20395 27047
rect 20395 27013 20404 27047
rect 20352 27004 20404 27013
rect 21824 27072 21876 27124
rect 22008 27072 22060 27124
rect 24584 27072 24636 27124
rect 24768 27072 24820 27124
rect 21548 27004 21600 27056
rect 20536 26979 20588 26988
rect 20536 26945 20545 26979
rect 20545 26945 20579 26979
rect 20579 26945 20588 26979
rect 20536 26936 20588 26945
rect 21088 26979 21140 26988
rect 21088 26945 21097 26979
rect 21097 26945 21131 26979
rect 21131 26945 21140 26979
rect 21088 26936 21140 26945
rect 25228 27004 25280 27056
rect 23020 26979 23072 26988
rect 23020 26945 23029 26979
rect 23029 26945 23063 26979
rect 23063 26945 23072 26979
rect 23020 26936 23072 26945
rect 24032 26979 24084 26988
rect 24032 26945 24041 26979
rect 24041 26945 24075 26979
rect 24075 26945 24084 26979
rect 24032 26936 24084 26945
rect 22284 26911 22336 26920
rect 22284 26877 22293 26911
rect 22293 26877 22327 26911
rect 22327 26877 22336 26911
rect 22284 26868 22336 26877
rect 23112 26911 23164 26920
rect 23112 26877 23121 26911
rect 23121 26877 23155 26911
rect 23155 26877 23164 26911
rect 23112 26868 23164 26877
rect 24768 26936 24820 26988
rect 24952 26936 25004 26988
rect 25044 26936 25096 26988
rect 25964 27072 26016 27124
rect 26332 27072 26384 27124
rect 30472 27072 30524 27124
rect 32036 27072 32088 27124
rect 32312 27115 32364 27124
rect 32312 27081 32321 27115
rect 32321 27081 32355 27115
rect 32355 27081 32364 27115
rect 32312 27072 32364 27081
rect 48136 27115 48188 27124
rect 48136 27081 48145 27115
rect 48145 27081 48179 27115
rect 48179 27081 48188 27115
rect 48136 27072 48188 27081
rect 27160 26936 27212 26988
rect 27436 26979 27488 26988
rect 27436 26945 27445 26979
rect 27445 26945 27479 26979
rect 27479 26945 27488 26979
rect 27436 26936 27488 26945
rect 28448 26979 28500 26988
rect 28448 26945 28457 26979
rect 28457 26945 28491 26979
rect 28491 26945 28500 26979
rect 28448 26936 28500 26945
rect 27344 26911 27396 26920
rect 22468 26800 22520 26852
rect 24952 26843 25004 26852
rect 24952 26809 24961 26843
rect 24961 26809 24995 26843
rect 24995 26809 25004 26843
rect 24952 26800 25004 26809
rect 27344 26877 27353 26911
rect 27353 26877 27387 26911
rect 27387 26877 27396 26911
rect 27344 26868 27396 26877
rect 31208 27004 31260 27056
rect 29828 26936 29880 26988
rect 30288 26979 30340 26988
rect 30288 26945 30297 26979
rect 30297 26945 30331 26979
rect 30331 26945 30340 26979
rect 30288 26936 30340 26945
rect 30472 26979 30524 26988
rect 30472 26945 30481 26979
rect 30481 26945 30515 26979
rect 30515 26945 30524 26979
rect 30472 26936 30524 26945
rect 30656 26936 30708 26988
rect 31116 26979 31168 26988
rect 31116 26945 31125 26979
rect 31125 26945 31159 26979
rect 31159 26945 31168 26979
rect 31116 26936 31168 26945
rect 32772 27004 32824 27056
rect 34060 27004 34112 27056
rect 32036 26868 32088 26920
rect 33048 26936 33100 26988
rect 39580 26936 39632 26988
rect 32772 26868 32824 26920
rect 30104 26800 30156 26852
rect 24860 26732 24912 26784
rect 30380 26775 30432 26784
rect 30380 26741 30389 26775
rect 30389 26741 30423 26775
rect 30423 26741 30432 26775
rect 30380 26732 30432 26741
rect 36360 26732 36412 26784
rect 39580 26732 39632 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 19616 26571 19668 26580
rect 19616 26537 19625 26571
rect 19625 26537 19659 26571
rect 19659 26537 19668 26571
rect 19616 26528 19668 26537
rect 20168 26571 20220 26580
rect 20168 26537 20177 26571
rect 20177 26537 20211 26571
rect 20211 26537 20220 26571
rect 20168 26528 20220 26537
rect 21088 26528 21140 26580
rect 22192 26528 22244 26580
rect 23112 26528 23164 26580
rect 25044 26571 25096 26580
rect 25044 26537 25053 26571
rect 25053 26537 25087 26571
rect 25087 26537 25096 26571
rect 25044 26528 25096 26537
rect 26516 26571 26568 26580
rect 26516 26537 26525 26571
rect 26525 26537 26559 26571
rect 26559 26537 26568 26571
rect 26516 26528 26568 26537
rect 29828 26571 29880 26580
rect 29828 26537 29837 26571
rect 29837 26537 29871 26571
rect 29871 26537 29880 26571
rect 29828 26528 29880 26537
rect 30656 26528 30708 26580
rect 33048 26528 33100 26580
rect 24032 26460 24084 26512
rect 22284 26392 22336 26444
rect 36544 26460 36596 26512
rect 19616 26324 19668 26376
rect 20536 26324 20588 26376
rect 21824 26324 21876 26376
rect 22928 26324 22980 26376
rect 25136 26324 25188 26376
rect 25780 26324 25832 26376
rect 30288 26392 30340 26444
rect 1584 26256 1636 26308
rect 10784 26256 10836 26308
rect 22468 26256 22520 26308
rect 26240 26324 26292 26376
rect 29828 26324 29880 26376
rect 31576 26392 31628 26444
rect 33600 26392 33652 26444
rect 27436 26256 27488 26308
rect 28448 26256 28500 26308
rect 31116 26256 31168 26308
rect 33232 26324 33284 26376
rect 48136 26367 48188 26376
rect 48136 26333 48145 26367
rect 48145 26333 48179 26367
rect 48179 26333 48188 26367
rect 48136 26324 48188 26333
rect 30472 26231 30524 26240
rect 30472 26197 30481 26231
rect 30481 26197 30515 26231
rect 30515 26197 30524 26231
rect 30472 26188 30524 26197
rect 31024 26188 31076 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 21824 26027 21876 26036
rect 21824 25993 21833 26027
rect 21833 25993 21867 26027
rect 21867 25993 21876 26027
rect 21824 25984 21876 25993
rect 30196 25984 30248 26036
rect 31024 26027 31076 26036
rect 31024 25993 31033 26027
rect 31033 25993 31067 26027
rect 31067 25993 31076 26027
rect 31024 25984 31076 25993
rect 32772 26027 32824 26036
rect 32772 25993 32781 26027
rect 32781 25993 32815 26027
rect 32815 25993 32824 26027
rect 32772 25984 32824 25993
rect 1584 25959 1636 25968
rect 1584 25925 1593 25959
rect 1593 25925 1627 25959
rect 1627 25925 1636 25959
rect 1584 25916 1636 25925
rect 48136 25959 48188 25968
rect 48136 25925 48145 25959
rect 48145 25925 48179 25959
rect 48179 25925 48188 25959
rect 48136 25916 48188 25925
rect 24584 25891 24636 25900
rect 24584 25857 24593 25891
rect 24593 25857 24627 25891
rect 24627 25857 24636 25891
rect 24584 25848 24636 25857
rect 24768 25891 24820 25900
rect 24768 25857 24777 25891
rect 24777 25857 24811 25891
rect 24811 25857 24820 25891
rect 24768 25848 24820 25857
rect 28172 25848 28224 25900
rect 30380 25848 30432 25900
rect 31116 25848 31168 25900
rect 31576 25848 31628 25900
rect 26148 25780 26200 25832
rect 27712 25780 27764 25832
rect 29828 25823 29880 25832
rect 29828 25789 29837 25823
rect 29837 25789 29871 25823
rect 29871 25789 29880 25823
rect 29828 25780 29880 25789
rect 20536 25687 20588 25696
rect 20536 25653 20545 25687
rect 20545 25653 20579 25687
rect 20579 25653 20588 25687
rect 20536 25644 20588 25653
rect 22468 25687 22520 25696
rect 22468 25653 22477 25687
rect 22477 25653 22511 25687
rect 22511 25653 22520 25687
rect 22468 25644 22520 25653
rect 24860 25644 24912 25696
rect 26240 25687 26292 25696
rect 26240 25653 26249 25687
rect 26249 25653 26283 25687
rect 26283 25653 26292 25687
rect 26240 25644 26292 25653
rect 32036 25644 32088 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 27344 25440 27396 25492
rect 28172 25483 28224 25492
rect 28172 25449 28181 25483
rect 28181 25449 28215 25483
rect 28215 25449 28224 25483
rect 28172 25440 28224 25449
rect 28264 25440 28316 25492
rect 29276 25440 29328 25492
rect 31116 25440 31168 25492
rect 31576 25440 31628 25492
rect 25780 25415 25832 25424
rect 25780 25381 25789 25415
rect 25789 25381 25823 25415
rect 25823 25381 25832 25415
rect 25780 25372 25832 25381
rect 26148 25372 26200 25424
rect 29828 25372 29880 25424
rect 24952 25347 25004 25356
rect 24952 25313 24961 25347
rect 24961 25313 24995 25347
rect 24995 25313 25004 25347
rect 24952 25304 25004 25313
rect 24860 25279 24912 25288
rect 24860 25245 24869 25279
rect 24869 25245 24903 25279
rect 24903 25245 24912 25279
rect 24860 25236 24912 25245
rect 26700 25279 26752 25288
rect 26700 25245 26709 25279
rect 26709 25245 26743 25279
rect 26743 25245 26752 25279
rect 26700 25236 26752 25245
rect 28080 25279 28132 25288
rect 28080 25245 28089 25279
rect 28089 25245 28123 25279
rect 28123 25245 28132 25279
rect 28080 25236 28132 25245
rect 28264 25279 28316 25288
rect 28264 25245 28273 25279
rect 28273 25245 28307 25279
rect 28307 25245 28316 25279
rect 28264 25236 28316 25245
rect 27988 25168 28040 25220
rect 23756 25100 23808 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 26148 24896 26200 24948
rect 28080 24939 28132 24948
rect 28080 24905 28089 24939
rect 28089 24905 28123 24939
rect 28123 24905 28132 24939
rect 28080 24896 28132 24905
rect 23756 24803 23808 24812
rect 23756 24769 23765 24803
rect 23765 24769 23799 24803
rect 23799 24769 23808 24803
rect 23756 24760 23808 24769
rect 23940 24803 23992 24812
rect 23940 24769 23949 24803
rect 23949 24769 23983 24803
rect 23983 24769 23992 24803
rect 23940 24760 23992 24769
rect 24584 24803 24636 24812
rect 24584 24769 24593 24803
rect 24593 24769 24627 24803
rect 24627 24769 24636 24803
rect 24584 24760 24636 24769
rect 23204 24692 23256 24744
rect 24768 24692 24820 24744
rect 25044 24803 25096 24812
rect 25044 24769 25053 24803
rect 25053 24769 25087 24803
rect 25087 24769 25096 24803
rect 25044 24760 25096 24769
rect 26700 24760 26752 24812
rect 27160 24803 27212 24812
rect 27160 24769 27169 24803
rect 27169 24769 27203 24803
rect 27203 24769 27212 24803
rect 27160 24760 27212 24769
rect 27988 24803 28040 24812
rect 27988 24769 27997 24803
rect 27997 24769 28031 24803
rect 28031 24769 28040 24803
rect 27988 24760 28040 24769
rect 28264 24692 28316 24744
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 8944 24352 8996 24404
rect 24584 24352 24636 24404
rect 23940 24216 23992 24268
rect 23756 24148 23808 24200
rect 26608 24352 26660 24404
rect 27988 24352 28040 24404
rect 39764 24352 39816 24404
rect 48136 24080 48188 24132
rect 1492 24055 1544 24064
rect 1492 24021 1501 24055
rect 1501 24021 1535 24055
rect 1535 24021 1544 24055
rect 1492 24012 1544 24021
rect 23756 24055 23808 24064
rect 23756 24021 23765 24055
rect 23765 24021 23799 24055
rect 23799 24021 23808 24055
rect 23756 24012 23808 24021
rect 27160 24012 27212 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 48136 23851 48188 23860
rect 48136 23817 48145 23851
rect 48145 23817 48179 23851
rect 48179 23817 48188 23851
rect 48136 23808 48188 23817
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 37004 21972 37056 22024
rect 1584 21904 1636 21956
rect 15752 21836 15804 21888
rect 48044 21879 48096 21888
rect 48044 21845 48053 21879
rect 48053 21845 48087 21879
rect 48087 21845 48096 21879
rect 48044 21836 48096 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 1584 21675 1636 21684
rect 1584 21641 1593 21675
rect 1593 21641 1627 21675
rect 1627 21641 1636 21675
rect 1584 21632 1636 21641
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 39396 20000 39448 20052
rect 1860 19771 1912 19780
rect 1860 19737 1869 19771
rect 1869 19737 1903 19771
rect 1903 19737 1912 19771
rect 1860 19728 1912 19737
rect 14004 19660 14056 19712
rect 48044 19703 48096 19712
rect 48044 19669 48053 19703
rect 48053 19669 48087 19703
rect 48087 19669 48096 19703
rect 48044 19660 48096 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 1860 19456 1912 19508
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 1584 18232 1636 18284
rect 41236 18232 41288 18284
rect 47676 18232 47728 18284
rect 9864 18028 9916 18080
rect 48044 18071 48096 18080
rect 48044 18037 48053 18071
rect 48053 18037 48087 18071
rect 48087 18037 48096 18071
rect 48044 18028 48096 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 47676 17867 47728 17876
rect 47676 17833 47685 17867
rect 47685 17833 47719 17867
rect 47719 17833 47728 17867
rect 47676 17824 47728 17833
rect 1584 17799 1636 17808
rect 1584 17765 1593 17799
rect 1593 17765 1627 17799
rect 1627 17765 1636 17799
rect 1584 17756 1636 17765
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 42064 16192 42116 16244
rect 1584 16056 1636 16108
rect 48136 16099 48188 16108
rect 48136 16065 48145 16099
rect 48145 16065 48179 16099
rect 48179 16065 48188 16099
rect 48136 16056 48188 16065
rect 39580 15852 39632 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 1584 15691 1636 15700
rect 1584 15657 1593 15691
rect 1593 15657 1627 15691
rect 1627 15657 1636 15691
rect 1584 15648 1636 15657
rect 48136 15691 48188 15700
rect 48136 15657 48145 15691
rect 48145 15657 48179 15691
rect 48179 15657 48188 15691
rect 48136 15648 48188 15657
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 47860 13923 47912 13932
rect 47860 13889 47869 13923
rect 47869 13889 47903 13923
rect 47903 13889 47912 13923
rect 47860 13880 47912 13889
rect 35624 13812 35676 13864
rect 48044 13719 48096 13728
rect 48044 13685 48053 13719
rect 48053 13685 48087 13719
rect 48087 13685 48096 13719
rect 48044 13676 48096 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 1400 13515 1452 13524
rect 1400 13481 1409 13515
rect 1409 13481 1443 13515
rect 1443 13481 1452 13515
rect 1400 13472 1452 13481
rect 47860 13472 47912 13524
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 47768 11840 47820 11892
rect 48136 11747 48188 11756
rect 1492 11611 1544 11620
rect 1492 11577 1501 11611
rect 1501 11577 1535 11611
rect 1535 11577 1544 11611
rect 1492 11568 1544 11577
rect 48136 11713 48145 11747
rect 48145 11713 48179 11747
rect 48179 11713 48188 11747
rect 48136 11704 48188 11713
rect 27436 11568 27488 11620
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 48136 11339 48188 11348
rect 48136 11305 48145 11339
rect 48145 11305 48179 11339
rect 48179 11305 48188 11339
rect 48136 11296 48188 11305
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 31668 10004 31720 10056
rect 1584 9936 1636 9988
rect 31116 9868 31168 9920
rect 48044 9911 48096 9920
rect 48044 9877 48053 9911
rect 48053 9877 48087 9911
rect 48087 9877 48096 9911
rect 48044 9868 48096 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 1584 9639 1636 9648
rect 1584 9605 1593 9639
rect 1593 9605 1627 9639
rect 1627 9605 1636 9639
rect 1584 9596 1636 9605
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 47952 8075 48004 8084
rect 47952 8041 47961 8075
rect 47961 8041 47995 8075
rect 47995 8041 48004 8075
rect 47952 8032 48004 8041
rect 14924 7828 14976 7880
rect 48044 7803 48096 7812
rect 48044 7769 48053 7803
rect 48053 7769 48087 7803
rect 48087 7769 48096 7803
rect 48044 7760 48096 7769
rect 1492 7735 1544 7744
rect 1492 7701 1501 7735
rect 1501 7701 1535 7735
rect 1535 7701 1544 7735
rect 1492 7692 1544 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 1584 5584 1636 5636
rect 11520 5516 11572 5568
rect 22468 5516 22520 5568
rect 48044 5627 48096 5636
rect 48044 5593 48053 5627
rect 48053 5593 48087 5627
rect 48087 5593 48096 5627
rect 48044 5584 48096 5593
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 1584 5355 1636 5364
rect 1584 5321 1593 5355
rect 1593 5321 1627 5355
rect 1627 5321 1636 5355
rect 1584 5312 1636 5321
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 39488 4088 39540 4140
rect 47768 4088 47820 4140
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 47308 3587 47360 3596
rect 47308 3553 47317 3587
rect 47317 3553 47351 3587
rect 47351 3553 47360 3587
rect 47308 3544 47360 3553
rect 15476 3408 15528 3460
rect 48320 3408 48372 3460
rect 1492 3383 1544 3392
rect 1492 3349 1501 3383
rect 1501 3349 1535 3383
rect 1535 3349 1544 3383
rect 1492 3340 1544 3349
rect 48044 3383 48096 3392
rect 48044 3349 48053 3383
rect 48053 3349 48087 3383
rect 48087 3349 48096 3383
rect 48044 3340 48096 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 32588 3136 32640 3188
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 48320 3000 48372 3052
rect 49608 3000 49660 3052
rect 4620 2932 4672 2984
rect 28816 2932 28868 2984
rect 46572 2975 46624 2984
rect 46572 2941 46581 2975
rect 46581 2941 46615 2975
rect 46615 2941 46624 2975
rect 46572 2932 46624 2941
rect 10968 2864 11020 2916
rect 11980 2907 12032 2916
rect 11980 2873 11989 2907
rect 11989 2873 12023 2907
rect 12023 2873 12032 2907
rect 11980 2864 12032 2873
rect 36084 2864 36136 2916
rect 20 2796 72 2848
rect 2136 2839 2188 2848
rect 2136 2805 2145 2839
rect 2145 2805 2179 2839
rect 2179 2805 2188 2839
rect 2136 2796 2188 2805
rect 9036 2796 9088 2848
rect 16764 2796 16816 2848
rect 18696 2796 18748 2848
rect 19708 2796 19760 2848
rect 20720 2796 20772 2848
rect 24492 2796 24544 2848
rect 28356 2839 28408 2848
rect 28356 2805 28365 2839
rect 28365 2805 28399 2839
rect 28399 2805 28408 2839
rect 28356 2796 28408 2805
rect 40040 2796 40092 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 9772 2592 9824 2644
rect 20904 2635 20956 2644
rect 20904 2601 20913 2635
rect 20913 2601 20947 2635
rect 20947 2601 20956 2635
rect 20904 2592 20956 2601
rect 9496 2524 9548 2576
rect 14556 2524 14608 2576
rect 23204 2592 23256 2644
rect 26240 2592 26292 2644
rect 36360 2635 36412 2644
rect 22560 2524 22612 2576
rect 2136 2431 2188 2440
rect 2136 2397 2145 2431
rect 2145 2397 2179 2431
rect 2179 2397 2188 2431
rect 2136 2388 2188 2397
rect 4620 2388 4672 2440
rect 5172 2388 5224 2440
rect 1308 2320 1360 2372
rect 7104 2320 7156 2372
rect 9036 2320 9088 2372
rect 11980 2388 12032 2440
rect 14832 2388 14884 2440
rect 15200 2431 15252 2440
rect 15200 2397 15209 2431
rect 15209 2397 15243 2431
rect 15243 2397 15252 2431
rect 15200 2388 15252 2397
rect 19708 2431 19760 2440
rect 19708 2397 19717 2431
rect 19717 2397 19751 2431
rect 19751 2397 19760 2431
rect 19708 2388 19760 2397
rect 12900 2320 12952 2372
rect 16764 2320 16816 2372
rect 20536 2456 20588 2508
rect 25504 2524 25556 2576
rect 36360 2601 36369 2635
rect 36369 2601 36403 2635
rect 36403 2601 36412 2635
rect 36360 2592 36412 2601
rect 45284 2635 45336 2644
rect 45284 2601 45293 2635
rect 45293 2601 45327 2635
rect 45327 2601 45336 2635
rect 45284 2592 45336 2601
rect 44180 2567 44232 2576
rect 20720 2431 20772 2440
rect 20720 2397 20729 2431
rect 20729 2397 20763 2431
rect 20763 2397 20772 2431
rect 20720 2388 20772 2397
rect 22560 2388 22612 2440
rect 23756 2320 23808 2372
rect 24492 2320 24544 2372
rect 28448 2456 28500 2508
rect 30656 2499 30708 2508
rect 30656 2465 30665 2499
rect 30665 2465 30699 2499
rect 30699 2465 30708 2499
rect 30656 2456 30708 2465
rect 28356 2320 28408 2372
rect 30288 2388 30340 2440
rect 32588 2431 32640 2440
rect 32588 2397 32597 2431
rect 32597 2397 32631 2431
rect 32631 2397 32640 2431
rect 32588 2388 32640 2397
rect 44180 2533 44189 2567
rect 44189 2533 44223 2567
rect 44223 2533 44232 2567
rect 44180 2524 44232 2533
rect 40040 2431 40092 2440
rect 40040 2397 40049 2431
rect 40049 2397 40083 2431
rect 40083 2397 40092 2431
rect 40040 2388 40092 2397
rect 36084 2320 36136 2372
rect 45284 2388 45336 2440
rect 46572 2388 46624 2440
rect 47768 2431 47820 2440
rect 47768 2397 47777 2431
rect 47777 2397 47811 2431
rect 47811 2397 47820 2431
rect 47768 2388 47820 2397
rect 43812 2320 43864 2372
rect 2320 2295 2372 2304
rect 2320 2261 2329 2295
rect 2329 2261 2363 2295
rect 2363 2261 2372 2295
rect 2320 2252 2372 2261
rect 3240 2252 3292 2304
rect 10968 2252 11020 2304
rect 14832 2252 14884 2304
rect 17224 2295 17276 2304
rect 17224 2261 17233 2295
rect 17233 2261 17267 2295
rect 17267 2261 17276 2295
rect 17224 2252 17276 2261
rect 24952 2295 25004 2304
rect 24952 2261 24961 2295
rect 24961 2261 24995 2295
rect 24995 2261 25004 2295
rect 24952 2252 25004 2261
rect 26424 2295 26476 2304
rect 26424 2261 26433 2295
rect 26433 2261 26467 2295
rect 26467 2261 26476 2295
rect 26424 2252 26476 2261
rect 32220 2252 32272 2304
rect 34152 2295 34204 2304
rect 34152 2261 34161 2295
rect 34161 2261 34195 2295
rect 34195 2261 34204 2295
rect 34152 2252 34204 2261
rect 38016 2252 38068 2304
rect 40224 2295 40276 2304
rect 40224 2261 40233 2295
rect 40233 2261 40267 2295
rect 40267 2261 40276 2295
rect 40224 2252 40276 2261
rect 41880 2295 41932 2304
rect 41880 2261 41889 2295
rect 41889 2261 41923 2295
rect 41923 2261 41932 2295
rect 41880 2252 41932 2261
rect 42616 2295 42668 2304
rect 42616 2261 42625 2295
rect 42625 2261 42659 2295
rect 42659 2261 42668 2295
rect 42616 2252 42668 2261
rect 45744 2252 45796 2304
rect 46848 2252 46900 2304
rect 47676 2252 47728 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 2320 2048 2372 2100
rect 32036 2048 32088 2100
rect 17224 1980 17276 2032
rect 27160 1980 27212 2032
rect 24952 1912 25004 1964
rect 33968 1912 34020 1964
rect 13360 1844 13412 1896
rect 40224 1844 40276 1896
rect 20352 1776 20404 1828
rect 42616 1980 42668 2032
<< metal2 >>
rect 18 49200 74 50000
rect 1950 49200 2006 50000
rect 3882 49314 3938 50000
rect 3882 49286 4016 49314
rect 3882 49200 3938 49286
rect 32 46918 60 49200
rect 1964 46918 1992 49200
rect 2778 48376 2834 48385
rect 2778 48311 2834 48320
rect 2688 47048 2740 47054
rect 2688 46990 2740 46996
rect 20 46912 72 46918
rect 20 46854 72 46860
rect 1952 46912 2004 46918
rect 1952 46854 2004 46860
rect 2504 46912 2556 46918
rect 2504 46854 2556 46860
rect 2516 46714 2544 46854
rect 2700 46714 2728 46990
rect 2504 46708 2556 46714
rect 2504 46650 2556 46656
rect 2688 46708 2740 46714
rect 2688 46650 2740 46656
rect 1400 46572 1452 46578
rect 1400 46514 1452 46520
rect 1412 46345 1440 46514
rect 2688 46368 2740 46374
rect 1398 46336 1454 46345
rect 2688 46310 2740 46316
rect 1398 46271 1454 46280
rect 1412 46170 1440 46271
rect 1400 46164 1452 46170
rect 1400 46106 1452 46112
rect 1676 45960 1728 45966
rect 1676 45902 1728 45908
rect 1688 45626 1716 45902
rect 1952 45824 2004 45830
rect 1952 45766 2004 45772
rect 1964 45626 1992 45766
rect 1676 45620 1728 45626
rect 1676 45562 1728 45568
rect 1952 45620 2004 45626
rect 1952 45562 2004 45568
rect 1400 44396 1452 44402
rect 1400 44338 1452 44344
rect 1412 44305 1440 44338
rect 1398 44296 1454 44305
rect 1398 44231 1454 44240
rect 1412 43994 1440 44231
rect 1676 44192 1728 44198
rect 1676 44134 1728 44140
rect 1400 43988 1452 43994
rect 1400 43930 1452 43936
rect 1492 42560 1544 42566
rect 1492 42502 1544 42508
rect 1504 42265 1532 42502
rect 1490 42256 1546 42265
rect 1490 42191 1546 42200
rect 1584 40452 1636 40458
rect 1584 40394 1636 40400
rect 1596 40225 1624 40394
rect 1582 40216 1638 40225
rect 1582 40151 1584 40160
rect 1636 40151 1638 40160
rect 1584 40122 1636 40128
rect 1584 38276 1636 38282
rect 1584 38218 1636 38224
rect 1596 38185 1624 38218
rect 1582 38176 1638 38185
rect 1582 38111 1638 38120
rect 1596 38010 1624 38111
rect 1584 38004 1636 38010
rect 1584 37946 1636 37952
rect 1490 36136 1546 36145
rect 1490 36071 1546 36080
rect 1504 36038 1532 36071
rect 1492 36032 1544 36038
rect 1492 35974 1544 35980
rect 1584 34604 1636 34610
rect 1584 34546 1636 34552
rect 1596 34134 1624 34546
rect 1584 34128 1636 34134
rect 1582 34096 1584 34105
rect 1636 34096 1638 34105
rect 1582 34031 1638 34040
rect 1688 33561 1716 44134
rect 2044 40452 2096 40458
rect 2044 40394 2096 40400
rect 1952 35012 2004 35018
rect 1952 34954 2004 34960
rect 1964 34746 1992 34954
rect 1952 34740 2004 34746
rect 1952 34682 2004 34688
rect 2056 33658 2084 40394
rect 2700 39001 2728 46310
rect 2792 45966 2820 48311
rect 3988 47054 4016 49286
rect 5814 49200 5870 50000
rect 7746 49314 7802 50000
rect 9678 49314 9734 50000
rect 7746 49286 7880 49314
rect 7746 49200 7802 49286
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 5828 47258 5856 49200
rect 5816 47252 5868 47258
rect 5816 47194 5868 47200
rect 7852 47054 7880 49286
rect 9678 49286 9812 49314
rect 9678 49200 9734 49286
rect 9588 47184 9640 47190
rect 9588 47126 9640 47132
rect 9128 47116 9180 47122
rect 9128 47058 9180 47064
rect 3976 47048 4028 47054
rect 3976 46990 4028 46996
rect 6828 47048 6880 47054
rect 6828 46990 6880 46996
rect 7840 47048 7892 47054
rect 7840 46990 7892 46996
rect 2872 46980 2924 46986
rect 2872 46922 2924 46928
rect 2780 45960 2832 45966
rect 2780 45902 2832 45908
rect 2686 38992 2742 39001
rect 2686 38927 2742 38936
rect 2044 33652 2096 33658
rect 2044 33594 2096 33600
rect 1674 33552 1730 33561
rect 1674 33487 1730 33496
rect 1584 32428 1636 32434
rect 1584 32370 1636 32376
rect 1596 32065 1624 32370
rect 1952 32224 2004 32230
rect 1952 32166 2004 32172
rect 1582 32056 1638 32065
rect 1582 31991 1584 32000
rect 1636 31991 1638 32000
rect 1584 31962 1636 31968
rect 1964 31958 1992 32166
rect 1952 31952 2004 31958
rect 1952 31894 2004 31900
rect 1584 30252 1636 30258
rect 1584 30194 1636 30200
rect 1596 30025 1624 30194
rect 1582 30016 1638 30025
rect 1582 29951 1638 29960
rect 1596 29850 1624 29951
rect 1584 29844 1636 29850
rect 1584 29786 1636 29792
rect 2884 28121 2912 46922
rect 6840 46374 6868 46990
rect 8024 46912 8076 46918
rect 8024 46854 8076 46860
rect 6828 46368 6880 46374
rect 6828 46310 6880 46316
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 6840 44810 6868 46310
rect 6828 44804 6880 44810
rect 6828 44746 6880 44752
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 8036 34105 8064 46854
rect 9140 35494 9168 47058
rect 9600 46646 9628 47126
rect 9784 47122 9812 49286
rect 11610 49200 11666 50000
rect 13542 49200 13598 50000
rect 15474 49200 15530 50000
rect 17406 49200 17462 50000
rect 19338 49200 19394 50000
rect 21270 49200 21326 50000
rect 23202 49200 23258 50000
rect 25134 49314 25190 50000
rect 25134 49286 25544 49314
rect 25134 49200 25190 49286
rect 9772 47116 9824 47122
rect 9772 47058 9824 47064
rect 9588 46640 9640 46646
rect 9588 46582 9640 46588
rect 9312 46368 9364 46374
rect 9312 46310 9364 46316
rect 9324 46102 9352 46310
rect 9312 46096 9364 46102
rect 9312 46038 9364 46044
rect 9680 45554 9732 45558
rect 9784 45554 9812 47058
rect 11624 47054 11652 49200
rect 13556 47258 13584 49200
rect 14280 47456 14332 47462
rect 14280 47398 14332 47404
rect 13544 47252 13596 47258
rect 13544 47194 13596 47200
rect 12348 47116 12400 47122
rect 12348 47058 12400 47064
rect 12532 47116 12584 47122
rect 12532 47058 12584 47064
rect 14188 47116 14240 47122
rect 14188 47058 14240 47064
rect 11612 47048 11664 47054
rect 11612 46990 11664 46996
rect 9864 46980 9916 46986
rect 9864 46922 9916 46928
rect 10876 46980 10928 46986
rect 10876 46922 10928 46928
rect 9876 46442 9904 46922
rect 10416 46912 10468 46918
rect 10416 46854 10468 46860
rect 10428 46714 10456 46854
rect 10416 46708 10468 46714
rect 10416 46650 10468 46656
rect 10888 46510 10916 46922
rect 10876 46504 10928 46510
rect 10876 46446 10928 46452
rect 9864 46436 9916 46442
rect 9864 46378 9916 46384
rect 10784 46436 10836 46442
rect 10784 46378 10836 46384
rect 10232 45824 10284 45830
rect 10232 45766 10284 45772
rect 9680 45552 9812 45554
rect 9732 45526 9812 45552
rect 9680 45494 9732 45500
rect 10244 44878 10272 45766
rect 10416 45280 10468 45286
rect 10416 45222 10468 45228
rect 10232 44872 10284 44878
rect 10232 44814 10284 44820
rect 9864 44736 9916 44742
rect 9864 44678 9916 44684
rect 9876 44402 9904 44678
rect 10428 44538 10456 45222
rect 10416 44532 10468 44538
rect 10416 44474 10468 44480
rect 9864 44396 9916 44402
rect 9864 44338 9916 44344
rect 9876 44198 9904 44338
rect 9864 44192 9916 44198
rect 9864 44134 9916 44140
rect 9876 43654 9904 44134
rect 9864 43648 9916 43654
rect 9864 43590 9916 43596
rect 9588 42764 9640 42770
rect 9588 42706 9640 42712
rect 9600 42566 9628 42706
rect 9588 42560 9640 42566
rect 9588 42502 9640 42508
rect 9600 41478 9628 42502
rect 9588 41472 9640 41478
rect 9588 41414 9640 41420
rect 9128 35488 9180 35494
rect 9128 35430 9180 35436
rect 9140 34746 9168 35430
rect 9128 34740 9180 34746
rect 9128 34682 9180 34688
rect 8022 34096 8078 34105
rect 8022 34031 8078 34040
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 8944 32224 8996 32230
rect 8944 32166 8996 32172
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 2870 28112 2926 28121
rect 2870 28047 2926 28056
rect 1490 27976 1546 27985
rect 1490 27911 1492 27920
rect 1544 27911 1546 27920
rect 1492 27882 1544 27888
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 1584 26308 1636 26314
rect 1584 26250 1636 26256
rect 1596 25974 1624 26250
rect 1584 25968 1636 25974
rect 1582 25936 1584 25945
rect 1636 25936 1638 25945
rect 1582 25871 1638 25880
rect 1596 25845 1624 25871
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 8956 24410 8984 32166
rect 8944 24404 8996 24410
rect 8944 24346 8996 24352
rect 1492 24064 1544 24070
rect 1492 24006 1544 24012
rect 1504 23905 1532 24006
rect 1490 23896 1546 23905
rect 1490 23831 1546 23840
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 1584 21956 1636 21962
rect 1584 21898 1636 21904
rect 1596 21865 1624 21898
rect 1582 21856 1638 21865
rect 1582 21791 1638 21800
rect 1596 21690 1624 21791
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 1858 19816 1914 19825
rect 1858 19751 1860 19760
rect 1912 19751 1914 19760
rect 1860 19722 1912 19728
rect 1872 19514 1900 19722
rect 1860 19508 1912 19514
rect 1860 19450 1912 19456
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 1584 18284 1636 18290
rect 1584 18226 1636 18232
rect 1596 17814 1624 18226
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 1584 17808 1636 17814
rect 1582 17776 1584 17785
rect 1636 17776 1638 17785
rect 1582 17711 1638 17720
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 1584 16108 1636 16114
rect 1584 16050 1636 16056
rect 1596 15745 1624 16050
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 1582 15736 1638 15745
rect 4214 15739 4522 15748
rect 1582 15671 1584 15680
rect 1636 15671 1638 15680
rect 1584 15642 1636 15648
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 13705 1440 13874
rect 1398 13696 1454 13705
rect 1398 13631 1454 13640
rect 1412 13530 1440 13631
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 1400 13524 1452 13530
rect 1400 13466 1452 13472
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 1490 11656 1546 11665
rect 1490 11591 1492 11600
rect 1544 11591 1546 11600
rect 1492 11562 1544 11568
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 1584 9988 1636 9994
rect 1584 9930 1636 9936
rect 1596 9654 1624 9930
rect 1584 9648 1636 9654
rect 1582 9616 1584 9625
rect 1636 9616 1638 9625
rect 1582 9551 1638 9560
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 1492 7744 1544 7750
rect 1492 7686 1544 7692
rect 1504 7585 1532 7686
rect 1490 7576 1546 7585
rect 1490 7511 1546 7520
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 9600 6914 9628 41414
rect 9772 34400 9824 34406
rect 9772 34342 9824 34348
rect 9784 33862 9812 34342
rect 9772 33856 9824 33862
rect 9772 33798 9824 33804
rect 9508 6886 9628 6914
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 1584 5636 1636 5642
rect 1584 5578 1636 5584
rect 1596 5545 1624 5578
rect 1582 5536 1638 5545
rect 1582 5471 1638 5480
rect 1596 5370 1624 5471
rect 1584 5364 1636 5370
rect 1584 5306 1636 5312
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 1490 3496 1546 3505
rect 1490 3431 1546 3440
rect 1504 3398 1532 3431
rect 1492 3392 1544 3398
rect 1492 3334 1544 3340
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 20 2848 72 2854
rect 20 2790 72 2796
rect 32 800 60 2790
rect 1308 2372 1360 2378
rect 1308 2314 1360 2320
rect 1320 800 1348 2314
rect 1412 1465 1440 2994
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 2136 2848 2188 2854
rect 2136 2790 2188 2796
rect 2148 2446 2176 2790
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2446 4660 2926
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 2136 2440 2188 2446
rect 2136 2382 2188 2388
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 2320 2304 2372 2310
rect 2320 2246 2372 2252
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 2332 2106 2360 2246
rect 2320 2100 2372 2106
rect 2320 2042 2372 2048
rect 1398 1456 1454 1465
rect 1398 1391 1454 1400
rect 3252 800 3280 2246
rect 5184 800 5212 2382
rect 9048 2378 9076 2790
rect 9508 2582 9536 6886
rect 9784 2650 9812 33798
rect 9876 18086 9904 43590
rect 10796 43450 10824 46378
rect 10888 44810 10916 46446
rect 11624 46170 11652 46990
rect 11612 46164 11664 46170
rect 11612 46106 11664 46112
rect 11704 45824 11756 45830
rect 11704 45766 11756 45772
rect 11888 45824 11940 45830
rect 11888 45766 11940 45772
rect 11152 45620 11204 45626
rect 11152 45562 11204 45568
rect 10876 44804 10928 44810
rect 10876 44746 10928 44752
rect 10888 43790 10916 44746
rect 10968 44192 11020 44198
rect 10968 44134 11020 44140
rect 10876 43784 10928 43790
rect 10876 43726 10928 43732
rect 10980 43722 11008 44134
rect 10968 43716 11020 43722
rect 10968 43658 11020 43664
rect 10784 43444 10836 43450
rect 10784 43386 10836 43392
rect 10796 42922 10824 43386
rect 10980 43382 11008 43658
rect 10968 43376 11020 43382
rect 10968 43318 11020 43324
rect 10796 42894 10916 42922
rect 10980 42906 11008 43318
rect 10888 42786 10916 42894
rect 10968 42900 11020 42906
rect 10968 42842 11020 42848
rect 10888 42758 11100 42786
rect 10784 42696 10836 42702
rect 10784 42638 10836 42644
rect 10796 42566 10824 42638
rect 10784 42560 10836 42566
rect 10784 42502 10836 42508
rect 10796 42022 10824 42502
rect 11072 42362 11100 42758
rect 11060 42356 11112 42362
rect 11060 42298 11112 42304
rect 10784 42016 10836 42022
rect 10784 41958 10836 41964
rect 10232 38752 10284 38758
rect 10232 38694 10284 38700
rect 10244 35834 10272 38694
rect 10324 37664 10376 37670
rect 10324 37606 10376 37612
rect 10336 37330 10364 37606
rect 10324 37324 10376 37330
rect 10324 37266 10376 37272
rect 10232 35828 10284 35834
rect 10232 35770 10284 35776
rect 10244 34746 10272 35770
rect 10232 34740 10284 34746
rect 10232 34682 10284 34688
rect 10244 34474 10272 34682
rect 10336 34542 10364 37266
rect 10324 34536 10376 34542
rect 10324 34478 10376 34484
rect 10232 34468 10284 34474
rect 10232 34410 10284 34416
rect 10244 34202 10272 34410
rect 10232 34196 10284 34202
rect 10232 34138 10284 34144
rect 10692 32564 10744 32570
rect 10692 32506 10744 32512
rect 10704 32026 10732 32506
rect 10692 32020 10744 32026
rect 10692 31962 10744 31968
rect 10796 26314 10824 41958
rect 11060 41540 11112 41546
rect 11060 41482 11112 41488
rect 11072 41138 11100 41482
rect 11060 41132 11112 41138
rect 11060 41074 11112 41080
rect 11072 40934 11100 41074
rect 11060 40928 11112 40934
rect 11060 40870 11112 40876
rect 10876 39364 10928 39370
rect 10876 39306 10928 39312
rect 10888 38758 10916 39306
rect 10876 38752 10928 38758
rect 10876 38694 10928 38700
rect 10968 37392 11020 37398
rect 10968 37334 11020 37340
rect 10980 36922 11008 37334
rect 10968 36916 11020 36922
rect 10888 36876 10968 36904
rect 10888 35290 10916 36876
rect 10968 36858 11020 36864
rect 11072 36802 11100 40870
rect 11164 39642 11192 45562
rect 11244 44736 11296 44742
rect 11244 44678 11296 44684
rect 11256 42702 11284 44678
rect 11716 43994 11744 45766
rect 11900 45558 11928 45766
rect 11888 45552 11940 45558
rect 11886 45520 11888 45529
rect 11940 45520 11942 45529
rect 11886 45455 11942 45464
rect 11900 45429 11928 45455
rect 12164 45280 12216 45286
rect 12164 45222 12216 45228
rect 12176 44334 12204 45222
rect 12164 44328 12216 44334
rect 12164 44270 12216 44276
rect 11704 43988 11756 43994
rect 11704 43930 11756 43936
rect 11796 43648 11848 43654
rect 11796 43590 11848 43596
rect 11244 42696 11296 42702
rect 11244 42638 11296 42644
rect 11808 42566 11836 43590
rect 11796 42560 11848 42566
rect 11796 42502 11848 42508
rect 11808 40118 11836 42502
rect 12072 42356 12124 42362
rect 12072 42298 12124 42304
rect 12084 40662 12112 42298
rect 12176 41546 12204 44270
rect 12256 42696 12308 42702
rect 12256 42638 12308 42644
rect 12268 42226 12296 42638
rect 12256 42220 12308 42226
rect 12256 42162 12308 42168
rect 12164 41540 12216 41546
rect 12164 41482 12216 41488
rect 12072 40656 12124 40662
rect 12072 40598 12124 40604
rect 11796 40112 11848 40118
rect 11796 40054 11848 40060
rect 12084 40050 12112 40598
rect 12072 40044 12124 40050
rect 12072 39986 12124 39992
rect 11152 39636 11204 39642
rect 11152 39578 11204 39584
rect 11164 38962 11192 39578
rect 12256 39296 12308 39302
rect 12256 39238 12308 39244
rect 11152 38956 11204 38962
rect 11152 38898 11204 38904
rect 11164 38554 11192 38898
rect 12268 38758 12296 39238
rect 12256 38752 12308 38758
rect 12256 38694 12308 38700
rect 11152 38548 11204 38554
rect 11152 38490 11204 38496
rect 10980 36774 11100 36802
rect 10876 35284 10928 35290
rect 10876 35226 10928 35232
rect 10876 33992 10928 33998
rect 10876 33934 10928 33940
rect 10888 33658 10916 33934
rect 10876 33652 10928 33658
rect 10876 33594 10928 33600
rect 10784 26308 10836 26314
rect 10784 26250 10836 26256
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 10980 2922 11008 36774
rect 11164 33590 11192 38490
rect 12268 38350 12296 38694
rect 12256 38344 12308 38350
rect 12256 38286 12308 38292
rect 11796 37460 11848 37466
rect 11796 37402 11848 37408
rect 11520 35080 11572 35086
rect 11520 35022 11572 35028
rect 11532 34406 11560 35022
rect 11520 34400 11572 34406
rect 11520 34342 11572 34348
rect 11532 34066 11560 34342
rect 11520 34060 11572 34066
rect 11520 34002 11572 34008
rect 11612 33992 11664 33998
rect 11612 33934 11664 33940
rect 11152 33584 11204 33590
rect 11152 33526 11204 33532
rect 11520 33516 11572 33522
rect 11520 33458 11572 33464
rect 11532 32910 11560 33458
rect 11624 33114 11652 33934
rect 11704 33584 11756 33590
rect 11704 33526 11756 33532
rect 11612 33108 11664 33114
rect 11612 33050 11664 33056
rect 11716 32910 11744 33526
rect 11520 32904 11572 32910
rect 11520 32846 11572 32852
rect 11704 32904 11756 32910
rect 11704 32846 11756 32852
rect 11532 5574 11560 32846
rect 11808 32026 11836 37402
rect 11888 36848 11940 36854
rect 11888 36790 11940 36796
rect 11900 36378 11928 36790
rect 11888 36372 11940 36378
rect 11888 36314 11940 36320
rect 11888 36100 11940 36106
rect 11888 36042 11940 36048
rect 11900 35494 11928 36042
rect 11888 35488 11940 35494
rect 11888 35430 11940 35436
rect 11900 33946 11928 35430
rect 11980 35080 12032 35086
rect 11980 35022 12032 35028
rect 11992 34746 12020 35022
rect 11980 34740 12032 34746
rect 11980 34682 12032 34688
rect 12072 34740 12124 34746
rect 12072 34682 12124 34688
rect 11992 34066 12020 34682
rect 11980 34060 12032 34066
rect 11980 34002 12032 34008
rect 12084 33998 12112 34682
rect 12072 33992 12124 33998
rect 11900 33918 12020 33946
rect 12072 33934 12124 33940
rect 11992 32978 12020 33918
rect 11980 32972 12032 32978
rect 11980 32914 12032 32920
rect 11992 32230 12020 32914
rect 11980 32224 12032 32230
rect 11980 32166 12032 32172
rect 11796 32020 11848 32026
rect 11796 31962 11848 31968
rect 11808 31793 11836 31962
rect 12360 31822 12388 47058
rect 12440 46368 12492 46374
rect 12440 46310 12492 46316
rect 12452 44810 12480 46310
rect 12544 45558 12572 47058
rect 14096 46912 14148 46918
rect 14096 46854 14148 46860
rect 12716 46640 12768 46646
rect 12714 46608 12716 46617
rect 12992 46640 13044 46646
rect 12768 46608 12770 46617
rect 13044 46600 13124 46628
rect 12992 46582 13044 46588
rect 12714 46543 12770 46552
rect 13096 46560 13124 46600
rect 13176 46572 13228 46578
rect 12728 46170 12756 46543
rect 13096 46532 13176 46560
rect 13176 46514 13228 46520
rect 13728 46572 13780 46578
rect 13728 46514 13780 46520
rect 13820 46572 13872 46578
rect 13820 46514 13872 46520
rect 12992 46504 13044 46510
rect 12992 46446 13044 46452
rect 12716 46164 12768 46170
rect 12716 46106 12768 46112
rect 12532 45552 12584 45558
rect 12532 45494 12584 45500
rect 12808 45484 12860 45490
rect 12808 45426 12860 45432
rect 12624 45280 12676 45286
rect 12624 45222 12676 45228
rect 12440 44804 12492 44810
rect 12440 44746 12492 44752
rect 12636 44538 12664 45222
rect 12820 44878 12848 45426
rect 13004 45354 13032 46446
rect 13452 46368 13504 46374
rect 13452 46310 13504 46316
rect 13464 46170 13492 46310
rect 13452 46164 13504 46170
rect 13452 46106 13504 46112
rect 13268 45484 13320 45490
rect 13268 45426 13320 45432
rect 12992 45348 13044 45354
rect 12992 45290 13044 45296
rect 13280 45082 13308 45426
rect 13268 45076 13320 45082
rect 13268 45018 13320 45024
rect 12808 44872 12860 44878
rect 12808 44814 12860 44820
rect 13268 44872 13320 44878
rect 13268 44814 13320 44820
rect 13360 44872 13412 44878
rect 13360 44814 13412 44820
rect 12820 44538 12848 44814
rect 13280 44538 13308 44814
rect 12624 44532 12676 44538
rect 12624 44474 12676 44480
rect 12808 44532 12860 44538
rect 12808 44474 12860 44480
rect 13268 44532 13320 44538
rect 13268 44474 13320 44480
rect 13268 44396 13320 44402
rect 13372 44384 13400 44814
rect 13320 44356 13400 44384
rect 13268 44338 13320 44344
rect 13464 44334 13492 46106
rect 13740 46034 13768 46514
rect 13728 46028 13780 46034
rect 13728 45970 13780 45976
rect 13832 44849 13860 46514
rect 14108 46442 14136 46854
rect 14096 46436 14148 46442
rect 14096 46378 14148 46384
rect 14108 45966 14136 46378
rect 14200 46170 14228 47058
rect 14292 47054 14320 47398
rect 15488 47258 15516 49200
rect 17224 47524 17276 47530
rect 17224 47466 17276 47472
rect 15476 47252 15528 47258
rect 15476 47194 15528 47200
rect 15752 47252 15804 47258
rect 15752 47194 15804 47200
rect 14740 47116 14792 47122
rect 14740 47058 14792 47064
rect 14280 47048 14332 47054
rect 14280 46990 14332 46996
rect 14292 46578 14320 46990
rect 14752 46578 14780 47058
rect 15764 47054 15792 47194
rect 17236 47190 17264 47466
rect 17224 47184 17276 47190
rect 17224 47126 17276 47132
rect 16856 47116 16908 47122
rect 16856 47058 16908 47064
rect 15752 47048 15804 47054
rect 15752 46990 15804 46996
rect 15292 46980 15344 46986
rect 15292 46922 15344 46928
rect 14280 46572 14332 46578
rect 14280 46514 14332 46520
rect 14740 46572 14792 46578
rect 14740 46514 14792 46520
rect 14188 46164 14240 46170
rect 14188 46106 14240 46112
rect 14096 45960 14148 45966
rect 14096 45902 14148 45908
rect 13912 45892 13964 45898
rect 13912 45834 13964 45840
rect 13924 45626 13952 45834
rect 13912 45620 13964 45626
rect 13912 45562 13964 45568
rect 13924 45490 13952 45562
rect 13912 45484 13964 45490
rect 13912 45426 13964 45432
rect 13818 44840 13874 44849
rect 13818 44775 13820 44784
rect 13872 44775 13874 44784
rect 13820 44746 13872 44752
rect 13832 44715 13860 44746
rect 13452 44328 13504 44334
rect 13452 44270 13504 44276
rect 12440 44260 12492 44266
rect 12440 44202 12492 44208
rect 12452 42362 12480 44202
rect 12990 43888 13046 43897
rect 12990 43823 13046 43832
rect 13084 43852 13136 43858
rect 12808 43784 12860 43790
rect 12808 43726 12860 43732
rect 12900 43784 12952 43790
rect 12900 43726 12952 43732
rect 12624 43172 12676 43178
rect 12624 43114 12676 43120
rect 12636 42838 12664 43114
rect 12624 42832 12676 42838
rect 12624 42774 12676 42780
rect 12440 42356 12492 42362
rect 12440 42298 12492 42304
rect 12452 40050 12480 42298
rect 12716 40928 12768 40934
rect 12716 40870 12768 40876
rect 12728 40730 12756 40870
rect 12716 40724 12768 40730
rect 12716 40666 12768 40672
rect 12728 40594 12756 40666
rect 12716 40588 12768 40594
rect 12716 40530 12768 40536
rect 12716 40112 12768 40118
rect 12716 40054 12768 40060
rect 12440 40044 12492 40050
rect 12440 39986 12492 39992
rect 12532 38344 12584 38350
rect 12532 38286 12584 38292
rect 12440 38208 12492 38214
rect 12440 38150 12492 38156
rect 12452 38010 12480 38150
rect 12440 38004 12492 38010
rect 12440 37946 12492 37952
rect 12440 37392 12492 37398
rect 12440 37334 12492 37340
rect 12452 37262 12480 37334
rect 12440 37256 12492 37262
rect 12440 37198 12492 37204
rect 12544 37126 12572 38286
rect 12532 37120 12584 37126
rect 12532 37062 12584 37068
rect 12440 36916 12492 36922
rect 12440 36858 12492 36864
rect 12452 36825 12480 36858
rect 12438 36816 12494 36825
rect 12438 36751 12494 36760
rect 12544 36650 12572 37062
rect 12532 36644 12584 36650
rect 12532 36586 12584 36592
rect 12440 35080 12492 35086
rect 12440 35022 12492 35028
rect 12452 34610 12480 35022
rect 12440 34604 12492 34610
rect 12440 34546 12492 34552
rect 12452 33114 12480 34546
rect 12440 33108 12492 33114
rect 12440 33050 12492 33056
rect 12544 31822 12572 36586
rect 12728 35834 12756 40054
rect 12820 39642 12848 43726
rect 12912 43450 12940 43726
rect 12900 43444 12952 43450
rect 12900 43386 12952 43392
rect 13004 43314 13032 43823
rect 13084 43794 13136 43800
rect 13096 43450 13124 43794
rect 13924 43450 13952 45426
rect 14004 44940 14056 44946
rect 14004 44882 14056 44888
rect 14016 44402 14044 44882
rect 14004 44396 14056 44402
rect 14004 44338 14056 44344
rect 14200 44282 14228 46106
rect 14280 45960 14332 45966
rect 14280 45902 14332 45908
rect 14292 45082 14320 45902
rect 14464 45892 14516 45898
rect 14464 45834 14516 45840
rect 14476 45558 14504 45834
rect 14464 45552 14516 45558
rect 14464 45494 14516 45500
rect 14464 45348 14516 45354
rect 14464 45290 14516 45296
rect 14280 45076 14332 45082
rect 14280 45018 14332 45024
rect 14476 44441 14504 45290
rect 14752 44878 14780 46514
rect 15304 46510 15332 46922
rect 15764 46646 15792 46990
rect 16488 46912 16540 46918
rect 16488 46854 16540 46860
rect 15752 46640 15804 46646
rect 15752 46582 15804 46588
rect 15292 46504 15344 46510
rect 15292 46446 15344 46452
rect 16500 45966 16528 46854
rect 16672 46572 16724 46578
rect 16672 46514 16724 46520
rect 16488 45960 16540 45966
rect 16488 45902 16540 45908
rect 16684 45898 16712 46514
rect 16764 46504 16816 46510
rect 16764 46446 16816 46452
rect 16776 45966 16804 46446
rect 16764 45960 16816 45966
rect 16764 45902 16816 45908
rect 16672 45892 16724 45898
rect 16672 45834 16724 45840
rect 16028 45824 16080 45830
rect 16028 45766 16080 45772
rect 16040 45286 16068 45766
rect 16776 45626 16804 45902
rect 16764 45620 16816 45626
rect 16764 45562 16816 45568
rect 16488 45484 16540 45490
rect 16488 45426 16540 45432
rect 16028 45280 16080 45286
rect 16028 45222 16080 45228
rect 14740 44872 14792 44878
rect 14646 44840 14702 44849
rect 14740 44814 14792 44820
rect 15108 44872 15160 44878
rect 15108 44814 15160 44820
rect 15476 44872 15528 44878
rect 15476 44814 15528 44820
rect 14646 44775 14648 44784
rect 14700 44775 14702 44784
rect 14648 44746 14700 44752
rect 14462 44432 14518 44441
rect 15120 44402 15148 44814
rect 15488 44402 15516 44814
rect 16040 44742 16068 45222
rect 16500 44878 16528 45426
rect 16580 45348 16632 45354
rect 16580 45290 16632 45296
rect 16592 44946 16620 45290
rect 16580 44940 16632 44946
rect 16580 44882 16632 44888
rect 16488 44872 16540 44878
rect 16488 44814 16540 44820
rect 16028 44736 16080 44742
rect 16028 44678 16080 44684
rect 16040 44538 16068 44678
rect 16028 44532 16080 44538
rect 16028 44474 16080 44480
rect 14462 44367 14518 44376
rect 15108 44396 15160 44402
rect 14200 44254 14320 44282
rect 14096 44192 14148 44198
rect 14096 44134 14148 44140
rect 14108 43994 14136 44134
rect 14096 43988 14148 43994
rect 14096 43930 14148 43936
rect 13084 43444 13136 43450
rect 13084 43386 13136 43392
rect 13912 43444 13964 43450
rect 13912 43386 13964 43392
rect 12992 43308 13044 43314
rect 12992 43250 13044 43256
rect 13096 42906 13124 43386
rect 13452 43240 13504 43246
rect 13452 43182 13504 43188
rect 13360 43172 13412 43178
rect 13360 43114 13412 43120
rect 13084 42900 13136 42906
rect 13084 42842 13136 42848
rect 12900 42764 12952 42770
rect 12900 42706 12952 42712
rect 12912 42566 12940 42706
rect 12992 42696 13044 42702
rect 12992 42638 13044 42644
rect 12900 42560 12952 42566
rect 12900 42502 12952 42508
rect 12912 40730 12940 42502
rect 13004 42226 13032 42638
rect 12992 42220 13044 42226
rect 12992 42162 13044 42168
rect 12900 40724 12952 40730
rect 12900 40666 12952 40672
rect 12808 39636 12860 39642
rect 12808 39578 12860 39584
rect 12900 39092 12952 39098
rect 12900 39034 12952 39040
rect 12912 38894 12940 39034
rect 12900 38888 12952 38894
rect 12900 38830 12952 38836
rect 12912 37738 12940 38830
rect 13176 38208 13228 38214
rect 13176 38150 13228 38156
rect 12900 37732 12952 37738
rect 12900 37674 12952 37680
rect 13188 37670 13216 38150
rect 13268 37936 13320 37942
rect 13268 37878 13320 37884
rect 13176 37664 13228 37670
rect 13176 37606 13228 37612
rect 13188 37194 13216 37606
rect 13176 37188 13228 37194
rect 13176 37130 13228 37136
rect 13188 36854 13216 37130
rect 13176 36848 13228 36854
rect 13176 36790 13228 36796
rect 12992 36168 13044 36174
rect 12992 36110 13044 36116
rect 12716 35828 12768 35834
rect 12716 35770 12768 35776
rect 13004 35766 13032 36110
rect 13280 35834 13308 37878
rect 13268 35828 13320 35834
rect 13268 35770 13320 35776
rect 12992 35760 13044 35766
rect 12992 35702 13044 35708
rect 12624 35148 12676 35154
rect 12624 35090 12676 35096
rect 12636 34678 12664 35090
rect 12808 35080 12860 35086
rect 12808 35022 12860 35028
rect 12716 34944 12768 34950
rect 12716 34886 12768 34892
rect 12624 34672 12676 34678
rect 12624 34614 12676 34620
rect 12728 34610 12756 34886
rect 12820 34746 12848 35022
rect 13268 35012 13320 35018
rect 13268 34954 13320 34960
rect 13280 34746 13308 34954
rect 12808 34740 12860 34746
rect 12808 34682 12860 34688
rect 13268 34740 13320 34746
rect 13268 34682 13320 34688
rect 12716 34604 12768 34610
rect 12716 34546 12768 34552
rect 12624 33856 12676 33862
rect 12624 33798 12676 33804
rect 12636 32434 12664 33798
rect 12728 33590 12756 34546
rect 13268 34060 13320 34066
rect 13268 34002 13320 34008
rect 12900 33992 12952 33998
rect 12900 33934 12952 33940
rect 12912 33590 12940 33934
rect 13280 33658 13308 34002
rect 13268 33652 13320 33658
rect 13268 33594 13320 33600
rect 12716 33584 12768 33590
rect 12716 33526 12768 33532
rect 12900 33584 12952 33590
rect 12900 33526 12952 33532
rect 12808 33516 12860 33522
rect 12808 33458 12860 33464
rect 12716 33312 12768 33318
rect 12716 33254 12768 33260
rect 12728 32434 12756 33254
rect 12820 32910 12848 33458
rect 12808 32904 12860 32910
rect 12912 32892 12940 33526
rect 12992 32904 13044 32910
rect 12912 32864 12992 32892
rect 12808 32846 12860 32852
rect 12992 32846 13044 32852
rect 12624 32428 12676 32434
rect 12624 32370 12676 32376
rect 12716 32428 12768 32434
rect 12716 32370 12768 32376
rect 12820 32298 12848 32846
rect 13176 32768 13228 32774
rect 13176 32710 13228 32716
rect 13188 32434 13216 32710
rect 13176 32428 13228 32434
rect 13176 32370 13228 32376
rect 12808 32292 12860 32298
rect 12808 32234 12860 32240
rect 12820 32026 12848 32234
rect 12808 32020 12860 32026
rect 12808 31962 12860 31968
rect 12348 31816 12400 31822
rect 11794 31784 11850 31793
rect 12348 31758 12400 31764
rect 12532 31816 12584 31822
rect 12532 31758 12584 31764
rect 11794 31719 11850 31728
rect 12360 31414 12388 31758
rect 12348 31408 12400 31414
rect 12348 31350 12400 31356
rect 12360 30734 12388 31350
rect 12544 31346 12572 31758
rect 12532 31340 12584 31346
rect 12532 31282 12584 31288
rect 12544 30734 12572 31282
rect 12992 31136 13044 31142
rect 12992 31078 13044 31084
rect 13004 30734 13032 31078
rect 12348 30728 12400 30734
rect 12348 30670 12400 30676
rect 12532 30728 12584 30734
rect 12532 30670 12584 30676
rect 12992 30728 13044 30734
rect 12992 30670 13044 30676
rect 12360 30394 12388 30670
rect 12544 30394 12572 30670
rect 12348 30388 12400 30394
rect 12348 30330 12400 30336
rect 12532 30388 12584 30394
rect 12532 30330 12584 30336
rect 13188 30258 13216 32370
rect 13268 32360 13320 32366
rect 13268 32302 13320 32308
rect 13280 30734 13308 32302
rect 13268 30728 13320 30734
rect 13268 30670 13320 30676
rect 13176 30252 13228 30258
rect 13176 30194 13228 30200
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11978 2952 12034 2961
rect 10968 2916 11020 2922
rect 11978 2887 11980 2896
rect 10968 2858 11020 2864
rect 12032 2887 12034 2896
rect 11980 2858 12032 2864
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 9496 2576 9548 2582
rect 9496 2518 9548 2524
rect 11992 2446 12020 2858
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 7104 2372 7156 2378
rect 7104 2314 7156 2320
rect 9036 2372 9088 2378
rect 9036 2314 9088 2320
rect 12900 2372 12952 2378
rect 12900 2314 12952 2320
rect 7116 800 7144 2314
rect 9048 800 9076 2314
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 10980 800 11008 2246
rect 12912 800 12940 2314
rect 13372 1902 13400 43114
rect 13464 42362 13492 43182
rect 13544 42764 13596 42770
rect 13544 42706 13596 42712
rect 13452 42356 13504 42362
rect 13452 42298 13504 42304
rect 13556 41818 13584 42706
rect 13820 42560 13872 42566
rect 13820 42502 13872 42508
rect 13544 41812 13596 41818
rect 13544 41754 13596 41760
rect 13544 41472 13596 41478
rect 13544 41414 13596 41420
rect 13556 41274 13584 41414
rect 13832 41274 13860 42502
rect 14108 42362 14136 43930
rect 14188 43104 14240 43110
rect 14188 43046 14240 43052
rect 14096 42356 14148 42362
rect 13924 42316 14096 42344
rect 13544 41268 13596 41274
rect 13544 41210 13596 41216
rect 13820 41268 13872 41274
rect 13820 41210 13872 41216
rect 13556 40934 13584 41210
rect 13544 40928 13596 40934
rect 13544 40870 13596 40876
rect 13832 40730 13860 41210
rect 13820 40724 13872 40730
rect 13820 40666 13872 40672
rect 13924 40186 13952 42316
rect 14096 42298 14148 42304
rect 14200 41818 14228 43046
rect 14188 41812 14240 41818
rect 14016 41772 14188 41800
rect 14016 41313 14044 41772
rect 14188 41754 14240 41760
rect 14292 41414 14320 44254
rect 14476 43994 14504 44367
rect 15292 44396 15344 44402
rect 15108 44338 15160 44344
rect 15212 44356 15292 44384
rect 15016 44328 15068 44334
rect 15016 44270 15068 44276
rect 14464 43988 14516 43994
rect 14464 43930 14516 43936
rect 14832 43852 14884 43858
rect 14832 43794 14884 43800
rect 14844 42702 14872 43794
rect 14924 43784 14976 43790
rect 14924 43726 14976 43732
rect 14936 43246 14964 43726
rect 14924 43240 14976 43246
rect 14924 43182 14976 43188
rect 14832 42696 14884 42702
rect 14832 42638 14884 42644
rect 14936 42634 14964 43182
rect 14924 42628 14976 42634
rect 14924 42570 14976 42576
rect 15028 42344 15056 44270
rect 15120 43926 15148 44338
rect 15108 43920 15160 43926
rect 15108 43862 15160 43868
rect 15212 43790 15240 44356
rect 15292 44338 15344 44344
rect 15476 44396 15528 44402
rect 15476 44338 15528 44344
rect 16040 43994 16068 44474
rect 16304 44464 16356 44470
rect 16304 44406 16356 44412
rect 16028 43988 16080 43994
rect 16028 43930 16080 43936
rect 16316 43790 16344 44406
rect 16500 44334 16528 44814
rect 16488 44328 16540 44334
rect 16488 44270 16540 44276
rect 16486 43888 16542 43897
rect 16486 43823 16542 43832
rect 16500 43790 16528 43823
rect 15200 43784 15252 43790
rect 15200 43726 15252 43732
rect 16304 43784 16356 43790
rect 16304 43726 16356 43732
rect 16488 43784 16540 43790
rect 16488 43726 16540 43732
rect 16580 43784 16632 43790
rect 16580 43726 16632 43732
rect 15212 43450 15240 43726
rect 15660 43716 15712 43722
rect 15660 43658 15712 43664
rect 15568 43648 15620 43654
rect 15568 43590 15620 43596
rect 15200 43444 15252 43450
rect 15200 43386 15252 43392
rect 15580 42702 15608 43590
rect 15672 43246 15700 43658
rect 15660 43240 15712 43246
rect 15660 43182 15712 43188
rect 15672 42906 15700 43182
rect 15844 43172 15896 43178
rect 15844 43114 15896 43120
rect 15660 42900 15712 42906
rect 15660 42842 15712 42848
rect 15856 42770 15884 43114
rect 16592 42838 16620 43726
rect 16764 43308 16816 43314
rect 16868 43296 16896 47058
rect 17040 47048 17092 47054
rect 17040 46990 17092 46996
rect 16948 46640 17000 46646
rect 16948 46582 17000 46588
rect 16960 43314 16988 46582
rect 17052 45082 17080 46990
rect 17420 46986 17448 49200
rect 19156 47728 19208 47734
rect 19156 47670 19208 47676
rect 17408 46980 17460 46986
rect 17408 46922 17460 46928
rect 18052 46572 18104 46578
rect 18052 46514 18104 46520
rect 18696 46572 18748 46578
rect 18696 46514 18748 46520
rect 18064 45830 18092 46514
rect 18512 46504 18564 46510
rect 18512 46446 18564 46452
rect 18236 46436 18288 46442
rect 18236 46378 18288 46384
rect 17684 45824 17736 45830
rect 17684 45766 17736 45772
rect 18052 45824 18104 45830
rect 18052 45766 18104 45772
rect 17696 45626 17724 45766
rect 17684 45620 17736 45626
rect 17684 45562 17736 45568
rect 18248 45490 18276 46378
rect 18420 46368 18472 46374
rect 18420 46310 18472 46316
rect 18432 46102 18460 46310
rect 18524 46170 18552 46446
rect 18708 46170 18736 46514
rect 18512 46164 18564 46170
rect 18512 46106 18564 46112
rect 18696 46164 18748 46170
rect 18696 46106 18748 46112
rect 18420 46096 18472 46102
rect 18420 46038 18472 46044
rect 18420 45892 18472 45898
rect 18420 45834 18472 45840
rect 18880 45892 18932 45898
rect 18880 45834 18932 45840
rect 18326 45520 18382 45529
rect 17592 45484 17644 45490
rect 17592 45426 17644 45432
rect 18236 45484 18288 45490
rect 18326 45455 18328 45464
rect 18236 45426 18288 45432
rect 18380 45455 18382 45464
rect 18328 45426 18380 45432
rect 17498 45384 17554 45393
rect 17498 45319 17554 45328
rect 17040 45076 17092 45082
rect 17040 45018 17092 45024
rect 17040 44940 17092 44946
rect 17040 44882 17092 44888
rect 17052 43314 17080 44882
rect 17512 44441 17540 45319
rect 17498 44432 17554 44441
rect 17498 44367 17500 44376
rect 17552 44367 17554 44376
rect 17500 44338 17552 44344
rect 16816 43268 16896 43296
rect 16764 43250 16816 43256
rect 16672 43104 16724 43110
rect 16672 43046 16724 43052
rect 16580 42832 16632 42838
rect 16580 42774 16632 42780
rect 15844 42764 15896 42770
rect 15844 42706 15896 42712
rect 15568 42696 15620 42702
rect 15568 42638 15620 42644
rect 15660 42560 15712 42566
rect 15660 42502 15712 42508
rect 15200 42356 15252 42362
rect 15028 42316 15200 42344
rect 15200 42298 15252 42304
rect 14740 41608 14792 41614
rect 14740 41550 14792 41556
rect 14108 41386 14320 41414
rect 14002 41304 14058 41313
rect 14002 41239 14058 41248
rect 14016 40474 14044 41239
rect 14108 40610 14136 41386
rect 14752 41274 14780 41550
rect 15108 41472 15160 41478
rect 15108 41414 15160 41420
rect 15212 41414 15240 42298
rect 15672 42226 15700 42502
rect 15660 42220 15712 42226
rect 15660 42162 15712 42168
rect 15568 41812 15620 41818
rect 15568 41754 15620 41760
rect 15120 41274 15148 41414
rect 15212 41386 15332 41414
rect 14740 41268 14792 41274
rect 14740 41210 14792 41216
rect 15108 41268 15160 41274
rect 15108 41210 15160 41216
rect 14108 40582 14228 40610
rect 14016 40446 14136 40474
rect 14004 40384 14056 40390
rect 14004 40326 14056 40332
rect 13912 40180 13964 40186
rect 13912 40122 13964 40128
rect 13820 39500 13872 39506
rect 13820 39442 13872 39448
rect 13636 39364 13688 39370
rect 13636 39306 13688 39312
rect 13648 39030 13676 39306
rect 13832 39098 13860 39442
rect 13820 39092 13872 39098
rect 13820 39034 13872 39040
rect 13636 39024 13688 39030
rect 13636 38966 13688 38972
rect 13452 38480 13504 38486
rect 13452 38422 13504 38428
rect 13464 37942 13492 38422
rect 13820 38276 13872 38282
rect 13820 38218 13872 38224
rect 13452 37936 13504 37942
rect 13452 37878 13504 37884
rect 13544 37936 13596 37942
rect 13544 37878 13596 37884
rect 13452 37256 13504 37262
rect 13452 37198 13504 37204
rect 13464 36786 13492 37198
rect 13556 36922 13584 37878
rect 13832 37466 13860 38218
rect 13912 37868 13964 37874
rect 13912 37810 13964 37816
rect 13820 37460 13872 37466
rect 13820 37402 13872 37408
rect 13924 37194 13952 37810
rect 13912 37188 13964 37194
rect 13912 37130 13964 37136
rect 13544 36916 13596 36922
rect 13544 36858 13596 36864
rect 13924 36854 13952 37130
rect 13912 36848 13964 36854
rect 13912 36790 13964 36796
rect 13452 36780 13504 36786
rect 13452 36722 13504 36728
rect 13544 36780 13596 36786
rect 13544 36722 13596 36728
rect 13556 35086 13584 36722
rect 13728 36032 13780 36038
rect 13728 35974 13780 35980
rect 13740 35562 13768 35974
rect 13820 35624 13872 35630
rect 13820 35566 13872 35572
rect 13728 35556 13780 35562
rect 13728 35498 13780 35504
rect 13544 35080 13596 35086
rect 13544 35022 13596 35028
rect 13832 34610 13860 35566
rect 13820 34604 13872 34610
rect 13820 34546 13872 34552
rect 13832 34066 13860 34546
rect 13820 34060 13872 34066
rect 13820 34002 13872 34008
rect 13452 33584 13504 33590
rect 13452 33526 13504 33532
rect 13464 32842 13492 33526
rect 13820 33516 13872 33522
rect 13820 33458 13872 33464
rect 13832 32910 13860 33458
rect 13820 32904 13872 32910
rect 13820 32846 13872 32852
rect 13452 32836 13504 32842
rect 13452 32778 13504 32784
rect 13464 31346 13492 32778
rect 13832 32502 13860 32846
rect 13820 32496 13872 32502
rect 13820 32438 13872 32444
rect 13544 32224 13596 32230
rect 13544 32166 13596 32172
rect 13556 31822 13584 32166
rect 13832 32042 13860 32438
rect 13648 32014 13860 32042
rect 13648 31822 13676 32014
rect 13728 31884 13780 31890
rect 13728 31826 13780 31832
rect 13544 31816 13596 31822
rect 13544 31758 13596 31764
rect 13636 31816 13688 31822
rect 13636 31758 13688 31764
rect 13740 31686 13768 31826
rect 13820 31816 13872 31822
rect 13820 31758 13872 31764
rect 13728 31680 13780 31686
rect 13728 31622 13780 31628
rect 13740 31346 13768 31622
rect 13832 31482 13860 31758
rect 13820 31476 13872 31482
rect 13820 31418 13872 31424
rect 13452 31340 13504 31346
rect 13452 31282 13504 31288
rect 13728 31340 13780 31346
rect 13728 31282 13780 31288
rect 13740 30938 13768 31282
rect 13728 30932 13780 30938
rect 13728 30874 13780 30880
rect 13832 30666 13860 31418
rect 13820 30660 13872 30666
rect 13820 30602 13872 30608
rect 14016 19718 14044 40326
rect 14108 38554 14136 40446
rect 14200 39914 14228 40582
rect 15120 40526 15148 41210
rect 15200 41132 15252 41138
rect 15200 41074 15252 41080
rect 15212 40662 15240 41074
rect 15200 40656 15252 40662
rect 15200 40598 15252 40604
rect 15016 40520 15068 40526
rect 15014 40488 15016 40497
rect 15108 40520 15160 40526
rect 15068 40488 15070 40497
rect 15108 40462 15160 40468
rect 15014 40423 15070 40432
rect 15304 40390 15332 41386
rect 15580 40730 15608 41754
rect 15672 41614 15700 42162
rect 15936 42152 15988 42158
rect 15936 42094 15988 42100
rect 15752 42016 15804 42022
rect 15752 41958 15804 41964
rect 15764 41818 15792 41958
rect 15752 41812 15804 41818
rect 15752 41754 15804 41760
rect 15948 41614 15976 42094
rect 15660 41608 15712 41614
rect 15660 41550 15712 41556
rect 15936 41608 15988 41614
rect 15936 41550 15988 41556
rect 15672 41206 15700 41550
rect 15660 41200 15712 41206
rect 15660 41142 15712 41148
rect 15948 41138 15976 41550
rect 16120 41540 16172 41546
rect 16120 41482 16172 41488
rect 16132 41274 16160 41482
rect 16120 41268 16172 41274
rect 16120 41210 16172 41216
rect 15936 41132 15988 41138
rect 15936 41074 15988 41080
rect 15660 41064 15712 41070
rect 15660 41006 15712 41012
rect 15568 40724 15620 40730
rect 15568 40666 15620 40672
rect 15292 40384 15344 40390
rect 15292 40326 15344 40332
rect 14832 40180 14884 40186
rect 14832 40122 14884 40128
rect 15476 40180 15528 40186
rect 15476 40122 15528 40128
rect 14648 40044 14700 40050
rect 14648 39986 14700 39992
rect 14280 39976 14332 39982
rect 14280 39918 14332 39924
rect 14188 39908 14240 39914
rect 14188 39850 14240 39856
rect 14292 39098 14320 39918
rect 14464 39500 14516 39506
rect 14464 39442 14516 39448
rect 14372 39364 14424 39370
rect 14372 39306 14424 39312
rect 14280 39092 14332 39098
rect 14280 39034 14332 39040
rect 14384 39030 14412 39306
rect 14188 39024 14240 39030
rect 14372 39024 14424 39030
rect 14240 38972 14320 38978
rect 14188 38966 14320 38972
rect 14372 38966 14424 38972
rect 14200 38950 14320 38966
rect 14476 38962 14504 39442
rect 14556 39296 14608 39302
rect 14556 39238 14608 39244
rect 14568 38962 14596 39238
rect 14292 38894 14320 38950
rect 14464 38956 14516 38962
rect 14464 38898 14516 38904
rect 14556 38956 14608 38962
rect 14556 38898 14608 38904
rect 14280 38888 14332 38894
rect 14280 38830 14332 38836
rect 14096 38548 14148 38554
rect 14096 38490 14148 38496
rect 14188 38004 14240 38010
rect 14188 37946 14240 37952
rect 14200 37262 14228 37946
rect 14292 37874 14320 38830
rect 14476 38554 14504 38898
rect 14464 38548 14516 38554
rect 14464 38490 14516 38496
rect 14660 38282 14688 39986
rect 14648 38276 14700 38282
rect 14648 38218 14700 38224
rect 14556 37936 14608 37942
rect 14556 37878 14608 37884
rect 14280 37868 14332 37874
rect 14280 37810 14332 37816
rect 14568 37777 14596 37878
rect 14554 37768 14610 37777
rect 14554 37703 14610 37712
rect 14188 37256 14240 37262
rect 14188 37198 14240 37204
rect 14096 37120 14148 37126
rect 14096 37062 14148 37068
rect 14108 36786 14136 37062
rect 14096 36780 14148 36786
rect 14096 36722 14148 36728
rect 14096 36100 14148 36106
rect 14096 36042 14148 36048
rect 14108 35494 14136 36042
rect 14096 35488 14148 35494
rect 14096 35430 14148 35436
rect 14108 35222 14136 35430
rect 14096 35216 14148 35222
rect 14096 35158 14148 35164
rect 14108 33454 14136 35158
rect 14096 33448 14148 33454
rect 14096 33390 14148 33396
rect 14200 32570 14228 37198
rect 14660 36922 14688 38218
rect 14844 37274 14872 40122
rect 15488 40089 15516 40122
rect 15474 40080 15530 40089
rect 15474 40015 15530 40024
rect 15016 39908 15068 39914
rect 15016 39850 15068 39856
rect 15028 38978 15056 39850
rect 15672 39846 15700 41006
rect 16592 40526 16620 42774
rect 16684 42226 16712 43046
rect 16764 42764 16816 42770
rect 16764 42706 16816 42712
rect 16672 42220 16724 42226
rect 16672 42162 16724 42168
rect 16776 42158 16804 42706
rect 16868 42702 16896 43268
rect 16948 43308 17000 43314
rect 16948 43250 17000 43256
rect 17040 43308 17092 43314
rect 17040 43250 17092 43256
rect 16856 42696 16908 42702
rect 16856 42638 16908 42644
rect 16960 42566 16988 43250
rect 17132 42628 17184 42634
rect 17132 42570 17184 42576
rect 16948 42560 17000 42566
rect 16948 42502 17000 42508
rect 16764 42152 16816 42158
rect 16764 42094 16816 42100
rect 16960 42106 16988 42502
rect 17144 42226 17172 42570
rect 17132 42220 17184 42226
rect 17132 42162 17184 42168
rect 16776 41614 16804 42094
rect 16960 42078 17172 42106
rect 16856 42016 16908 42022
rect 16856 41958 16908 41964
rect 16764 41608 16816 41614
rect 16764 41550 16816 41556
rect 16764 41472 16816 41478
rect 16764 41414 16816 41420
rect 16776 41070 16804 41414
rect 16868 41138 16896 41958
rect 16948 41608 17000 41614
rect 16948 41550 17000 41556
rect 16960 41274 16988 41550
rect 17144 41528 17172 42078
rect 17224 41540 17276 41546
rect 17144 41500 17224 41528
rect 16948 41268 17000 41274
rect 16948 41210 17000 41216
rect 16856 41132 16908 41138
rect 16856 41074 16908 41080
rect 16764 41064 16816 41070
rect 16764 41006 16816 41012
rect 16580 40520 16632 40526
rect 16580 40462 16632 40468
rect 17040 40384 17092 40390
rect 17040 40326 17092 40332
rect 17052 40186 17080 40326
rect 17040 40180 17092 40186
rect 17040 40122 17092 40128
rect 17144 39982 17172 41500
rect 17224 41482 17276 41488
rect 17604 41206 17632 45426
rect 17960 44736 18012 44742
rect 17960 44678 18012 44684
rect 17972 44146 18000 44678
rect 18142 44432 18198 44441
rect 18052 44396 18104 44402
rect 18142 44367 18144 44376
rect 18052 44338 18104 44344
rect 18196 44367 18198 44376
rect 18144 44338 18196 44344
rect 17880 44118 18000 44146
rect 17880 43858 17908 44118
rect 17960 43988 18012 43994
rect 17960 43930 18012 43936
rect 17868 43852 17920 43858
rect 17868 43794 17920 43800
rect 17972 43382 18000 43930
rect 18064 43432 18092 44338
rect 18156 43897 18184 44338
rect 18236 44192 18288 44198
rect 18236 44134 18288 44140
rect 18142 43888 18198 43897
rect 18142 43823 18198 43832
rect 18248 43790 18276 44134
rect 18236 43784 18288 43790
rect 18236 43726 18288 43732
rect 18340 43636 18368 45426
rect 18432 45422 18460 45834
rect 18604 45484 18656 45490
rect 18604 45426 18656 45432
rect 18420 45416 18472 45422
rect 18420 45358 18472 45364
rect 18248 43608 18368 43636
rect 18064 43404 18184 43432
rect 17960 43376 18012 43382
rect 18012 43324 18092 43330
rect 17960 43318 18092 43324
rect 17684 43308 17736 43314
rect 17972 43302 18092 43318
rect 17684 43250 17736 43256
rect 17696 41818 17724 43250
rect 17868 43240 17920 43246
rect 17866 43208 17868 43217
rect 17920 43208 17922 43217
rect 17866 43143 17922 43152
rect 17960 43172 18012 43178
rect 17960 43114 18012 43120
rect 17972 42702 18000 43114
rect 17960 42696 18012 42702
rect 17960 42638 18012 42644
rect 17960 42560 18012 42566
rect 17960 42502 18012 42508
rect 17972 42226 18000 42502
rect 17960 42220 18012 42226
rect 17960 42162 18012 42168
rect 17684 41812 17736 41818
rect 17684 41754 17736 41760
rect 17972 41478 18000 42162
rect 17960 41472 18012 41478
rect 17960 41414 18012 41420
rect 17972 41290 18000 41414
rect 17880 41262 18000 41290
rect 17592 41200 17644 41206
rect 17592 41142 17644 41148
rect 17604 40662 17632 41142
rect 17880 40730 17908 41262
rect 18064 41154 18092 43302
rect 18156 42702 18184 43404
rect 18144 42696 18196 42702
rect 18144 42638 18196 42644
rect 18156 42294 18184 42638
rect 18144 42288 18196 42294
rect 18144 42230 18196 42236
rect 18144 41268 18196 41274
rect 18144 41210 18196 41216
rect 17972 41126 18092 41154
rect 18156 41138 18184 41210
rect 18144 41132 18196 41138
rect 17868 40724 17920 40730
rect 17868 40666 17920 40672
rect 17592 40656 17644 40662
rect 17592 40598 17644 40604
rect 17604 40118 17632 40598
rect 17868 40520 17920 40526
rect 17866 40488 17868 40497
rect 17920 40488 17922 40497
rect 17866 40423 17922 40432
rect 17224 40112 17276 40118
rect 17592 40112 17644 40118
rect 17224 40054 17276 40060
rect 17406 40080 17462 40089
rect 17040 39976 17092 39982
rect 17040 39918 17092 39924
rect 17132 39976 17184 39982
rect 17132 39918 17184 39924
rect 15660 39840 15712 39846
rect 15660 39782 15712 39788
rect 16304 39840 16356 39846
rect 16304 39782 16356 39788
rect 15028 38962 15424 38978
rect 15016 38956 15436 38962
rect 15068 38950 15384 38956
rect 15016 38898 15068 38904
rect 15384 38898 15436 38904
rect 15028 37754 15056 38898
rect 15672 38486 15700 39782
rect 15752 39432 15804 39438
rect 15752 39374 15804 39380
rect 16120 39432 16172 39438
rect 16120 39374 16172 39380
rect 15660 38480 15712 38486
rect 15660 38422 15712 38428
rect 15764 38418 15792 39374
rect 16132 39098 16160 39374
rect 16212 39296 16264 39302
rect 16212 39238 16264 39244
rect 15844 39092 15896 39098
rect 15844 39034 15896 39040
rect 16120 39092 16172 39098
rect 16120 39034 16172 39040
rect 15856 38876 15884 39034
rect 16028 38956 16080 38962
rect 16028 38898 16080 38904
rect 15936 38888 15988 38894
rect 15856 38848 15936 38876
rect 15936 38830 15988 38836
rect 16040 38486 16068 38898
rect 16028 38480 16080 38486
rect 16028 38422 16080 38428
rect 15752 38412 15804 38418
rect 15752 38354 15804 38360
rect 15108 38344 15160 38350
rect 15292 38344 15344 38350
rect 15160 38292 15240 38298
rect 15108 38286 15240 38292
rect 15292 38286 15344 38292
rect 15120 38270 15240 38286
rect 15212 37874 15240 38270
rect 15200 37868 15252 37874
rect 15200 37810 15252 37816
rect 14936 37738 15056 37754
rect 14924 37732 15056 37738
rect 14976 37726 15056 37732
rect 14924 37674 14976 37680
rect 15028 37482 15056 37726
rect 15106 37496 15162 37505
rect 15028 37454 15106 37482
rect 15212 37466 15240 37810
rect 15304 37806 15332 38286
rect 15476 38276 15528 38282
rect 15476 38218 15528 38224
rect 15488 37874 15516 38218
rect 15476 37868 15528 37874
rect 15476 37810 15528 37816
rect 15292 37800 15344 37806
rect 15292 37742 15344 37748
rect 15106 37431 15162 37440
rect 15200 37460 15252 37466
rect 14844 37246 14964 37274
rect 14648 36916 14700 36922
rect 14648 36858 14700 36864
rect 14280 35692 14332 35698
rect 14280 35634 14332 35640
rect 14292 34542 14320 35634
rect 14464 35488 14516 35494
rect 14464 35430 14516 35436
rect 14476 34610 14504 35430
rect 14556 34944 14608 34950
rect 14556 34886 14608 34892
rect 14568 34746 14596 34886
rect 14556 34740 14608 34746
rect 14556 34682 14608 34688
rect 14464 34604 14516 34610
rect 14464 34546 14516 34552
rect 14740 34604 14792 34610
rect 14740 34546 14792 34552
rect 14280 34536 14332 34542
rect 14280 34478 14332 34484
rect 14292 33998 14320 34478
rect 14280 33992 14332 33998
rect 14280 33934 14332 33940
rect 14476 33862 14504 34546
rect 14752 34202 14780 34546
rect 14832 34400 14884 34406
rect 14832 34342 14884 34348
rect 14740 34196 14792 34202
rect 14740 34138 14792 34144
rect 14844 33998 14872 34342
rect 14832 33992 14884 33998
rect 14832 33934 14884 33940
rect 14464 33856 14516 33862
rect 14464 33798 14516 33804
rect 14476 33522 14504 33798
rect 14464 33516 14516 33522
rect 14464 33458 14516 33464
rect 14740 32768 14792 32774
rect 14740 32710 14792 32716
rect 14188 32564 14240 32570
rect 14188 32506 14240 32512
rect 14200 32366 14228 32506
rect 14752 32366 14780 32710
rect 14188 32360 14240 32366
rect 14740 32360 14792 32366
rect 14240 32320 14412 32348
rect 14188 32302 14240 32308
rect 14188 31816 14240 31822
rect 14188 31758 14240 31764
rect 14200 31278 14228 31758
rect 14384 31754 14412 32320
rect 14740 32302 14792 32308
rect 14832 32224 14884 32230
rect 14832 32166 14884 32172
rect 14844 31822 14872 32166
rect 14832 31816 14884 31822
rect 14832 31758 14884 31764
rect 14384 31726 14596 31754
rect 14188 31272 14240 31278
rect 14188 31214 14240 31220
rect 14004 19712 14056 19718
rect 14004 19654 14056 19660
rect 14568 2582 14596 31726
rect 14832 31340 14884 31346
rect 14832 31282 14884 31288
rect 14844 30802 14872 31282
rect 14832 30796 14884 30802
rect 14832 30738 14884 30744
rect 14832 29028 14884 29034
rect 14832 28970 14884 28976
rect 14556 2576 14608 2582
rect 14556 2518 14608 2524
rect 14844 2446 14872 28970
rect 14936 7886 14964 37246
rect 15016 37256 15068 37262
rect 15014 37224 15016 37233
rect 15068 37224 15070 37233
rect 15014 37159 15070 37168
rect 15120 36786 15148 37431
rect 15200 37402 15252 37408
rect 15212 37126 15240 37402
rect 15200 37120 15252 37126
rect 15200 37062 15252 37068
rect 15108 36780 15160 36786
rect 15108 36722 15160 36728
rect 15304 36650 15332 37742
rect 15764 37670 15792 38354
rect 16040 38214 16068 38422
rect 16224 38282 16252 39238
rect 16212 38276 16264 38282
rect 16212 38218 16264 38224
rect 16028 38208 16080 38214
rect 16028 38150 16080 38156
rect 16120 38208 16172 38214
rect 16120 38150 16172 38156
rect 16132 37670 16160 38150
rect 15752 37664 15804 37670
rect 15752 37606 15804 37612
rect 16028 37664 16080 37670
rect 16028 37606 16080 37612
rect 16120 37664 16172 37670
rect 16120 37606 16172 37612
rect 15934 37360 15990 37369
rect 15934 37295 15990 37304
rect 15384 37256 15436 37262
rect 15384 37198 15436 37204
rect 15396 36854 15424 37198
rect 15384 36848 15436 36854
rect 15384 36790 15436 36796
rect 15842 36680 15898 36689
rect 15292 36644 15344 36650
rect 15842 36615 15898 36624
rect 15292 36586 15344 36592
rect 15856 36582 15884 36615
rect 15844 36576 15896 36582
rect 15844 36518 15896 36524
rect 15948 36378 15976 37295
rect 16040 36564 16068 37606
rect 16316 37398 16344 39782
rect 17052 39642 17080 39918
rect 17236 39846 17264 40054
rect 17592 40054 17644 40060
rect 17972 40066 18000 41126
rect 18144 41074 18196 41080
rect 18156 40526 18184 41074
rect 18144 40520 18196 40526
rect 18144 40462 18196 40468
rect 17972 40038 18092 40066
rect 17406 40015 17462 40024
rect 17420 39982 17448 40015
rect 17408 39976 17460 39982
rect 17408 39918 17460 39924
rect 18064 39846 18092 40038
rect 17224 39840 17276 39846
rect 17224 39782 17276 39788
rect 18052 39840 18104 39846
rect 18052 39782 18104 39788
rect 16948 39636 17000 39642
rect 16948 39578 17000 39584
rect 17040 39636 17092 39642
rect 17040 39578 17092 39584
rect 16960 39438 16988 39578
rect 17960 39500 18012 39506
rect 17960 39442 18012 39448
rect 16396 39432 16448 39438
rect 16396 39374 16448 39380
rect 16948 39432 17000 39438
rect 16948 39374 17000 39380
rect 17776 39432 17828 39438
rect 17776 39374 17828 39380
rect 16408 38894 16436 39374
rect 17316 39364 17368 39370
rect 17316 39306 17368 39312
rect 16396 38888 16448 38894
rect 16396 38830 16448 38836
rect 17040 38752 17092 38758
rect 17040 38694 17092 38700
rect 17052 38554 17080 38694
rect 16672 38548 16724 38554
rect 16672 38490 16724 38496
rect 17040 38548 17092 38554
rect 17040 38490 17092 38496
rect 16488 38412 16540 38418
rect 16488 38354 16540 38360
rect 16500 37942 16528 38354
rect 16488 37936 16540 37942
rect 16488 37878 16540 37884
rect 16500 37466 16528 37878
rect 16684 37874 16712 38490
rect 16856 38344 16908 38350
rect 16856 38286 16908 38292
rect 16868 38010 16896 38286
rect 17040 38208 17092 38214
rect 17040 38150 17092 38156
rect 16856 38004 16908 38010
rect 16856 37946 16908 37952
rect 17052 37913 17080 38150
rect 17224 38004 17276 38010
rect 17224 37946 17276 37952
rect 17038 37904 17094 37913
rect 16672 37868 16724 37874
rect 16672 37810 16724 37816
rect 16948 37868 17000 37874
rect 17038 37839 17094 37848
rect 16948 37810 17000 37816
rect 16578 37632 16634 37641
rect 16578 37567 16634 37576
rect 16488 37460 16540 37466
rect 16488 37402 16540 37408
rect 16304 37392 16356 37398
rect 16304 37334 16356 37340
rect 16120 36576 16172 36582
rect 16040 36544 16120 36564
rect 16172 36544 16174 36553
rect 16040 36536 16118 36544
rect 15936 36372 15988 36378
rect 15936 36314 15988 36320
rect 15568 36236 15620 36242
rect 15568 36178 15620 36184
rect 15384 35692 15436 35698
rect 15384 35634 15436 35640
rect 15396 34950 15424 35634
rect 15476 35624 15528 35630
rect 15476 35566 15528 35572
rect 15488 35068 15516 35566
rect 15580 35290 15608 36178
rect 15660 36168 15712 36174
rect 15660 36110 15712 36116
rect 15568 35284 15620 35290
rect 15568 35226 15620 35232
rect 15568 35080 15620 35086
rect 15488 35040 15568 35068
rect 15568 35022 15620 35028
rect 15384 34944 15436 34950
rect 15384 34886 15436 34892
rect 15292 34536 15344 34542
rect 15292 34478 15344 34484
rect 15016 33992 15068 33998
rect 15016 33934 15068 33940
rect 15028 33522 15056 33934
rect 15304 33522 15332 34478
rect 15384 34468 15436 34474
rect 15384 34410 15436 34416
rect 15396 33980 15424 34410
rect 15580 34202 15608 35022
rect 15672 34746 15700 36110
rect 16040 36106 16068 36536
rect 16118 36479 16174 36488
rect 16592 36106 16620 37567
rect 16960 37466 16988 37810
rect 17236 37738 17264 37946
rect 17224 37732 17276 37738
rect 17224 37674 17276 37680
rect 16948 37460 17000 37466
rect 16948 37402 17000 37408
rect 16948 37324 17000 37330
rect 16948 37266 17000 37272
rect 16960 37126 16988 37266
rect 17224 37188 17276 37194
rect 17224 37130 17276 37136
rect 16948 37120 17000 37126
rect 16948 37062 17000 37068
rect 16856 36916 16908 36922
rect 16856 36858 16908 36864
rect 16868 36174 16896 36858
rect 16960 36582 16988 37062
rect 16948 36576 17000 36582
rect 16948 36518 17000 36524
rect 16856 36168 16908 36174
rect 16856 36110 16908 36116
rect 16028 36100 16080 36106
rect 16028 36042 16080 36048
rect 16580 36100 16632 36106
rect 16580 36042 16632 36048
rect 16592 35698 16620 36042
rect 16672 36032 16724 36038
rect 16672 35974 16724 35980
rect 16580 35692 16632 35698
rect 16580 35634 16632 35640
rect 15844 35148 15896 35154
rect 15844 35090 15896 35096
rect 15660 34740 15712 34746
rect 15712 34700 15792 34728
rect 15660 34682 15712 34688
rect 15568 34196 15620 34202
rect 15568 34138 15620 34144
rect 15476 33992 15528 33998
rect 15396 33952 15476 33980
rect 15396 33658 15424 33952
rect 15476 33934 15528 33940
rect 15384 33652 15436 33658
rect 15384 33594 15436 33600
rect 15016 33516 15068 33522
rect 15016 33458 15068 33464
rect 15292 33516 15344 33522
rect 15292 33458 15344 33464
rect 15660 33516 15712 33522
rect 15660 33458 15712 33464
rect 15304 32994 15332 33458
rect 15568 33312 15620 33318
rect 15568 33254 15620 33260
rect 15212 32966 15332 32994
rect 15212 32230 15240 32966
rect 15580 32910 15608 33254
rect 15292 32904 15344 32910
rect 15292 32846 15344 32852
rect 15568 32904 15620 32910
rect 15568 32846 15620 32852
rect 15304 32502 15332 32846
rect 15292 32496 15344 32502
rect 15292 32438 15344 32444
rect 15200 32224 15252 32230
rect 15200 32166 15252 32172
rect 15672 32026 15700 33458
rect 15764 32978 15792 34700
rect 15856 34610 15884 35090
rect 16684 35086 16712 35974
rect 16868 35698 16896 36110
rect 16856 35692 16908 35698
rect 16856 35634 16908 35640
rect 16672 35080 16724 35086
rect 16672 35022 16724 35028
rect 15936 34944 15988 34950
rect 15936 34886 15988 34892
rect 15844 34604 15896 34610
rect 15844 34546 15896 34552
rect 15752 32972 15804 32978
rect 15752 32914 15804 32920
rect 15948 32910 15976 34886
rect 16856 34740 16908 34746
rect 16856 34682 16908 34688
rect 16580 34672 16632 34678
rect 16580 34614 16632 34620
rect 16592 33998 16620 34614
rect 16672 34536 16724 34542
rect 16672 34478 16724 34484
rect 16764 34536 16816 34542
rect 16764 34478 16816 34484
rect 16684 34134 16712 34478
rect 16672 34128 16724 34134
rect 16672 34070 16724 34076
rect 16580 33992 16632 33998
rect 16580 33934 16632 33940
rect 16776 33386 16804 34478
rect 16868 34202 16896 34682
rect 16856 34196 16908 34202
rect 16856 34138 16908 34144
rect 16580 33380 16632 33386
rect 16580 33322 16632 33328
rect 16764 33380 16816 33386
rect 16764 33322 16816 33328
rect 15936 32904 15988 32910
rect 15936 32846 15988 32852
rect 16592 32026 16620 33322
rect 16672 32904 16724 32910
rect 16672 32846 16724 32852
rect 16684 32570 16712 32846
rect 16672 32564 16724 32570
rect 16672 32506 16724 32512
rect 16856 32428 16908 32434
rect 16856 32370 16908 32376
rect 16672 32292 16724 32298
rect 16672 32234 16724 32240
rect 15660 32020 15712 32026
rect 15660 31962 15712 31968
rect 16580 32020 16632 32026
rect 16580 31962 16632 31968
rect 15200 31952 15252 31958
rect 15200 31894 15252 31900
rect 15016 31748 15068 31754
rect 15016 31690 15068 31696
rect 15028 31482 15056 31690
rect 15212 31482 15240 31894
rect 15382 31784 15438 31793
rect 15382 31719 15384 31728
rect 15436 31719 15438 31728
rect 15384 31690 15436 31696
rect 15016 31476 15068 31482
rect 15016 31418 15068 31424
rect 15200 31476 15252 31482
rect 15200 31418 15252 31424
rect 16488 31476 16540 31482
rect 16488 31418 16540 31424
rect 15844 31408 15896 31414
rect 15028 31346 15332 31362
rect 15844 31350 15896 31356
rect 15016 31340 15332 31346
rect 15068 31334 15332 31340
rect 15016 31282 15068 31288
rect 15200 31272 15252 31278
rect 15200 31214 15252 31220
rect 15212 30938 15240 31214
rect 15200 30932 15252 30938
rect 15200 30874 15252 30880
rect 15304 30666 15332 31334
rect 15568 30864 15620 30870
rect 15568 30806 15620 30812
rect 15292 30660 15344 30666
rect 15292 30602 15344 30608
rect 15304 30258 15332 30602
rect 15384 30388 15436 30394
rect 15384 30330 15436 30336
rect 15292 30252 15344 30258
rect 15292 30194 15344 30200
rect 15304 29782 15332 30194
rect 15396 29850 15424 30330
rect 15580 30258 15608 30806
rect 15856 30666 15884 31350
rect 16500 31142 16528 31418
rect 16396 31136 16448 31142
rect 16396 31078 16448 31084
rect 16488 31136 16540 31142
rect 16488 31078 16540 31084
rect 15844 30660 15896 30666
rect 15844 30602 15896 30608
rect 16028 30660 16080 30666
rect 16028 30602 16080 30608
rect 15856 30394 15884 30602
rect 15844 30388 15896 30394
rect 15844 30330 15896 30336
rect 15568 30252 15620 30258
rect 15568 30194 15620 30200
rect 16040 29850 16068 30602
rect 16304 30252 16356 30258
rect 16304 30194 16356 30200
rect 15384 29844 15436 29850
rect 15384 29786 15436 29792
rect 16028 29844 16080 29850
rect 16028 29786 16080 29792
rect 15292 29776 15344 29782
rect 15292 29718 15344 29724
rect 15304 28014 15332 29718
rect 15396 28762 15424 29786
rect 16316 29782 16344 30194
rect 16304 29776 16356 29782
rect 16304 29718 16356 29724
rect 16408 29696 16436 31078
rect 16684 30258 16712 32234
rect 16868 30938 16896 32370
rect 16960 32212 16988 36518
rect 17236 36242 17264 37130
rect 17224 36236 17276 36242
rect 17224 36178 17276 36184
rect 17224 35692 17276 35698
rect 17224 35634 17276 35640
rect 17040 35148 17092 35154
rect 17040 35090 17092 35096
rect 17052 32910 17080 35090
rect 17132 35080 17184 35086
rect 17132 35022 17184 35028
rect 17144 33114 17172 35022
rect 17132 33108 17184 33114
rect 17132 33050 17184 33056
rect 17040 32904 17092 32910
rect 17040 32846 17092 32852
rect 17040 32224 17092 32230
rect 16960 32184 17040 32212
rect 17040 32166 17092 32172
rect 16856 30932 16908 30938
rect 16856 30874 16908 30880
rect 16856 30728 16908 30734
rect 16856 30670 16908 30676
rect 16672 30252 16724 30258
rect 16672 30194 16724 30200
rect 16580 30184 16632 30190
rect 16580 30126 16632 30132
rect 16488 29708 16540 29714
rect 16408 29668 16488 29696
rect 16488 29650 16540 29656
rect 16592 29578 16620 30126
rect 16580 29572 16632 29578
rect 16580 29514 16632 29520
rect 15476 29504 15528 29510
rect 15476 29446 15528 29452
rect 15488 29034 15516 29446
rect 16120 29164 16172 29170
rect 16120 29106 16172 29112
rect 15476 29028 15528 29034
rect 15476 28970 15528 28976
rect 15384 28756 15436 28762
rect 15384 28698 15436 28704
rect 15292 28008 15344 28014
rect 15292 27950 15344 27956
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 15488 3466 15516 28970
rect 16132 28422 16160 29106
rect 16684 28558 16712 30194
rect 16868 29646 16896 30670
rect 16948 30252 17000 30258
rect 16948 30194 17000 30200
rect 16960 29850 16988 30194
rect 16948 29844 17000 29850
rect 16948 29786 17000 29792
rect 17052 29730 17080 32166
rect 17144 31822 17172 33050
rect 17132 31816 17184 31822
rect 17132 31758 17184 31764
rect 16960 29702 17080 29730
rect 16856 29640 16908 29646
rect 16856 29582 16908 29588
rect 16868 29306 16896 29582
rect 16856 29300 16908 29306
rect 16856 29242 16908 29248
rect 16960 29034 16988 29702
rect 17040 29640 17092 29646
rect 17040 29582 17092 29588
rect 17052 29306 17080 29582
rect 17040 29300 17092 29306
rect 17040 29242 17092 29248
rect 17236 29170 17264 35634
rect 17328 34474 17356 39306
rect 17788 39098 17816 39374
rect 17776 39092 17828 39098
rect 17776 39034 17828 39040
rect 17592 38344 17644 38350
rect 17590 38312 17592 38321
rect 17644 38312 17646 38321
rect 17590 38247 17646 38256
rect 17972 38214 18000 39442
rect 18064 39438 18092 39782
rect 18052 39432 18104 39438
rect 18052 39374 18104 39380
rect 18248 38842 18276 43608
rect 18616 43466 18644 45426
rect 18694 43752 18750 43761
rect 18694 43687 18696 43696
rect 18748 43687 18750 43696
rect 18696 43658 18748 43664
rect 18616 43438 18736 43466
rect 18326 43344 18382 43353
rect 18326 43279 18328 43288
rect 18380 43279 18382 43288
rect 18512 43308 18564 43314
rect 18328 43250 18380 43256
rect 18512 43250 18564 43256
rect 18340 42158 18368 43250
rect 18524 42906 18552 43250
rect 18604 43172 18656 43178
rect 18604 43114 18656 43120
rect 18512 42900 18564 42906
rect 18512 42842 18564 42848
rect 18512 42628 18564 42634
rect 18512 42570 18564 42576
rect 18328 42152 18380 42158
rect 18328 42094 18380 42100
rect 18420 42152 18472 42158
rect 18420 42094 18472 42100
rect 18432 41818 18460 42094
rect 18420 41812 18472 41818
rect 18420 41754 18472 41760
rect 18524 41614 18552 42570
rect 18512 41608 18564 41614
rect 18512 41550 18564 41556
rect 18420 41540 18472 41546
rect 18420 41482 18472 41488
rect 18432 41138 18460 41482
rect 18616 41177 18644 43114
rect 18602 41168 18658 41177
rect 18420 41132 18472 41138
rect 18602 41103 18658 41112
rect 18420 41074 18472 41080
rect 18328 41064 18380 41070
rect 18328 41006 18380 41012
rect 18340 40594 18368 41006
rect 18432 40662 18460 41074
rect 18512 40996 18564 41002
rect 18512 40938 18564 40944
rect 18420 40656 18472 40662
rect 18420 40598 18472 40604
rect 18328 40588 18380 40594
rect 18328 40530 18380 40536
rect 18524 40526 18552 40938
rect 18708 40730 18736 43438
rect 18788 42560 18840 42566
rect 18788 42502 18840 42508
rect 18800 42090 18828 42502
rect 18788 42084 18840 42090
rect 18788 42026 18840 42032
rect 18800 41682 18828 42026
rect 18788 41676 18840 41682
rect 18788 41618 18840 41624
rect 18892 41206 18920 45834
rect 19168 45354 19196 47670
rect 19352 47036 19380 49200
rect 21088 47796 21140 47802
rect 21088 47738 21140 47744
rect 19616 47592 19668 47598
rect 19616 47534 19668 47540
rect 19628 47258 19656 47534
rect 19616 47252 19668 47258
rect 19616 47194 19668 47200
rect 21100 47190 21128 47738
rect 21180 47660 21232 47666
rect 21180 47602 21232 47608
rect 21192 47258 21220 47602
rect 21180 47252 21232 47258
rect 21180 47194 21232 47200
rect 21088 47184 21140 47190
rect 21088 47126 21140 47132
rect 20260 47116 20312 47122
rect 20260 47058 20312 47064
rect 19432 47048 19484 47054
rect 19352 47008 19432 47036
rect 19432 46990 19484 46996
rect 19444 46714 19472 46990
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 19432 46708 19484 46714
rect 19432 46650 19484 46656
rect 19340 46640 19392 46646
rect 19340 46582 19392 46588
rect 19352 45529 19380 46582
rect 20076 46572 20128 46578
rect 20076 46514 20128 46520
rect 19982 46472 20038 46481
rect 19982 46407 19984 46416
rect 20036 46407 20038 46416
rect 19984 46378 20036 46384
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 19338 45520 19394 45529
rect 19338 45455 19394 45464
rect 19352 45354 19380 45455
rect 19156 45348 19208 45354
rect 19156 45290 19208 45296
rect 19340 45348 19392 45354
rect 19340 45290 19392 45296
rect 19248 44872 19300 44878
rect 19248 44814 19300 44820
rect 19156 44736 19208 44742
rect 19156 44678 19208 44684
rect 18972 44328 19024 44334
rect 18972 44270 19024 44276
rect 18984 43994 19012 44270
rect 18972 43988 19024 43994
rect 18972 43930 19024 43936
rect 19168 41682 19196 44678
rect 19260 44538 19288 44814
rect 19340 44736 19392 44742
rect 19340 44678 19392 44684
rect 19248 44532 19300 44538
rect 19248 44474 19300 44480
rect 19248 44396 19300 44402
rect 19248 44338 19300 44344
rect 19260 43450 19288 44338
rect 19248 43444 19300 43450
rect 19248 43386 19300 43392
rect 19352 42702 19380 44678
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19432 43716 19484 43722
rect 19432 43658 19484 43664
rect 19444 43330 19472 43658
rect 19984 43648 20036 43654
rect 19984 43590 20036 43596
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19444 43302 19564 43330
rect 19432 43240 19484 43246
rect 19432 43182 19484 43188
rect 19340 42696 19392 42702
rect 19340 42638 19392 42644
rect 19352 42226 19380 42638
rect 19340 42220 19392 42226
rect 19340 42162 19392 42168
rect 19340 42084 19392 42090
rect 19340 42026 19392 42032
rect 19156 41676 19208 41682
rect 19156 41618 19208 41624
rect 18880 41200 18932 41206
rect 18880 41142 18932 41148
rect 19352 41154 19380 42026
rect 19444 41818 19472 43182
rect 19536 42906 19564 43302
rect 19996 43246 20024 43590
rect 19984 43240 20036 43246
rect 19984 43182 20036 43188
rect 19984 43104 20036 43110
rect 19984 43046 20036 43052
rect 19524 42900 19576 42906
rect 19524 42842 19576 42848
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 19996 42294 20024 43046
rect 19984 42288 20036 42294
rect 19984 42230 20036 42236
rect 19996 42090 20024 42230
rect 19984 42084 20036 42090
rect 19984 42026 20036 42032
rect 19432 41812 19484 41818
rect 19432 41754 19484 41760
rect 19432 41608 19484 41614
rect 19432 41550 19484 41556
rect 19444 41449 19472 41550
rect 19430 41440 19486 41449
rect 19430 41375 19486 41384
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19708 41268 19760 41274
rect 19760 41228 19932 41256
rect 19708 41210 19760 41216
rect 18696 40724 18748 40730
rect 18696 40666 18748 40672
rect 18788 40724 18840 40730
rect 18788 40666 18840 40672
rect 18512 40520 18564 40526
rect 18512 40462 18564 40468
rect 18800 40458 18828 40666
rect 18892 40526 18920 41142
rect 19352 41138 19656 41154
rect 19064 41132 19116 41138
rect 19064 41074 19116 41080
rect 19248 41132 19300 41138
rect 19352 41132 19668 41138
rect 19352 41126 19616 41132
rect 19248 41074 19300 41080
rect 19616 41074 19668 41080
rect 19076 40594 19104 41074
rect 19260 40934 19288 41074
rect 19432 41064 19484 41070
rect 19432 41006 19484 41012
rect 19156 40928 19208 40934
rect 19156 40870 19208 40876
rect 19248 40928 19300 40934
rect 19248 40870 19300 40876
rect 19064 40588 19116 40594
rect 19064 40530 19116 40536
rect 18880 40520 18932 40526
rect 18880 40462 18932 40468
rect 18328 40452 18380 40458
rect 18328 40394 18380 40400
rect 18788 40452 18840 40458
rect 18788 40394 18840 40400
rect 18340 39914 18368 40394
rect 18892 39982 18920 40462
rect 19076 40390 19104 40530
rect 19064 40384 19116 40390
rect 19064 40326 19116 40332
rect 19168 40118 19196 40870
rect 19444 40730 19472 41006
rect 19432 40724 19484 40730
rect 19432 40666 19484 40672
rect 19338 40216 19394 40225
rect 19338 40151 19394 40160
rect 19352 40118 19380 40151
rect 19156 40112 19208 40118
rect 19156 40054 19208 40060
rect 19340 40112 19392 40118
rect 19340 40054 19392 40060
rect 18880 39976 18932 39982
rect 19444 39953 19472 40666
rect 19524 40656 19576 40662
rect 19524 40598 19576 40604
rect 19536 40390 19564 40598
rect 19800 40588 19852 40594
rect 19800 40530 19852 40536
rect 19812 40390 19840 40530
rect 19524 40384 19576 40390
rect 19524 40326 19576 40332
rect 19800 40384 19852 40390
rect 19904 40372 19932 41228
rect 19996 41206 20024 42026
rect 20088 41274 20116 46514
rect 20168 45892 20220 45898
rect 20168 45834 20220 45840
rect 20180 44402 20208 45834
rect 20168 44396 20220 44402
rect 20168 44338 20220 44344
rect 20076 41268 20128 41274
rect 20076 41210 20128 41216
rect 19984 41200 20036 41206
rect 19984 41142 20036 41148
rect 20076 40996 20128 41002
rect 20076 40938 20128 40944
rect 20088 40730 20116 40938
rect 20076 40724 20128 40730
rect 20076 40666 20128 40672
rect 20076 40588 20128 40594
rect 20076 40530 20128 40536
rect 19904 40344 20024 40372
rect 19800 40326 19852 40332
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19996 39982 20024 40344
rect 20088 40118 20116 40530
rect 20272 40186 20300 47058
rect 21284 46986 21312 49200
rect 22008 47524 22060 47530
rect 22008 47466 22060 47472
rect 21732 47048 21784 47054
rect 21732 46990 21784 46996
rect 20352 46980 20404 46986
rect 20352 46922 20404 46928
rect 20996 46980 21048 46986
rect 20996 46922 21048 46928
rect 21272 46980 21324 46986
rect 21272 46922 21324 46928
rect 20364 44334 20392 46922
rect 20812 46912 20864 46918
rect 20812 46854 20864 46860
rect 20718 46608 20774 46617
rect 20718 46543 20720 46552
rect 20772 46543 20774 46552
rect 20720 46514 20772 46520
rect 20732 45558 20760 46514
rect 20720 45552 20772 45558
rect 20720 45494 20772 45500
rect 20824 45490 20852 46854
rect 20904 46708 20956 46714
rect 20904 46650 20956 46656
rect 20916 46034 20944 46650
rect 21008 46374 21036 46922
rect 21640 46640 21692 46646
rect 21640 46582 21692 46588
rect 21180 46572 21232 46578
rect 21180 46514 21232 46520
rect 20996 46368 21048 46374
rect 20996 46310 21048 46316
rect 20904 46028 20956 46034
rect 20904 45970 20956 45976
rect 20996 45552 21048 45558
rect 20916 45512 20996 45540
rect 20812 45484 20864 45490
rect 20812 45426 20864 45432
rect 20444 45280 20496 45286
rect 20444 45222 20496 45228
rect 20456 44946 20484 45222
rect 20536 45076 20588 45082
rect 20536 45018 20588 45024
rect 20444 44940 20496 44946
rect 20444 44882 20496 44888
rect 20548 44878 20576 45018
rect 20916 44878 20944 45512
rect 20996 45494 21048 45500
rect 21088 45484 21140 45490
rect 21192 45472 21220 46514
rect 21456 45824 21508 45830
rect 21456 45766 21508 45772
rect 21140 45444 21312 45472
rect 21088 45426 21140 45432
rect 20996 45416 21048 45422
rect 21100 45393 21128 45426
rect 20996 45358 21048 45364
rect 21086 45384 21142 45393
rect 20536 44872 20588 44878
rect 20536 44814 20588 44820
rect 20904 44872 20956 44878
rect 20904 44814 20956 44820
rect 21008 44742 21036 45358
rect 21086 45319 21142 45328
rect 21180 45348 21232 45354
rect 21180 45290 21232 45296
rect 20720 44736 20772 44742
rect 20996 44736 21048 44742
rect 20772 44684 20852 44690
rect 20720 44678 20852 44684
rect 21048 44684 21128 44690
rect 20996 44678 21128 44684
rect 20732 44662 20852 44678
rect 21008 44662 21128 44678
rect 20718 44568 20774 44577
rect 20718 44503 20774 44512
rect 20732 44402 20760 44503
rect 20720 44396 20772 44402
rect 20720 44338 20772 44344
rect 20352 44328 20404 44334
rect 20352 44270 20404 44276
rect 20824 44198 20852 44662
rect 20812 44192 20864 44198
rect 20812 44134 20864 44140
rect 20536 43988 20588 43994
rect 20536 43930 20588 43936
rect 20628 43988 20680 43994
rect 20628 43930 20680 43936
rect 20352 43240 20404 43246
rect 20352 43182 20404 43188
rect 20364 42770 20392 43182
rect 20352 42764 20404 42770
rect 20352 42706 20404 42712
rect 20548 42362 20576 43930
rect 20640 43382 20668 43930
rect 20824 43926 20852 44134
rect 20812 43920 20864 43926
rect 20812 43862 20864 43868
rect 20720 43648 20772 43654
rect 20720 43590 20772 43596
rect 20628 43376 20680 43382
rect 20628 43318 20680 43324
rect 20732 43314 20760 43590
rect 20824 43382 20852 43862
rect 20812 43376 20864 43382
rect 21100 43330 21128 44662
rect 21192 44402 21220 45290
rect 21180 44396 21232 44402
rect 21180 44338 21232 44344
rect 21180 43852 21232 43858
rect 21180 43794 21232 43800
rect 20812 43318 20864 43324
rect 20720 43308 20772 43314
rect 20720 43250 20772 43256
rect 21008 43302 21128 43330
rect 20732 42906 20760 43250
rect 20720 42900 20772 42906
rect 20720 42842 20772 42848
rect 20536 42356 20588 42362
rect 20588 42316 20668 42344
rect 20536 42298 20588 42304
rect 20536 41676 20588 41682
rect 20536 41618 20588 41624
rect 20352 41608 20404 41614
rect 20352 41550 20404 41556
rect 20364 41274 20392 41550
rect 20352 41268 20404 41274
rect 20352 41210 20404 41216
rect 20442 41168 20498 41177
rect 20442 41103 20444 41112
rect 20496 41103 20498 41112
rect 20444 41074 20496 41080
rect 20548 40526 20576 41618
rect 20536 40520 20588 40526
rect 20536 40462 20588 40468
rect 20640 40202 20668 42316
rect 21008 42294 21036 43302
rect 21192 42362 21220 43794
rect 21284 43722 21312 45444
rect 21272 43716 21324 43722
rect 21272 43658 21324 43664
rect 21180 42356 21232 42362
rect 21180 42298 21232 42304
rect 20996 42288 21048 42294
rect 20996 42230 21048 42236
rect 20904 42220 20956 42226
rect 20904 42162 20956 42168
rect 21180 42220 21232 42226
rect 21284 42208 21312 43658
rect 21468 43654 21496 45766
rect 21652 45558 21680 46582
rect 21744 45937 21772 46990
rect 22020 46934 22048 47466
rect 23216 47258 23244 49200
rect 23204 47252 23256 47258
rect 23204 47194 23256 47200
rect 22192 47048 22244 47054
rect 22192 46990 22244 46996
rect 24400 47048 24452 47054
rect 24400 46990 24452 46996
rect 24584 47048 24636 47054
rect 24584 46990 24636 46996
rect 24952 47048 25004 47054
rect 24952 46990 25004 46996
rect 22020 46906 22140 46934
rect 22112 46646 22140 46906
rect 22100 46640 22152 46646
rect 22100 46582 22152 46588
rect 21824 46572 21876 46578
rect 21824 46514 21876 46520
rect 21730 45928 21786 45937
rect 21730 45863 21786 45872
rect 21744 45626 21772 45863
rect 21732 45620 21784 45626
rect 21732 45562 21784 45568
rect 21640 45552 21692 45558
rect 21640 45494 21692 45500
rect 21836 45422 21864 46514
rect 22204 46442 22232 46990
rect 22284 46980 22336 46986
rect 22284 46922 22336 46928
rect 22192 46436 22244 46442
rect 22192 46378 22244 46384
rect 22204 46034 22232 46378
rect 22008 46028 22060 46034
rect 22008 45970 22060 45976
rect 22192 46028 22244 46034
rect 22192 45970 22244 45976
rect 21916 45960 21968 45966
rect 21916 45902 21968 45908
rect 21824 45416 21876 45422
rect 21824 45358 21876 45364
rect 21640 45076 21692 45082
rect 21640 45018 21692 45024
rect 21652 44946 21680 45018
rect 21640 44940 21692 44946
rect 21640 44882 21692 44888
rect 21652 44198 21680 44882
rect 21732 44872 21784 44878
rect 21732 44814 21784 44820
rect 21744 44538 21772 44814
rect 21732 44532 21784 44538
rect 21732 44474 21784 44480
rect 21824 44396 21876 44402
rect 21928 44384 21956 45902
rect 22020 45422 22048 45970
rect 22100 45960 22152 45966
rect 22100 45902 22152 45908
rect 22112 45626 22140 45902
rect 22192 45824 22244 45830
rect 22192 45766 22244 45772
rect 22100 45620 22152 45626
rect 22100 45562 22152 45568
rect 22008 45416 22060 45422
rect 22008 45358 22060 45364
rect 22020 44946 22048 45358
rect 22112 45082 22140 45562
rect 22204 45558 22232 45766
rect 22192 45552 22244 45558
rect 22192 45494 22244 45500
rect 22296 45490 22324 46922
rect 24412 46714 24440 46990
rect 24400 46708 24452 46714
rect 24400 46650 24452 46656
rect 24400 46572 24452 46578
rect 24400 46514 24452 46520
rect 22928 46504 22980 46510
rect 22928 46446 22980 46452
rect 23572 46504 23624 46510
rect 23572 46446 23624 46452
rect 22940 45558 22968 46446
rect 23388 46164 23440 46170
rect 23388 46106 23440 46112
rect 22928 45552 22980 45558
rect 23204 45552 23256 45558
rect 22928 45494 22980 45500
rect 23124 45512 23204 45540
rect 22284 45484 22336 45490
rect 22284 45426 22336 45432
rect 22100 45076 22152 45082
rect 22100 45018 22152 45024
rect 22192 45008 22244 45014
rect 22192 44950 22244 44956
rect 22008 44940 22060 44946
rect 22008 44882 22060 44888
rect 22008 44736 22060 44742
rect 22008 44678 22060 44684
rect 22020 44402 22048 44678
rect 21876 44356 21956 44384
rect 22008 44396 22060 44402
rect 21824 44338 21876 44344
rect 22008 44338 22060 44344
rect 21640 44192 21692 44198
rect 21640 44134 21692 44140
rect 22008 43852 22060 43858
rect 22008 43794 22060 43800
rect 21548 43784 21600 43790
rect 21548 43726 21600 43732
rect 21456 43648 21508 43654
rect 21456 43590 21508 43596
rect 21468 42226 21496 43590
rect 21560 43450 21588 43726
rect 21548 43444 21600 43450
rect 21548 43386 21600 43392
rect 22020 43314 22048 43794
rect 22204 43722 22232 44950
rect 22296 44878 22324 45426
rect 22284 44872 22336 44878
rect 22284 44814 22336 44820
rect 22284 44532 22336 44538
rect 22284 44474 22336 44480
rect 22296 44334 22324 44474
rect 23124 44334 23152 45512
rect 23204 45494 23256 45500
rect 23204 45280 23256 45286
rect 23204 45222 23256 45228
rect 23216 44810 23244 45222
rect 23204 44804 23256 44810
rect 23204 44746 23256 44752
rect 22284 44328 22336 44334
rect 22284 44270 22336 44276
rect 23112 44328 23164 44334
rect 23112 44270 23164 44276
rect 22296 43790 22324 44270
rect 22928 44192 22980 44198
rect 22928 44134 22980 44140
rect 22284 43784 22336 43790
rect 22284 43726 22336 43732
rect 22744 43784 22796 43790
rect 22744 43726 22796 43732
rect 22192 43716 22244 43722
rect 22192 43658 22244 43664
rect 22100 43648 22152 43654
rect 22100 43590 22152 43596
rect 22468 43648 22520 43654
rect 22468 43590 22520 43596
rect 22008 43308 22060 43314
rect 22008 43250 22060 43256
rect 21916 43104 21968 43110
rect 21916 43046 21968 43052
rect 21640 42900 21692 42906
rect 21640 42842 21692 42848
rect 21548 42696 21600 42702
rect 21548 42638 21600 42644
rect 21560 42226 21588 42638
rect 21456 42220 21508 42226
rect 21232 42180 21312 42208
rect 21376 42180 21456 42208
rect 21180 42162 21232 42168
rect 20720 42016 20772 42022
rect 20720 41958 20772 41964
rect 20732 41818 20760 41958
rect 20720 41812 20772 41818
rect 20720 41754 20772 41760
rect 20260 40180 20312 40186
rect 20260 40122 20312 40128
rect 20456 40174 20668 40202
rect 20076 40112 20128 40118
rect 20076 40054 20128 40060
rect 19984 39976 20036 39982
rect 18880 39918 18932 39924
rect 19430 39944 19486 39953
rect 18328 39908 18380 39914
rect 19984 39918 20036 39924
rect 19430 39879 19486 39888
rect 18328 39850 18380 39856
rect 18420 39840 18472 39846
rect 18420 39782 18472 39788
rect 19432 39840 19484 39846
rect 19432 39782 19484 39788
rect 18328 39500 18380 39506
rect 18328 39442 18380 39448
rect 18064 38814 18276 38842
rect 17960 38208 18012 38214
rect 17960 38150 18012 38156
rect 17868 37868 17920 37874
rect 17788 37828 17868 37856
rect 17684 37800 17736 37806
rect 17684 37742 17736 37748
rect 17500 37256 17552 37262
rect 17500 37198 17552 37204
rect 17512 36174 17540 37198
rect 17696 36174 17724 37742
rect 17788 37126 17816 37828
rect 17868 37810 17920 37816
rect 18064 37466 18092 38814
rect 18340 38758 18368 39442
rect 18328 38752 18380 38758
rect 18328 38694 18380 38700
rect 18144 38412 18196 38418
rect 18144 38354 18196 38360
rect 18236 38412 18288 38418
rect 18236 38354 18288 38360
rect 18156 38282 18184 38354
rect 18144 38276 18196 38282
rect 18144 38218 18196 38224
rect 18144 38004 18196 38010
rect 18144 37946 18196 37952
rect 18156 37738 18184 37946
rect 18248 37738 18276 38354
rect 18144 37732 18196 37738
rect 18144 37674 18196 37680
rect 18236 37732 18288 37738
rect 18236 37674 18288 37680
rect 18052 37460 18104 37466
rect 18052 37402 18104 37408
rect 17776 37120 17828 37126
rect 17776 37062 17828 37068
rect 17788 36242 17816 37062
rect 17960 36848 18012 36854
rect 17960 36790 18012 36796
rect 17776 36236 17828 36242
rect 17776 36178 17828 36184
rect 17500 36168 17552 36174
rect 17500 36110 17552 36116
rect 17684 36168 17736 36174
rect 17684 36110 17736 36116
rect 17512 35834 17540 36110
rect 17972 36038 18000 36790
rect 17960 36032 18012 36038
rect 17960 35974 18012 35980
rect 18064 35850 18092 37402
rect 18236 36372 18288 36378
rect 18236 36314 18288 36320
rect 17500 35828 17552 35834
rect 17500 35770 17552 35776
rect 17972 35822 18092 35850
rect 17500 35624 17552 35630
rect 17500 35566 17552 35572
rect 17316 34468 17368 34474
rect 17316 34410 17368 34416
rect 17512 32910 17540 35566
rect 17972 35562 18000 35822
rect 18248 35766 18276 36314
rect 18340 36258 18368 38694
rect 18432 37330 18460 39782
rect 18880 39432 18932 39438
rect 18880 39374 18932 39380
rect 18892 39030 18920 39374
rect 19444 39302 19472 39782
rect 19340 39296 19392 39302
rect 19340 39238 19392 39244
rect 19432 39296 19484 39302
rect 19432 39238 19484 39244
rect 19352 39030 19380 39238
rect 19444 39098 19472 39238
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19432 39092 19484 39098
rect 19432 39034 19484 39040
rect 18880 39024 18932 39030
rect 18880 38966 18932 38972
rect 19340 39024 19392 39030
rect 19340 38966 19392 38972
rect 18604 38956 18656 38962
rect 18604 38898 18656 38904
rect 18616 38486 18644 38898
rect 18604 38480 18656 38486
rect 18604 38422 18656 38428
rect 18512 38344 18564 38350
rect 18510 38312 18512 38321
rect 18564 38312 18566 38321
rect 18510 38247 18566 38256
rect 18696 37800 18748 37806
rect 18694 37768 18696 37777
rect 18748 37768 18750 37777
rect 18616 37726 18694 37754
rect 18420 37324 18472 37330
rect 18420 37266 18472 37272
rect 18512 37256 18564 37262
rect 18512 37198 18564 37204
rect 18524 36786 18552 37198
rect 18616 36786 18644 37726
rect 18892 37754 18920 38966
rect 19248 38888 19300 38894
rect 19248 38830 19300 38836
rect 19156 38752 19208 38758
rect 19156 38694 19208 38700
rect 19168 38486 19196 38694
rect 19260 38554 19288 38830
rect 19352 38826 19380 38966
rect 20076 38956 20128 38962
rect 20076 38898 20128 38904
rect 19340 38820 19392 38826
rect 19340 38762 19392 38768
rect 19248 38548 19300 38554
rect 19248 38490 19300 38496
rect 19156 38480 19208 38486
rect 19156 38422 19208 38428
rect 18972 38276 19024 38282
rect 18972 38218 19024 38224
rect 18984 37874 19012 38218
rect 18972 37868 19024 37874
rect 18972 37810 19024 37816
rect 18892 37726 19104 37754
rect 18694 37703 18750 37712
rect 19076 37398 19104 37726
rect 19352 37482 19380 38762
rect 19616 38752 19668 38758
rect 19616 38694 19668 38700
rect 19628 38321 19656 38694
rect 19892 38344 19944 38350
rect 19614 38312 19670 38321
rect 19944 38304 20024 38332
rect 19892 38286 19944 38292
rect 19614 38247 19670 38256
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19892 37664 19944 37670
rect 19890 37632 19892 37641
rect 19944 37632 19946 37641
rect 19890 37567 19946 37576
rect 19156 37460 19208 37466
rect 19352 37454 19472 37482
rect 19156 37402 19208 37408
rect 19064 37392 19116 37398
rect 19064 37334 19116 37340
rect 18880 37188 18932 37194
rect 18880 37130 18932 37136
rect 18696 36848 18748 36854
rect 18696 36790 18748 36796
rect 18512 36780 18564 36786
rect 18512 36722 18564 36728
rect 18604 36780 18656 36786
rect 18604 36722 18656 36728
rect 18524 36378 18552 36722
rect 18708 36718 18736 36790
rect 18892 36786 18920 37130
rect 18880 36780 18932 36786
rect 18880 36722 18932 36728
rect 18696 36712 18748 36718
rect 18602 36680 18658 36689
rect 18696 36654 18748 36660
rect 18602 36615 18658 36624
rect 18512 36372 18564 36378
rect 18512 36314 18564 36320
rect 18340 36230 18460 36258
rect 18328 36100 18380 36106
rect 18328 36042 18380 36048
rect 18236 35760 18288 35766
rect 18236 35702 18288 35708
rect 17960 35556 18012 35562
rect 17960 35498 18012 35504
rect 17972 34678 18000 35498
rect 18248 35290 18276 35702
rect 18340 35494 18368 36042
rect 18432 35630 18460 36230
rect 18512 36032 18564 36038
rect 18512 35974 18564 35980
rect 18524 35698 18552 35974
rect 18512 35692 18564 35698
rect 18512 35634 18564 35640
rect 18420 35624 18472 35630
rect 18420 35566 18472 35572
rect 18328 35488 18380 35494
rect 18328 35430 18380 35436
rect 18340 35290 18368 35430
rect 18236 35284 18288 35290
rect 18236 35226 18288 35232
rect 18328 35284 18380 35290
rect 18328 35226 18380 35232
rect 18524 35086 18552 35634
rect 18144 35080 18196 35086
rect 18144 35022 18196 35028
rect 18512 35080 18564 35086
rect 18512 35022 18564 35028
rect 18052 34944 18104 34950
rect 18052 34886 18104 34892
rect 17960 34672 18012 34678
rect 17960 34614 18012 34620
rect 17960 34400 18012 34406
rect 17960 34342 18012 34348
rect 17972 34202 18000 34342
rect 17960 34196 18012 34202
rect 17960 34138 18012 34144
rect 18064 33522 18092 34886
rect 18156 33658 18184 35022
rect 18420 33992 18472 33998
rect 18420 33934 18472 33940
rect 18144 33652 18196 33658
rect 18144 33594 18196 33600
rect 18156 33522 18184 33594
rect 18052 33516 18104 33522
rect 18052 33458 18104 33464
rect 18144 33516 18196 33522
rect 18144 33458 18196 33464
rect 18328 33516 18380 33522
rect 18328 33458 18380 33464
rect 18064 33402 18092 33458
rect 18064 33374 18276 33402
rect 18144 33312 18196 33318
rect 18144 33254 18196 33260
rect 17868 33108 17920 33114
rect 17868 33050 17920 33056
rect 17316 32904 17368 32910
rect 17316 32846 17368 32852
rect 17500 32904 17552 32910
rect 17500 32846 17552 32852
rect 17328 32434 17356 32846
rect 17408 32564 17460 32570
rect 17408 32506 17460 32512
rect 17316 32428 17368 32434
rect 17316 32370 17368 32376
rect 17420 31822 17448 32506
rect 17512 32366 17540 32846
rect 17880 32502 17908 33050
rect 18156 32910 18184 33254
rect 17960 32904 18012 32910
rect 17960 32846 18012 32852
rect 18144 32904 18196 32910
rect 18144 32846 18196 32852
rect 17868 32496 17920 32502
rect 17868 32438 17920 32444
rect 17500 32360 17552 32366
rect 17500 32302 17552 32308
rect 17972 32298 18000 32846
rect 18052 32768 18104 32774
rect 18052 32710 18104 32716
rect 17960 32292 18012 32298
rect 17960 32234 18012 32240
rect 17592 32224 17644 32230
rect 17592 32166 17644 32172
rect 17408 31816 17460 31822
rect 17408 31758 17460 31764
rect 17500 31748 17552 31754
rect 17500 31690 17552 31696
rect 17408 31680 17460 31686
rect 17408 31622 17460 31628
rect 17316 31340 17368 31346
rect 17316 31282 17368 31288
rect 17328 30870 17356 31282
rect 17420 30938 17448 31622
rect 17512 31346 17540 31690
rect 17604 31686 17632 32166
rect 17868 31816 17920 31822
rect 17868 31758 17920 31764
rect 17592 31680 17644 31686
rect 17592 31622 17644 31628
rect 17880 31482 17908 31758
rect 17972 31686 18000 32234
rect 17960 31680 18012 31686
rect 17960 31622 18012 31628
rect 17868 31476 17920 31482
rect 17868 31418 17920 31424
rect 18064 31346 18092 32710
rect 18156 31804 18184 32846
rect 18248 32366 18276 33374
rect 18340 32434 18368 33458
rect 18432 33454 18460 33934
rect 18512 33856 18564 33862
rect 18512 33798 18564 33804
rect 18524 33522 18552 33798
rect 18512 33516 18564 33522
rect 18512 33458 18564 33464
rect 18420 33448 18472 33454
rect 18616 33402 18644 36615
rect 18708 36106 18736 36654
rect 18696 36100 18748 36106
rect 18696 36042 18748 36048
rect 18786 35728 18842 35737
rect 19076 35698 19104 37334
rect 19168 36038 19196 37402
rect 19248 37324 19300 37330
rect 19300 37284 19380 37312
rect 19248 37266 19300 37272
rect 19352 36786 19380 37284
rect 19340 36780 19392 36786
rect 19340 36722 19392 36728
rect 19340 36644 19392 36650
rect 19340 36586 19392 36592
rect 19352 36378 19380 36586
rect 19340 36372 19392 36378
rect 19340 36314 19392 36320
rect 19444 36174 19472 37454
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19706 36816 19762 36825
rect 19706 36751 19708 36760
rect 19760 36751 19762 36760
rect 19892 36780 19944 36786
rect 19708 36722 19760 36728
rect 19996 36768 20024 38304
rect 19944 36740 20024 36768
rect 19892 36722 19944 36728
rect 19720 36650 19748 36722
rect 19904 36689 19932 36722
rect 19890 36680 19946 36689
rect 19708 36644 19760 36650
rect 19890 36615 19946 36624
rect 19708 36586 19760 36592
rect 20088 36582 20116 38898
rect 20272 38654 20300 40122
rect 20352 40044 20404 40050
rect 20352 39986 20404 39992
rect 20364 39506 20392 39986
rect 20456 39846 20484 40174
rect 20536 40112 20588 40118
rect 20536 40054 20588 40060
rect 20718 40080 20774 40089
rect 20444 39840 20496 39846
rect 20444 39782 20496 39788
rect 20352 39500 20404 39506
rect 20352 39442 20404 39448
rect 20180 38626 20300 38654
rect 20180 38350 20208 38626
rect 20364 38554 20392 39442
rect 20548 39370 20576 40054
rect 20718 40015 20774 40024
rect 20628 39976 20680 39982
rect 20628 39918 20680 39924
rect 20640 39438 20668 39918
rect 20628 39432 20680 39438
rect 20628 39374 20680 39380
rect 20536 39364 20588 39370
rect 20536 39306 20588 39312
rect 20548 38554 20576 39306
rect 20640 39030 20668 39374
rect 20732 39302 20760 40015
rect 20812 39840 20864 39846
rect 20812 39782 20864 39788
rect 20824 39370 20852 39782
rect 20812 39364 20864 39370
rect 20812 39306 20864 39312
rect 20720 39296 20772 39302
rect 20720 39238 20772 39244
rect 20628 39024 20680 39030
rect 20628 38966 20680 38972
rect 20812 38956 20864 38962
rect 20812 38898 20864 38904
rect 20824 38826 20852 38898
rect 20812 38820 20864 38826
rect 20812 38762 20864 38768
rect 20352 38548 20404 38554
rect 20352 38490 20404 38496
rect 20536 38548 20588 38554
rect 20536 38490 20588 38496
rect 20168 38344 20220 38350
rect 20168 38286 20220 38292
rect 20180 37346 20208 38286
rect 20364 37874 20392 38490
rect 20444 38344 20496 38350
rect 20444 38286 20496 38292
rect 20352 37868 20404 37874
rect 20352 37810 20404 37816
rect 20180 37318 20300 37346
rect 20364 37330 20392 37810
rect 20168 37120 20220 37126
rect 20166 37088 20168 37097
rect 20220 37088 20222 37097
rect 20166 37023 20222 37032
rect 20272 36650 20300 37318
rect 20352 37324 20404 37330
rect 20352 37266 20404 37272
rect 20456 37240 20484 38286
rect 20548 37466 20576 38490
rect 20720 38344 20772 38350
rect 20720 38286 20772 38292
rect 20628 37664 20680 37670
rect 20628 37606 20680 37612
rect 20536 37460 20588 37466
rect 20536 37402 20588 37408
rect 20444 37234 20496 37240
rect 20444 37176 20496 37182
rect 20536 37234 20588 37240
rect 20536 37176 20588 37182
rect 20260 36644 20312 36650
rect 20260 36586 20312 36592
rect 20076 36576 20128 36582
rect 20076 36518 20128 36524
rect 19984 36236 20036 36242
rect 19984 36178 20036 36184
rect 19432 36168 19484 36174
rect 19432 36110 19484 36116
rect 19156 36032 19208 36038
rect 19156 35974 19208 35980
rect 19444 35698 19472 36110
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19800 35828 19852 35834
rect 19996 35816 20024 36178
rect 19800 35770 19852 35776
rect 19904 35788 20024 35816
rect 18786 35663 18842 35672
rect 18972 35692 19024 35698
rect 18800 34950 18828 35663
rect 18972 35634 19024 35640
rect 19064 35692 19116 35698
rect 19064 35634 19116 35640
rect 19432 35692 19484 35698
rect 19432 35634 19484 35640
rect 18880 35624 18932 35630
rect 18880 35566 18932 35572
rect 18892 35290 18920 35566
rect 18880 35284 18932 35290
rect 18880 35226 18932 35232
rect 18788 34944 18840 34950
rect 18788 34886 18840 34892
rect 18800 34678 18828 34886
rect 18788 34672 18840 34678
rect 18788 34614 18840 34620
rect 18696 33924 18748 33930
rect 18696 33866 18748 33872
rect 18708 33590 18736 33866
rect 18984 33862 19012 35634
rect 19076 34134 19104 35634
rect 19444 35290 19472 35634
rect 19432 35284 19484 35290
rect 19432 35226 19484 35232
rect 19444 35018 19472 35226
rect 19812 35086 19840 35770
rect 19904 35698 19932 35788
rect 19892 35692 19944 35698
rect 19892 35634 19944 35640
rect 19984 35692 20036 35698
rect 19984 35634 20036 35640
rect 19904 35290 19932 35634
rect 19892 35284 19944 35290
rect 19892 35226 19944 35232
rect 19996 35154 20024 35634
rect 19984 35148 20036 35154
rect 19984 35090 20036 35096
rect 19800 35080 19852 35086
rect 19800 35022 19852 35028
rect 19432 35012 19484 35018
rect 19432 34954 19484 34960
rect 19340 34944 19392 34950
rect 19340 34886 19392 34892
rect 19352 34746 19380 34886
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19996 34746 20024 35090
rect 20076 35012 20128 35018
rect 20076 34954 20128 34960
rect 19340 34740 19392 34746
rect 19340 34682 19392 34688
rect 19984 34740 20036 34746
rect 19984 34682 20036 34688
rect 19248 34604 19300 34610
rect 19248 34546 19300 34552
rect 19340 34604 19392 34610
rect 19340 34546 19392 34552
rect 19064 34128 19116 34134
rect 19064 34070 19116 34076
rect 19260 34066 19288 34546
rect 19248 34060 19300 34066
rect 19248 34002 19300 34008
rect 18972 33856 19024 33862
rect 18972 33798 19024 33804
rect 19260 33658 19288 34002
rect 19352 33998 19380 34546
rect 19432 34536 19484 34542
rect 19432 34478 19484 34484
rect 19340 33992 19392 33998
rect 19340 33934 19392 33940
rect 19248 33652 19300 33658
rect 19248 33594 19300 33600
rect 18696 33584 18748 33590
rect 18696 33526 18748 33532
rect 18708 33454 18736 33526
rect 19260 33454 19288 33594
rect 18420 33390 18472 33396
rect 18432 33289 18460 33390
rect 18524 33374 18644 33402
rect 18696 33448 18748 33454
rect 18696 33390 18748 33396
rect 19248 33448 19300 33454
rect 19248 33390 19300 33396
rect 18880 33380 18932 33386
rect 18418 33280 18474 33289
rect 18418 33215 18474 33224
rect 18328 32428 18380 32434
rect 18328 32370 18380 32376
rect 18236 32360 18288 32366
rect 18236 32302 18288 32308
rect 18328 31816 18380 31822
rect 18156 31776 18328 31804
rect 18328 31758 18380 31764
rect 18524 31754 18552 33374
rect 18880 33322 18932 33328
rect 18892 33046 18920 33322
rect 18880 33040 18932 33046
rect 18880 32982 18932 32988
rect 18788 32768 18840 32774
rect 18788 32710 18840 32716
rect 18800 32416 18828 32710
rect 18708 32388 18828 32416
rect 18524 31726 18644 31754
rect 17500 31340 17552 31346
rect 17500 31282 17552 31288
rect 18052 31340 18104 31346
rect 18052 31282 18104 31288
rect 17408 30932 17460 30938
rect 17408 30874 17460 30880
rect 17316 30864 17368 30870
rect 17316 30806 17368 30812
rect 17328 30666 17356 30806
rect 17512 30802 17540 31282
rect 17500 30796 17552 30802
rect 17500 30738 17552 30744
rect 18064 30734 18092 31282
rect 18052 30728 18104 30734
rect 18052 30670 18104 30676
rect 17316 30660 17368 30666
rect 17316 30602 17368 30608
rect 17328 30394 17356 30602
rect 18064 30394 18092 30670
rect 17316 30388 17368 30394
rect 17316 30330 17368 30336
rect 18052 30388 18104 30394
rect 18052 30330 18104 30336
rect 17776 30048 17828 30054
rect 17776 29990 17828 29996
rect 17960 30048 18012 30054
rect 17960 29990 18012 29996
rect 17788 29850 17816 29990
rect 17776 29844 17828 29850
rect 17776 29786 17828 29792
rect 17684 29572 17736 29578
rect 17684 29514 17736 29520
rect 17696 29306 17724 29514
rect 17684 29300 17736 29306
rect 17684 29242 17736 29248
rect 17224 29164 17276 29170
rect 17224 29106 17276 29112
rect 17592 29164 17644 29170
rect 17592 29106 17644 29112
rect 16948 29028 17000 29034
rect 16948 28970 17000 28976
rect 17604 28558 17632 29106
rect 17696 28558 17724 29242
rect 17972 29170 18000 29990
rect 18616 29646 18644 31726
rect 18708 30938 18736 32388
rect 18892 31958 18920 32982
rect 19352 32978 19380 33934
rect 19340 32972 19392 32978
rect 19340 32914 19392 32920
rect 19352 32434 19380 32914
rect 19444 32570 19472 34478
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 20088 33674 20116 34954
rect 19996 33646 20116 33674
rect 19996 32910 20024 33646
rect 20076 33584 20128 33590
rect 20076 33526 20128 33532
rect 19984 32904 20036 32910
rect 19984 32846 20036 32852
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19432 32564 19484 32570
rect 19432 32506 19484 32512
rect 19340 32428 19392 32434
rect 19340 32370 19392 32376
rect 19352 32026 19380 32370
rect 19340 32020 19392 32026
rect 19340 31962 19392 31968
rect 18880 31952 18932 31958
rect 18880 31894 18932 31900
rect 19444 31822 19472 32506
rect 19996 32434 20024 32846
rect 19984 32428 20036 32434
rect 19984 32370 20036 32376
rect 18788 31816 18840 31822
rect 19432 31816 19484 31822
rect 18788 31758 18840 31764
rect 19352 31776 19432 31804
rect 18696 30932 18748 30938
rect 18696 30874 18748 30880
rect 18604 29640 18656 29646
rect 18604 29582 18656 29588
rect 18420 29504 18472 29510
rect 18420 29446 18472 29452
rect 18432 29238 18460 29446
rect 18420 29232 18472 29238
rect 18420 29174 18472 29180
rect 17960 29164 18012 29170
rect 17960 29106 18012 29112
rect 17776 29028 17828 29034
rect 17776 28970 17828 28976
rect 17788 28694 17816 28970
rect 17776 28688 17828 28694
rect 17776 28630 17828 28636
rect 17972 28558 18000 29106
rect 18236 29096 18288 29102
rect 18236 29038 18288 29044
rect 16672 28552 16724 28558
rect 16672 28494 16724 28500
rect 17592 28552 17644 28558
rect 17592 28494 17644 28500
rect 17684 28552 17736 28558
rect 17684 28494 17736 28500
rect 17960 28552 18012 28558
rect 17960 28494 18012 28500
rect 15752 28416 15804 28422
rect 15752 28358 15804 28364
rect 16120 28416 16172 28422
rect 16120 28358 16172 28364
rect 17960 28416 18012 28422
rect 17960 28358 18012 28364
rect 15764 21894 15792 28358
rect 17972 27946 18000 28358
rect 18248 28082 18276 29038
rect 18328 28756 18380 28762
rect 18328 28698 18380 28704
rect 18340 28150 18368 28698
rect 18432 28218 18460 29174
rect 18420 28212 18472 28218
rect 18420 28154 18472 28160
rect 18328 28144 18380 28150
rect 18328 28086 18380 28092
rect 18236 28076 18288 28082
rect 18236 28018 18288 28024
rect 17960 27940 18012 27946
rect 17960 27882 18012 27888
rect 18616 27878 18644 29582
rect 18800 29170 18828 31758
rect 19352 31754 19380 31776
rect 19432 31758 19484 31764
rect 19260 31726 19380 31754
rect 19260 31414 19288 31726
rect 19338 31648 19394 31657
rect 19338 31583 19394 31592
rect 19248 31408 19300 31414
rect 19248 31350 19300 31356
rect 18972 31340 19024 31346
rect 18972 31282 19024 31288
rect 18984 29850 19012 31282
rect 19352 30274 19380 31583
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19996 31482 20024 32370
rect 19984 31476 20036 31482
rect 19984 31418 20036 31424
rect 19892 31340 19944 31346
rect 19892 31282 19944 31288
rect 19800 31136 19852 31142
rect 19800 31078 19852 31084
rect 19812 30870 19840 31078
rect 19800 30864 19852 30870
rect 19800 30806 19852 30812
rect 19432 30728 19484 30734
rect 19432 30670 19484 30676
rect 19444 30394 19472 30670
rect 19904 30648 19932 31282
rect 20088 31210 20116 33526
rect 20168 33448 20220 33454
rect 20168 33390 20220 33396
rect 20180 33114 20208 33390
rect 20168 33108 20220 33114
rect 20168 33050 20220 33056
rect 20166 31784 20222 31793
rect 20272 31770 20300 36586
rect 20456 36378 20484 37176
rect 20548 36922 20576 37176
rect 20640 37126 20668 37606
rect 20628 37120 20680 37126
rect 20628 37062 20680 37068
rect 20536 36916 20588 36922
rect 20536 36858 20588 36864
rect 20640 36854 20668 37062
rect 20732 36922 20760 38286
rect 20824 37670 20852 38762
rect 20812 37664 20864 37670
rect 20812 37606 20864 37612
rect 20824 37398 20852 37606
rect 20812 37392 20864 37398
rect 20812 37334 20864 37340
rect 20720 36916 20772 36922
rect 20720 36858 20772 36864
rect 20628 36848 20680 36854
rect 20628 36790 20680 36796
rect 20536 36780 20588 36786
rect 20536 36722 20588 36728
rect 20548 36650 20576 36722
rect 20628 36712 20680 36718
rect 20628 36654 20680 36660
rect 20536 36644 20588 36650
rect 20536 36586 20588 36592
rect 20548 36553 20576 36586
rect 20534 36544 20590 36553
rect 20534 36479 20590 36488
rect 20444 36372 20496 36378
rect 20444 36314 20496 36320
rect 20548 36258 20576 36479
rect 20456 36230 20576 36258
rect 20456 36174 20484 36230
rect 20640 36174 20668 36654
rect 20444 36168 20496 36174
rect 20444 36110 20496 36116
rect 20628 36168 20680 36174
rect 20628 36110 20680 36116
rect 20456 36009 20484 36110
rect 20442 36000 20498 36009
rect 20442 35935 20498 35944
rect 20812 35692 20864 35698
rect 20812 35634 20864 35640
rect 20824 35290 20852 35634
rect 20812 35284 20864 35290
rect 20812 35226 20864 35232
rect 20720 35080 20772 35086
rect 20720 35022 20772 35028
rect 20732 34542 20760 35022
rect 20720 34536 20772 34542
rect 20720 34478 20772 34484
rect 20444 34060 20496 34066
rect 20444 34002 20496 34008
rect 20456 32910 20484 34002
rect 20536 33856 20588 33862
rect 20536 33798 20588 33804
rect 20548 33522 20576 33798
rect 20536 33516 20588 33522
rect 20536 33458 20588 33464
rect 20732 33114 20760 34478
rect 20720 33108 20772 33114
rect 20720 33050 20772 33056
rect 20444 32904 20496 32910
rect 20444 32846 20496 32852
rect 20456 32298 20484 32846
rect 20444 32292 20496 32298
rect 20444 32234 20496 32240
rect 20222 31742 20300 31770
rect 20166 31719 20222 31728
rect 20076 31204 20128 31210
rect 20076 31146 20128 31152
rect 19984 31136 20036 31142
rect 19984 31078 20036 31084
rect 19996 30938 20024 31078
rect 19984 30932 20036 30938
rect 19984 30874 20036 30880
rect 20076 30932 20128 30938
rect 20076 30874 20128 30880
rect 19904 30620 20024 30648
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19432 30388 19484 30394
rect 19432 30330 19484 30336
rect 19260 30258 19380 30274
rect 19248 30252 19380 30258
rect 19300 30246 19380 30252
rect 19524 30252 19576 30258
rect 19248 30194 19300 30200
rect 19524 30194 19576 30200
rect 18972 29844 19024 29850
rect 18972 29786 19024 29792
rect 19156 29572 19208 29578
rect 19156 29514 19208 29520
rect 18880 29300 18932 29306
rect 18880 29242 18932 29248
rect 18788 29164 18840 29170
rect 18788 29106 18840 29112
rect 18800 28150 18828 29106
rect 18892 28762 18920 29242
rect 19168 29170 19196 29514
rect 19064 29164 19116 29170
rect 19064 29106 19116 29112
rect 19156 29164 19208 29170
rect 19156 29106 19208 29112
rect 19076 28762 19104 29106
rect 18880 28756 18932 28762
rect 18880 28698 18932 28704
rect 19064 28756 19116 28762
rect 19064 28698 19116 28704
rect 18788 28144 18840 28150
rect 18788 28086 18840 28092
rect 19260 27946 19288 30194
rect 19340 30184 19392 30190
rect 19340 30126 19392 30132
rect 19352 29782 19380 30126
rect 19432 30116 19484 30122
rect 19432 30058 19484 30064
rect 19340 29776 19392 29782
rect 19340 29718 19392 29724
rect 19352 29646 19380 29718
rect 19340 29640 19392 29646
rect 19340 29582 19392 29588
rect 19352 29306 19380 29582
rect 19444 29510 19472 30058
rect 19536 29646 19564 30194
rect 19524 29640 19576 29646
rect 19524 29582 19576 29588
rect 19432 29504 19484 29510
rect 19432 29446 19484 29452
rect 19340 29300 19392 29306
rect 19340 29242 19392 29248
rect 19444 29186 19472 29446
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19352 29158 19472 29186
rect 19524 29164 19576 29170
rect 19352 28558 19380 29158
rect 19800 29164 19852 29170
rect 19576 29124 19800 29152
rect 19524 29106 19576 29112
rect 19800 29106 19852 29112
rect 19996 28966 20024 30620
rect 20088 30598 20116 30874
rect 20076 30592 20128 30598
rect 20076 30534 20128 30540
rect 20088 30190 20116 30534
rect 20076 30184 20128 30190
rect 20076 30126 20128 30132
rect 20088 29850 20116 30126
rect 20076 29844 20128 29850
rect 20076 29786 20128 29792
rect 20180 29646 20208 31719
rect 20456 31142 20484 32234
rect 20720 32224 20772 32230
rect 20720 32166 20772 32172
rect 20812 32224 20864 32230
rect 20812 32166 20864 32172
rect 20732 31890 20760 32166
rect 20824 31958 20852 32166
rect 20812 31952 20864 31958
rect 20812 31894 20864 31900
rect 20720 31884 20772 31890
rect 20720 31826 20772 31832
rect 20444 31136 20496 31142
rect 20444 31078 20496 31084
rect 20444 30864 20496 30870
rect 20444 30806 20496 30812
rect 20536 30864 20588 30870
rect 20536 30806 20588 30812
rect 20352 30660 20404 30666
rect 20352 30602 20404 30608
rect 20076 29640 20128 29646
rect 20076 29582 20128 29588
rect 20168 29640 20220 29646
rect 20168 29582 20220 29588
rect 20088 29102 20116 29582
rect 20260 29504 20312 29510
rect 20260 29446 20312 29452
rect 20076 29096 20128 29102
rect 20076 29038 20128 29044
rect 19984 28960 20036 28966
rect 19984 28902 20036 28908
rect 19340 28552 19392 28558
rect 19340 28494 19392 28500
rect 19248 27940 19300 27946
rect 19248 27882 19300 27888
rect 19352 27878 19380 28494
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19708 28076 19760 28082
rect 19708 28018 19760 28024
rect 19892 28076 19944 28082
rect 19892 28018 19944 28024
rect 19432 27940 19484 27946
rect 19432 27882 19484 27888
rect 18604 27872 18656 27878
rect 18604 27814 18656 27820
rect 19340 27872 19392 27878
rect 19340 27814 19392 27820
rect 18616 27606 18644 27814
rect 19444 27674 19472 27882
rect 19432 27668 19484 27674
rect 19432 27610 19484 27616
rect 18604 27600 18656 27606
rect 18604 27542 18656 27548
rect 18616 27130 18644 27542
rect 19720 27470 19748 28018
rect 19904 27470 19932 28018
rect 20088 27674 20116 29038
rect 20272 28558 20300 29446
rect 20364 28694 20392 30602
rect 20456 29696 20484 30806
rect 20548 30394 20576 30806
rect 20628 30660 20680 30666
rect 20628 30602 20680 30608
rect 20536 30388 20588 30394
rect 20536 30330 20588 30336
rect 20640 30258 20668 30602
rect 20628 30252 20680 30258
rect 20628 30194 20680 30200
rect 20628 30048 20680 30054
rect 20628 29990 20680 29996
rect 20536 29708 20588 29714
rect 20456 29668 20536 29696
rect 20456 28762 20484 29668
rect 20536 29650 20588 29656
rect 20640 29646 20668 29990
rect 20628 29640 20680 29646
rect 20626 29608 20628 29617
rect 20680 29608 20682 29617
rect 20626 29543 20682 29552
rect 20628 29232 20680 29238
rect 20628 29174 20680 29180
rect 20536 28960 20588 28966
rect 20536 28902 20588 28908
rect 20444 28756 20496 28762
rect 20444 28698 20496 28704
rect 20352 28688 20404 28694
rect 20352 28630 20404 28636
rect 20548 28626 20576 28902
rect 20536 28620 20588 28626
rect 20536 28562 20588 28568
rect 20640 28558 20668 29174
rect 20260 28552 20312 28558
rect 20260 28494 20312 28500
rect 20628 28552 20680 28558
rect 20628 28494 20680 28500
rect 20640 28218 20668 28494
rect 20628 28212 20680 28218
rect 20628 28154 20680 28160
rect 20076 27668 20128 27674
rect 20076 27610 20128 27616
rect 19708 27464 19760 27470
rect 19708 27406 19760 27412
rect 19892 27464 19944 27470
rect 19944 27424 20024 27452
rect 19892 27406 19944 27412
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19996 27130 20024 27424
rect 20168 27396 20220 27402
rect 20168 27338 20220 27344
rect 18604 27124 18656 27130
rect 18604 27066 18656 27072
rect 19984 27124 20036 27130
rect 19984 27066 20036 27072
rect 19616 27056 19668 27062
rect 19616 26998 19668 27004
rect 19628 26586 19656 26998
rect 20180 26586 20208 27338
rect 20536 27328 20588 27334
rect 20536 27270 20588 27276
rect 20350 27160 20406 27169
rect 20350 27095 20406 27104
rect 20364 27062 20392 27095
rect 20352 27056 20404 27062
rect 20352 26998 20404 27004
rect 19616 26580 19668 26586
rect 19616 26522 19668 26528
rect 20168 26580 20220 26586
rect 20168 26522 20220 26528
rect 19628 26382 19656 26522
rect 19616 26376 19668 26382
rect 19616 26318 19668 26324
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 15752 21888 15804 21894
rect 15752 21830 15804 21836
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 15476 3460 15528 3466
rect 15476 3402 15528 3408
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 16764 2848 16816 2854
rect 16764 2790 16816 2796
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 19708 2848 19760 2854
rect 19708 2790 19760 2796
rect 15198 2544 15254 2553
rect 15198 2479 15254 2488
rect 15212 2446 15240 2479
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 16776 2378 16804 2790
rect 16764 2372 16816 2378
rect 16764 2314 16816 2320
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 13360 1896 13412 1902
rect 13360 1838 13412 1844
rect 14844 800 14872 2246
rect 16776 800 16804 2314
rect 17224 2304 17276 2310
rect 17224 2246 17276 2252
rect 17236 2038 17264 2246
rect 17224 2032 17276 2038
rect 17224 1974 17276 1980
rect 18708 800 18736 2790
rect 19720 2446 19748 2790
rect 19708 2440 19760 2446
rect 19708 2382 19760 2388
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 20364 1834 20392 26998
rect 20548 26994 20576 27270
rect 20536 26988 20588 26994
rect 20536 26930 20588 26936
rect 20548 26382 20576 26930
rect 20536 26376 20588 26382
rect 20536 26318 20588 26324
rect 20548 25702 20576 26318
rect 20536 25696 20588 25702
rect 20536 25638 20588 25644
rect 20548 2514 20576 25638
rect 20720 2848 20772 2854
rect 20720 2790 20772 2796
rect 20536 2508 20588 2514
rect 20536 2450 20588 2456
rect 20732 2446 20760 2790
rect 20916 2650 20944 42162
rect 21376 41682 21404 42180
rect 21456 42162 21508 42168
rect 21548 42220 21600 42226
rect 21548 42162 21600 42168
rect 21652 42022 21680 42842
rect 21928 42770 21956 43046
rect 22112 42770 22140 43590
rect 21916 42764 21968 42770
rect 21916 42706 21968 42712
rect 22100 42764 22152 42770
rect 22100 42706 22152 42712
rect 21824 42696 21876 42702
rect 21824 42638 21876 42644
rect 21836 42362 21864 42638
rect 21824 42356 21876 42362
rect 21824 42298 21876 42304
rect 21732 42288 21784 42294
rect 21732 42230 21784 42236
rect 21640 42016 21692 42022
rect 21640 41958 21692 41964
rect 21364 41676 21416 41682
rect 21364 41618 21416 41624
rect 21744 41614 21772 42230
rect 21928 42158 21956 42706
rect 22006 42664 22062 42673
rect 22006 42599 22008 42608
rect 22060 42599 22062 42608
rect 22008 42570 22060 42576
rect 22192 42560 22244 42566
rect 22192 42502 22244 42508
rect 22008 42220 22060 42226
rect 22008 42162 22060 42168
rect 21916 42152 21968 42158
rect 21916 42094 21968 42100
rect 21916 42016 21968 42022
rect 21916 41958 21968 41964
rect 21732 41608 21784 41614
rect 21732 41550 21784 41556
rect 21088 41472 21140 41478
rect 21088 41414 21140 41420
rect 21100 41313 21128 41414
rect 21086 41304 21142 41313
rect 21086 41239 21142 41248
rect 21100 40526 21128 41239
rect 21744 41070 21772 41550
rect 21822 41304 21878 41313
rect 21822 41239 21878 41248
rect 21836 41138 21864 41239
rect 21824 41132 21876 41138
rect 21824 41074 21876 41080
rect 21272 41064 21324 41070
rect 21272 41006 21324 41012
rect 21732 41064 21784 41070
rect 21732 41006 21784 41012
rect 21284 40526 21312 41006
rect 21088 40520 21140 40526
rect 21088 40462 21140 40468
rect 21272 40520 21324 40526
rect 21272 40462 21324 40468
rect 21836 40225 21864 41074
rect 21928 40526 21956 41958
rect 22020 41274 22048 42162
rect 22008 41268 22060 41274
rect 22008 41210 22060 41216
rect 21916 40520 21968 40526
rect 21916 40462 21968 40468
rect 21822 40216 21878 40225
rect 21822 40151 21878 40160
rect 22020 40050 22048 41210
rect 22098 40488 22154 40497
rect 22204 40458 22232 42502
rect 22480 42226 22508 43590
rect 22756 42634 22784 43726
rect 22836 43716 22888 43722
rect 22836 43658 22888 43664
rect 22848 42634 22876 43658
rect 22744 42628 22796 42634
rect 22744 42570 22796 42576
rect 22836 42628 22888 42634
rect 22836 42570 22888 42576
rect 22560 42560 22612 42566
rect 22560 42502 22612 42508
rect 22572 42226 22600 42502
rect 22284 42220 22336 42226
rect 22284 42162 22336 42168
rect 22468 42220 22520 42226
rect 22468 42162 22520 42168
rect 22560 42220 22612 42226
rect 22560 42162 22612 42168
rect 22296 41818 22324 42162
rect 22374 41984 22430 41993
rect 22374 41919 22430 41928
rect 22284 41812 22336 41818
rect 22284 41754 22336 41760
rect 22282 41168 22338 41177
rect 22282 41103 22338 41112
rect 22098 40423 22154 40432
rect 22192 40452 22244 40458
rect 21180 40044 21232 40050
rect 21180 39986 21232 39992
rect 22008 40044 22060 40050
rect 22008 39986 22060 39992
rect 21192 39642 21220 39986
rect 22006 39944 22062 39953
rect 22006 39879 22062 39888
rect 21824 39840 21876 39846
rect 21824 39782 21876 39788
rect 21180 39636 21232 39642
rect 21180 39578 21232 39584
rect 21836 39506 21864 39782
rect 21824 39500 21876 39506
rect 21824 39442 21876 39448
rect 20996 39092 21048 39098
rect 20996 39034 21048 39040
rect 21008 38978 21036 39034
rect 21008 38950 21128 38978
rect 21100 38758 21128 38950
rect 21916 38956 21968 38962
rect 21916 38898 21968 38904
rect 21088 38752 21140 38758
rect 21088 38694 21140 38700
rect 21928 38554 21956 38898
rect 22020 38894 22048 39879
rect 22112 39438 22140 40423
rect 22192 40394 22244 40400
rect 22204 39982 22232 40394
rect 22192 39976 22244 39982
rect 22192 39918 22244 39924
rect 22296 39846 22324 41103
rect 22284 39840 22336 39846
rect 22284 39782 22336 39788
rect 22100 39432 22152 39438
rect 22100 39374 22152 39380
rect 22008 38888 22060 38894
rect 22060 38848 22140 38876
rect 22008 38830 22060 38836
rect 21916 38548 21968 38554
rect 21916 38490 21968 38496
rect 21824 38480 21876 38486
rect 21876 38428 22048 38434
rect 21824 38422 22048 38428
rect 21836 38406 22048 38422
rect 21916 38344 21968 38350
rect 21916 38286 21968 38292
rect 21824 38208 21876 38214
rect 21824 38150 21876 38156
rect 21456 38004 21508 38010
rect 21456 37946 21508 37952
rect 21468 37262 21496 37946
rect 21836 37806 21864 38150
rect 21732 37800 21784 37806
rect 21732 37742 21784 37748
rect 21824 37800 21876 37806
rect 21824 37742 21876 37748
rect 21640 37732 21692 37738
rect 21640 37674 21692 37680
rect 21652 37398 21680 37674
rect 21640 37392 21692 37398
rect 21640 37334 21692 37340
rect 21548 37324 21600 37330
rect 21548 37266 21600 37272
rect 21456 37256 21508 37262
rect 21456 37198 21508 37204
rect 21560 37097 21588 37266
rect 21744 37262 21772 37742
rect 21824 37664 21876 37670
rect 21824 37606 21876 37612
rect 21836 37466 21864 37606
rect 21824 37460 21876 37466
rect 21824 37402 21876 37408
rect 21732 37256 21784 37262
rect 21732 37198 21784 37204
rect 21546 37088 21602 37097
rect 21546 37023 21602 37032
rect 21732 36304 21784 36310
rect 21732 36246 21784 36252
rect 21456 36236 21508 36242
rect 21456 36178 21508 36184
rect 21468 36145 21496 36178
rect 21454 36136 21510 36145
rect 21454 36071 21510 36080
rect 21456 36032 21508 36038
rect 21456 35974 21508 35980
rect 21468 35698 21496 35974
rect 21456 35692 21508 35698
rect 21456 35634 21508 35640
rect 21088 35148 21140 35154
rect 21088 35090 21140 35096
rect 21456 35148 21508 35154
rect 21456 35090 21508 35096
rect 21100 34610 21128 35090
rect 21272 34672 21324 34678
rect 21272 34614 21324 34620
rect 21088 34604 21140 34610
rect 21088 34546 21140 34552
rect 20996 33924 21048 33930
rect 20996 33866 21048 33872
rect 21008 32910 21036 33866
rect 21100 33590 21128 34546
rect 21088 33584 21140 33590
rect 21088 33526 21140 33532
rect 21284 33386 21312 34614
rect 21468 33998 21496 35090
rect 21548 35080 21600 35086
rect 21548 35022 21600 35028
rect 21640 35080 21692 35086
rect 21640 35022 21692 35028
rect 21560 33998 21588 35022
rect 21652 34746 21680 35022
rect 21640 34740 21692 34746
rect 21640 34682 21692 34688
rect 21652 34202 21680 34682
rect 21640 34196 21692 34202
rect 21640 34138 21692 34144
rect 21456 33992 21508 33998
rect 21456 33934 21508 33940
rect 21548 33992 21600 33998
rect 21548 33934 21600 33940
rect 21272 33380 21324 33386
rect 21272 33322 21324 33328
rect 20996 32904 21048 32910
rect 20996 32846 21048 32852
rect 21008 32434 21036 32846
rect 21468 32434 21496 33934
rect 21744 32910 21772 36246
rect 21928 35834 21956 38286
rect 22020 37670 22048 38406
rect 22008 37664 22060 37670
rect 22008 37606 22060 37612
rect 22112 37466 22140 38848
rect 22296 38350 22324 39782
rect 22388 39642 22416 41919
rect 22572 41614 22600 42162
rect 22560 41608 22612 41614
rect 22560 41550 22612 41556
rect 22744 41132 22796 41138
rect 22744 41074 22796 41080
rect 22756 40594 22784 41074
rect 22744 40588 22796 40594
rect 22744 40530 22796 40536
rect 22376 39636 22428 39642
rect 22376 39578 22428 39584
rect 22652 39500 22704 39506
rect 22652 39442 22704 39448
rect 22284 38344 22336 38350
rect 22284 38286 22336 38292
rect 22468 37868 22520 37874
rect 22468 37810 22520 37816
rect 22192 37800 22244 37806
rect 22192 37742 22244 37748
rect 22100 37460 22152 37466
rect 22100 37402 22152 37408
rect 22100 37324 22152 37330
rect 22204 37312 22232 37742
rect 22152 37284 22232 37312
rect 22100 37266 22152 37272
rect 22112 36922 22140 37266
rect 22192 37120 22244 37126
rect 22192 37062 22244 37068
rect 22100 36916 22152 36922
rect 22100 36858 22152 36864
rect 21916 35828 21968 35834
rect 21916 35770 21968 35776
rect 22204 34542 22232 37062
rect 22480 36854 22508 37810
rect 22664 36922 22692 39442
rect 22744 38752 22796 38758
rect 22744 38694 22796 38700
rect 22756 38554 22784 38694
rect 22744 38548 22796 38554
rect 22744 38490 22796 38496
rect 22836 38548 22888 38554
rect 22836 38490 22888 38496
rect 22848 38282 22876 38490
rect 22836 38276 22888 38282
rect 22836 38218 22888 38224
rect 22836 37120 22888 37126
rect 22836 37062 22888 37068
rect 22652 36916 22704 36922
rect 22652 36858 22704 36864
rect 22468 36848 22520 36854
rect 22468 36790 22520 36796
rect 22848 36718 22876 37062
rect 22284 36712 22336 36718
rect 22284 36654 22336 36660
rect 22376 36712 22428 36718
rect 22376 36654 22428 36660
rect 22836 36712 22888 36718
rect 22836 36654 22888 36660
rect 22296 35290 22324 36654
rect 22388 35698 22416 36654
rect 22744 36372 22796 36378
rect 22744 36314 22796 36320
rect 22756 36174 22784 36314
rect 22848 36242 22876 36654
rect 22836 36236 22888 36242
rect 22836 36178 22888 36184
rect 22744 36168 22796 36174
rect 22744 36110 22796 36116
rect 22756 36038 22784 36110
rect 22468 36032 22520 36038
rect 22468 35974 22520 35980
rect 22744 36032 22796 36038
rect 22744 35974 22796 35980
rect 22376 35692 22428 35698
rect 22376 35634 22428 35640
rect 22388 35494 22416 35634
rect 22376 35488 22428 35494
rect 22376 35430 22428 35436
rect 22284 35284 22336 35290
rect 22284 35226 22336 35232
rect 22376 34604 22428 34610
rect 22376 34546 22428 34552
rect 22192 34536 22244 34542
rect 22192 34478 22244 34484
rect 22008 34400 22060 34406
rect 22008 34342 22060 34348
rect 21914 33280 21970 33289
rect 21914 33215 21970 33224
rect 21928 32910 21956 33215
rect 21732 32904 21784 32910
rect 21732 32846 21784 32852
rect 21916 32904 21968 32910
rect 21916 32846 21968 32852
rect 20996 32428 21048 32434
rect 20996 32370 21048 32376
rect 21456 32428 21508 32434
rect 21456 32370 21508 32376
rect 21008 31346 21036 32370
rect 21088 31816 21140 31822
rect 21088 31758 21140 31764
rect 21100 31482 21128 31758
rect 21088 31476 21140 31482
rect 21088 31418 21140 31424
rect 21468 31414 21496 32370
rect 21744 31822 21772 32846
rect 21824 32836 21876 32842
rect 21824 32778 21876 32784
rect 21836 32502 21864 32778
rect 21824 32496 21876 32502
rect 21824 32438 21876 32444
rect 21732 31816 21784 31822
rect 21732 31758 21784 31764
rect 21456 31408 21508 31414
rect 21456 31350 21508 31356
rect 20996 31340 21048 31346
rect 20996 31282 21048 31288
rect 21008 30938 21036 31282
rect 21468 30938 21496 31350
rect 20996 30932 21048 30938
rect 20996 30874 21048 30880
rect 21456 30932 21508 30938
rect 21456 30874 21508 30880
rect 21180 30796 21232 30802
rect 21180 30738 21232 30744
rect 20996 30592 21048 30598
rect 20996 30534 21048 30540
rect 21008 30258 21036 30534
rect 21192 30326 21220 30738
rect 21272 30728 21324 30734
rect 21272 30670 21324 30676
rect 21180 30320 21232 30326
rect 21180 30262 21232 30268
rect 20996 30252 21048 30258
rect 20996 30194 21048 30200
rect 21192 29850 21220 30262
rect 21284 30258 21312 30670
rect 21744 30598 21772 31758
rect 21928 31754 21956 32846
rect 22020 32502 22048 34342
rect 22204 33114 22232 34478
rect 22284 33584 22336 33590
rect 22284 33526 22336 33532
rect 22192 33108 22244 33114
rect 22192 33050 22244 33056
rect 22008 32496 22060 32502
rect 22008 32438 22060 32444
rect 21916 31748 21968 31754
rect 21916 31690 21968 31696
rect 21732 30592 21784 30598
rect 21732 30534 21784 30540
rect 21272 30252 21324 30258
rect 21272 30194 21324 30200
rect 21180 29844 21232 29850
rect 21180 29786 21232 29792
rect 20996 29640 21048 29646
rect 21928 29594 21956 31690
rect 22020 31346 22048 32438
rect 22100 32428 22152 32434
rect 22100 32370 22152 32376
rect 22112 31686 22140 32370
rect 22204 32230 22232 33050
rect 22296 32774 22324 33526
rect 22388 32910 22416 34546
rect 22480 33590 22508 35974
rect 22560 35692 22612 35698
rect 22560 35634 22612 35640
rect 22572 35222 22600 35634
rect 22744 35488 22796 35494
rect 22744 35430 22796 35436
rect 22560 35216 22612 35222
rect 22560 35158 22612 35164
rect 22756 35154 22784 35430
rect 22744 35148 22796 35154
rect 22744 35090 22796 35096
rect 22560 35080 22612 35086
rect 22560 35022 22612 35028
rect 22572 34202 22600 35022
rect 22560 34196 22612 34202
rect 22940 34184 22968 44134
rect 23400 43790 23428 46106
rect 23584 45898 23612 46446
rect 23572 45892 23624 45898
rect 23572 45834 23624 45840
rect 23584 45490 23612 45834
rect 23572 45484 23624 45490
rect 23572 45426 23624 45432
rect 24412 45422 24440 46514
rect 24596 46374 24624 46990
rect 24964 46578 24992 46990
rect 25516 46578 25544 49286
rect 27066 49200 27122 50000
rect 28998 49200 29054 50000
rect 30930 49200 30986 50000
rect 32862 49200 32918 50000
rect 34794 49200 34850 50000
rect 36726 49314 36782 50000
rect 36726 49286 37228 49314
rect 36726 49200 36782 49286
rect 26240 47660 26292 47666
rect 26240 47602 26292 47608
rect 26424 47660 26476 47666
rect 26424 47602 26476 47608
rect 26252 47530 26280 47602
rect 26240 47524 26292 47530
rect 26240 47466 26292 47472
rect 26436 47258 26464 47602
rect 26884 47524 26936 47530
rect 26884 47466 26936 47472
rect 26424 47252 26476 47258
rect 26424 47194 26476 47200
rect 26148 46912 26200 46918
rect 26148 46854 26200 46860
rect 25964 46640 26016 46646
rect 25964 46582 26016 46588
rect 24952 46572 25004 46578
rect 24952 46514 25004 46520
rect 25228 46572 25280 46578
rect 25228 46514 25280 46520
rect 25504 46572 25556 46578
rect 25504 46514 25556 46520
rect 24584 46368 24636 46374
rect 24584 46310 24636 46316
rect 24492 45960 24544 45966
rect 24490 45928 24492 45937
rect 24544 45928 24546 45937
rect 24490 45863 24546 45872
rect 24492 45824 24544 45830
rect 24492 45766 24544 45772
rect 24504 45490 24532 45766
rect 24492 45484 24544 45490
rect 24492 45426 24544 45432
rect 24032 45416 24084 45422
rect 24032 45358 24084 45364
rect 24400 45416 24452 45422
rect 24400 45358 24452 45364
rect 23480 45280 23532 45286
rect 23480 45222 23532 45228
rect 23940 45280 23992 45286
rect 23940 45222 23992 45228
rect 23492 45014 23520 45222
rect 23480 45008 23532 45014
rect 23480 44950 23532 44956
rect 23480 44736 23532 44742
rect 23480 44678 23532 44684
rect 23756 44736 23808 44742
rect 23756 44678 23808 44684
rect 23492 44334 23520 44678
rect 23768 44538 23796 44678
rect 23756 44532 23808 44538
rect 23756 44474 23808 44480
rect 23768 44402 23796 44474
rect 23952 44402 23980 45222
rect 24044 45082 24072 45358
rect 24596 45082 24624 46310
rect 24964 46034 24992 46514
rect 24952 46028 25004 46034
rect 24952 45970 25004 45976
rect 24768 45960 24820 45966
rect 24768 45902 24820 45908
rect 24032 45076 24084 45082
rect 24032 45018 24084 45024
rect 24584 45076 24636 45082
rect 24584 45018 24636 45024
rect 24780 44470 24808 45902
rect 25136 45892 25188 45898
rect 25136 45834 25188 45840
rect 25044 45416 25096 45422
rect 25044 45358 25096 45364
rect 24860 45348 24912 45354
rect 24860 45290 24912 45296
rect 24768 44464 24820 44470
rect 24768 44406 24820 44412
rect 24872 44402 24900 45290
rect 25056 44878 25084 45358
rect 25044 44872 25096 44878
rect 25044 44814 25096 44820
rect 23756 44396 23808 44402
rect 23676 44356 23756 44384
rect 23480 44328 23532 44334
rect 23480 44270 23532 44276
rect 23388 43784 23440 43790
rect 23388 43726 23440 43732
rect 23204 43648 23256 43654
rect 23204 43590 23256 43596
rect 23216 42906 23244 43590
rect 23388 43308 23440 43314
rect 23388 43250 23440 43256
rect 23204 42900 23256 42906
rect 23204 42842 23256 42848
rect 23112 41744 23164 41750
rect 23112 41686 23164 41692
rect 23124 41478 23152 41686
rect 23112 41472 23164 41478
rect 23112 41414 23164 41420
rect 23020 41268 23072 41274
rect 23020 41210 23072 41216
rect 23032 40526 23060 41210
rect 23020 40520 23072 40526
rect 23020 40462 23072 40468
rect 23020 40044 23072 40050
rect 23020 39986 23072 39992
rect 23032 38962 23060 39986
rect 23124 39098 23152 41414
rect 23216 40186 23244 42842
rect 23296 42288 23348 42294
rect 23296 42230 23348 42236
rect 23204 40180 23256 40186
rect 23204 40122 23256 40128
rect 23216 39250 23244 40122
rect 23308 39386 23336 42230
rect 23400 39506 23428 43250
rect 23480 42764 23532 42770
rect 23676 42752 23704 44356
rect 23940 44396 23992 44402
rect 23756 44338 23808 44344
rect 23860 44356 23940 44384
rect 23756 43648 23808 43654
rect 23756 43590 23808 43596
rect 23768 43382 23796 43590
rect 23756 43376 23808 43382
rect 23756 43318 23808 43324
rect 23532 42724 23704 42752
rect 23480 42706 23532 42712
rect 23756 42696 23808 42702
rect 23860 42684 23888 44356
rect 23940 44338 23992 44344
rect 24860 44396 24912 44402
rect 24912 44356 24992 44384
rect 24860 44338 24912 44344
rect 24768 44328 24820 44334
rect 24768 44270 24820 44276
rect 23940 44192 23992 44198
rect 23940 44134 23992 44140
rect 24400 44192 24452 44198
rect 24780 44180 24808 44270
rect 24780 44152 24900 44180
rect 24400 44134 24452 44140
rect 23808 42656 23888 42684
rect 23756 42638 23808 42644
rect 23952 41614 23980 44134
rect 24124 43716 24176 43722
rect 24124 43658 24176 43664
rect 24032 43308 24084 43314
rect 24032 43250 24084 43256
rect 24044 42770 24072 43250
rect 24032 42764 24084 42770
rect 24032 42706 24084 42712
rect 24032 42628 24084 42634
rect 24032 42570 24084 42576
rect 24044 42362 24072 42570
rect 24032 42356 24084 42362
rect 24032 42298 24084 42304
rect 23940 41608 23992 41614
rect 23940 41550 23992 41556
rect 23480 41472 23532 41478
rect 23480 41414 23532 41420
rect 23492 41206 23520 41414
rect 23480 41200 23532 41206
rect 23480 41142 23532 41148
rect 23848 41064 23900 41070
rect 23848 41006 23900 41012
rect 23860 40662 23888 41006
rect 24032 40996 24084 41002
rect 24032 40938 24084 40944
rect 23848 40656 23900 40662
rect 23848 40598 23900 40604
rect 23756 40520 23808 40526
rect 23756 40462 23808 40468
rect 23664 40384 23716 40390
rect 23664 40326 23716 40332
rect 23676 40186 23704 40326
rect 23664 40180 23716 40186
rect 23664 40122 23716 40128
rect 23572 40044 23624 40050
rect 23572 39986 23624 39992
rect 23388 39500 23440 39506
rect 23440 39460 23520 39488
rect 23388 39442 23440 39448
rect 23308 39358 23428 39386
rect 23216 39222 23336 39250
rect 23112 39092 23164 39098
rect 23164 39052 23244 39080
rect 23112 39034 23164 39040
rect 23020 38956 23072 38962
rect 23072 38916 23152 38944
rect 23020 38898 23072 38904
rect 23020 38480 23072 38486
rect 23020 38422 23072 38428
rect 23032 37262 23060 38422
rect 23124 38214 23152 38916
rect 23216 38554 23244 39052
rect 23308 39030 23336 39222
rect 23296 39024 23348 39030
rect 23296 38966 23348 38972
rect 23204 38548 23256 38554
rect 23204 38490 23256 38496
rect 23308 38350 23336 38966
rect 23296 38344 23348 38350
rect 23296 38286 23348 38292
rect 23112 38208 23164 38214
rect 23296 38208 23348 38214
rect 23112 38150 23164 38156
rect 23216 38168 23296 38196
rect 23124 37806 23152 38150
rect 23216 38010 23244 38168
rect 23296 38150 23348 38156
rect 23204 38004 23256 38010
rect 23204 37946 23256 37952
rect 23296 37936 23348 37942
rect 23294 37904 23296 37913
rect 23348 37904 23350 37913
rect 23294 37839 23350 37848
rect 23112 37800 23164 37806
rect 23112 37742 23164 37748
rect 23124 37398 23152 37742
rect 23112 37392 23164 37398
rect 23112 37334 23164 37340
rect 23400 37330 23428 39358
rect 23492 38350 23520 39460
rect 23584 39098 23612 39986
rect 23572 39092 23624 39098
rect 23572 39034 23624 39040
rect 23664 38888 23716 38894
rect 23664 38830 23716 38836
rect 23480 38344 23532 38350
rect 23480 38286 23532 38292
rect 23676 38162 23704 38830
rect 23584 38134 23704 38162
rect 23388 37324 23440 37330
rect 23388 37266 23440 37272
rect 23020 37256 23072 37262
rect 23020 37198 23072 37204
rect 23032 36718 23060 37198
rect 23400 36786 23428 37266
rect 23388 36780 23440 36786
rect 23388 36722 23440 36728
rect 23584 36718 23612 38134
rect 23020 36712 23072 36718
rect 23020 36654 23072 36660
rect 23572 36712 23624 36718
rect 23572 36654 23624 36660
rect 23480 36032 23532 36038
rect 23480 35974 23532 35980
rect 23664 36032 23716 36038
rect 23664 35974 23716 35980
rect 23018 35864 23074 35873
rect 23018 35799 23074 35808
rect 23032 35154 23060 35799
rect 23020 35148 23072 35154
rect 23020 35090 23072 35096
rect 23112 35080 23164 35086
rect 23112 35022 23164 35028
rect 23124 34746 23152 35022
rect 23112 34740 23164 34746
rect 23112 34682 23164 34688
rect 23492 34678 23520 35974
rect 23572 35488 23624 35494
rect 23572 35430 23624 35436
rect 23480 34672 23532 34678
rect 23480 34614 23532 34620
rect 23480 34536 23532 34542
rect 23584 34490 23612 35430
rect 23676 34610 23704 35974
rect 23768 35562 23796 40462
rect 24044 40390 24072 40938
rect 24032 40384 24084 40390
rect 24032 40326 24084 40332
rect 23938 40216 23994 40225
rect 23938 40151 23994 40160
rect 23952 40118 23980 40151
rect 23940 40112 23992 40118
rect 23940 40054 23992 40060
rect 24044 39982 24072 40326
rect 24032 39976 24084 39982
rect 24032 39918 24084 39924
rect 23940 39568 23992 39574
rect 23940 39510 23992 39516
rect 23846 38584 23902 38593
rect 23846 38519 23848 38528
rect 23900 38519 23902 38528
rect 23848 38490 23900 38496
rect 23860 38010 23888 38490
rect 23848 38004 23900 38010
rect 23848 37946 23900 37952
rect 23860 37641 23888 37946
rect 23846 37632 23902 37641
rect 23846 37567 23902 37576
rect 23860 37398 23888 37567
rect 23952 37466 23980 39510
rect 24032 39024 24084 39030
rect 24032 38966 24084 38972
rect 24044 37874 24072 38966
rect 24032 37868 24084 37874
rect 24032 37810 24084 37816
rect 24030 37768 24086 37777
rect 24030 37703 24086 37712
rect 23940 37460 23992 37466
rect 23940 37402 23992 37408
rect 23848 37392 23900 37398
rect 23848 37334 23900 37340
rect 23848 37256 23900 37262
rect 23848 37198 23900 37204
rect 23860 36922 23888 37198
rect 23848 36916 23900 36922
rect 23848 36858 23900 36864
rect 23952 36854 23980 37402
rect 24044 36961 24072 37703
rect 24136 37670 24164 43658
rect 24412 43178 24440 44134
rect 24768 43920 24820 43926
rect 24768 43862 24820 43868
rect 24492 43852 24544 43858
rect 24492 43794 24544 43800
rect 24504 43246 24532 43794
rect 24780 43382 24808 43862
rect 24872 43722 24900 44152
rect 24964 43790 24992 44356
rect 25044 44192 25096 44198
rect 25044 44134 25096 44140
rect 24952 43784 25004 43790
rect 24952 43726 25004 43732
rect 24860 43716 24912 43722
rect 24860 43658 24912 43664
rect 24768 43376 24820 43382
rect 24768 43318 24820 43324
rect 24492 43240 24544 43246
rect 24492 43182 24544 43188
rect 24400 43172 24452 43178
rect 24400 43114 24452 43120
rect 24412 42226 24440 43114
rect 24504 42770 24532 43182
rect 24492 42764 24544 42770
rect 24492 42706 24544 42712
rect 24400 42220 24452 42226
rect 24400 42162 24452 42168
rect 24504 41682 24532 42706
rect 24676 42696 24728 42702
rect 24780 42684 24808 43318
rect 24860 42696 24912 42702
rect 24780 42656 24860 42684
rect 24676 42638 24728 42644
rect 24860 42638 24912 42644
rect 24584 42560 24636 42566
rect 24584 42502 24636 42508
rect 24596 42226 24624 42502
rect 24584 42220 24636 42226
rect 24584 42162 24636 42168
rect 24492 41676 24544 41682
rect 24492 41618 24544 41624
rect 24688 41614 24716 42638
rect 24860 42560 24912 42566
rect 24860 42502 24912 42508
rect 24872 42362 24900 42502
rect 24860 42356 24912 42362
rect 24860 42298 24912 42304
rect 25056 42242 25084 44134
rect 24872 42214 25084 42242
rect 24676 41608 24728 41614
rect 24676 41550 24728 41556
rect 24216 41472 24268 41478
rect 24216 41414 24268 41420
rect 24228 40526 24256 41414
rect 24308 41268 24360 41274
rect 24308 41210 24360 41216
rect 24216 40520 24268 40526
rect 24216 40462 24268 40468
rect 24228 39438 24256 40462
rect 24216 39432 24268 39438
rect 24216 39374 24268 39380
rect 24228 38026 24256 39374
rect 24320 38962 24348 41210
rect 24400 41132 24452 41138
rect 24400 41074 24452 41080
rect 24492 41132 24544 41138
rect 24492 41074 24544 41080
rect 24308 38956 24360 38962
rect 24308 38898 24360 38904
rect 24320 38214 24348 38898
rect 24308 38208 24360 38214
rect 24308 38150 24360 38156
rect 24228 37998 24348 38026
rect 24412 38010 24440 41074
rect 24504 39642 24532 41074
rect 24674 41032 24730 41041
rect 24674 40967 24676 40976
rect 24728 40967 24730 40976
rect 24676 40938 24728 40944
rect 24584 40928 24636 40934
rect 24584 40870 24636 40876
rect 24768 40928 24820 40934
rect 24768 40870 24820 40876
rect 24596 40526 24624 40870
rect 24780 40730 24808 40870
rect 24768 40724 24820 40730
rect 24768 40666 24820 40672
rect 24584 40520 24636 40526
rect 24584 40462 24636 40468
rect 24492 39636 24544 39642
rect 24492 39578 24544 39584
rect 24596 39506 24624 40462
rect 24872 40458 24900 42214
rect 24952 41132 25004 41138
rect 24952 41074 25004 41080
rect 24964 40730 24992 41074
rect 24952 40724 25004 40730
rect 24952 40666 25004 40672
rect 24768 40452 24820 40458
rect 24768 40394 24820 40400
rect 24860 40452 24912 40458
rect 24860 40394 24912 40400
rect 24780 40186 24808 40394
rect 24768 40180 24820 40186
rect 24768 40122 24820 40128
rect 24676 39840 24728 39846
rect 24676 39782 24728 39788
rect 24584 39500 24636 39506
rect 24584 39442 24636 39448
rect 24492 38888 24544 38894
rect 24492 38830 24544 38836
rect 24216 37868 24268 37874
rect 24216 37810 24268 37816
rect 24124 37664 24176 37670
rect 24124 37606 24176 37612
rect 24124 37392 24176 37398
rect 24124 37334 24176 37340
rect 24030 36952 24086 36961
rect 24030 36887 24086 36896
rect 23940 36848 23992 36854
rect 23940 36790 23992 36796
rect 24044 35834 24072 36887
rect 24136 36786 24164 37334
rect 24124 36780 24176 36786
rect 24124 36722 24176 36728
rect 24032 35828 24084 35834
rect 24032 35770 24084 35776
rect 23756 35556 23808 35562
rect 23756 35498 23808 35504
rect 24044 34610 24072 35770
rect 24228 35766 24256 37810
rect 24320 37777 24348 37998
rect 24400 38004 24452 38010
rect 24400 37946 24452 37952
rect 24504 37874 24532 38830
rect 24584 38752 24636 38758
rect 24584 38694 24636 38700
rect 24492 37868 24544 37874
rect 24492 37810 24544 37816
rect 24596 37806 24624 38694
rect 24688 38049 24716 39782
rect 24872 39574 24900 40394
rect 24860 39568 24912 39574
rect 24860 39510 24912 39516
rect 24964 39284 24992 40666
rect 25044 40520 25096 40526
rect 25044 40462 25096 40468
rect 25056 39914 25084 40462
rect 25044 39908 25096 39914
rect 25044 39850 25096 39856
rect 25044 39296 25096 39302
rect 24964 39256 25044 39284
rect 25044 39238 25096 39244
rect 24860 39024 24912 39030
rect 24860 38966 24912 38972
rect 24768 38956 24820 38962
rect 24768 38898 24820 38904
rect 24780 38758 24808 38898
rect 24768 38752 24820 38758
rect 24768 38694 24820 38700
rect 24768 38344 24820 38350
rect 24768 38286 24820 38292
rect 24674 38040 24730 38049
rect 24674 37975 24730 37984
rect 24688 37874 24716 37975
rect 24676 37868 24728 37874
rect 24676 37810 24728 37816
rect 24400 37800 24452 37806
rect 24306 37768 24362 37777
rect 24400 37742 24452 37748
rect 24584 37800 24636 37806
rect 24584 37742 24636 37748
rect 24306 37703 24362 37712
rect 24412 37670 24440 37742
rect 24400 37664 24452 37670
rect 24400 37606 24452 37612
rect 24308 37392 24360 37398
rect 24308 37334 24360 37340
rect 24490 37360 24546 37369
rect 24320 36038 24348 37334
rect 24490 37295 24492 37304
rect 24544 37295 24546 37304
rect 24492 37266 24544 37272
rect 24400 37256 24452 37262
rect 24452 37204 24532 37210
rect 24400 37198 24532 37204
rect 24412 37182 24532 37198
rect 24308 36032 24360 36038
rect 24308 35974 24360 35980
rect 24216 35760 24268 35766
rect 24216 35702 24268 35708
rect 24504 35601 24532 37182
rect 24596 36786 24624 37742
rect 24780 37466 24808 38286
rect 24872 37874 24900 38966
rect 24952 38344 25004 38350
rect 24952 38286 25004 38292
rect 24860 37868 24912 37874
rect 24860 37810 24912 37816
rect 24860 37732 24912 37738
rect 24860 37674 24912 37680
rect 24768 37460 24820 37466
rect 24768 37402 24820 37408
rect 24676 36916 24728 36922
rect 24676 36858 24728 36864
rect 24584 36780 24636 36786
rect 24584 36722 24636 36728
rect 24688 35834 24716 36858
rect 24768 36848 24820 36854
rect 24768 36790 24820 36796
rect 24780 36038 24808 36790
rect 24768 36032 24820 36038
rect 24768 35974 24820 35980
rect 24676 35828 24728 35834
rect 24676 35770 24728 35776
rect 24676 35692 24728 35698
rect 24676 35634 24728 35640
rect 24490 35592 24546 35601
rect 24400 35556 24452 35562
rect 24490 35527 24546 35536
rect 24400 35498 24452 35504
rect 23664 34604 23716 34610
rect 23664 34546 23716 34552
rect 24032 34604 24084 34610
rect 24032 34546 24084 34552
rect 24216 34604 24268 34610
rect 24216 34546 24268 34552
rect 23532 34484 23612 34490
rect 23480 34478 23612 34484
rect 23492 34462 23612 34478
rect 22560 34138 22612 34144
rect 22756 34156 22968 34184
rect 22468 33584 22520 33590
rect 22468 33526 22520 33532
rect 22376 32904 22428 32910
rect 22652 32904 22704 32910
rect 22428 32864 22508 32892
rect 22376 32846 22428 32852
rect 22284 32768 22336 32774
rect 22284 32710 22336 32716
rect 22296 32434 22324 32710
rect 22284 32428 22336 32434
rect 22284 32370 22336 32376
rect 22480 32366 22508 32864
rect 22652 32846 22704 32852
rect 22664 32570 22692 32846
rect 22652 32564 22704 32570
rect 22652 32506 22704 32512
rect 22468 32360 22520 32366
rect 22468 32302 22520 32308
rect 22284 32292 22336 32298
rect 22284 32234 22336 32240
rect 22192 32224 22244 32230
rect 22192 32166 22244 32172
rect 22296 31958 22324 32234
rect 22664 31958 22692 32506
rect 22284 31952 22336 31958
rect 22652 31952 22704 31958
rect 22284 31894 22336 31900
rect 22572 31900 22652 31906
rect 22572 31894 22704 31900
rect 22376 31884 22428 31890
rect 22376 31826 22428 31832
rect 22572 31878 22692 31894
rect 22100 31680 22152 31686
rect 22100 31622 22152 31628
rect 22112 31414 22140 31622
rect 22100 31408 22152 31414
rect 22100 31350 22152 31356
rect 22008 31340 22060 31346
rect 22008 31282 22060 31288
rect 22006 31240 22062 31249
rect 22006 31175 22062 31184
rect 22020 31142 22048 31175
rect 22008 31136 22060 31142
rect 22008 31078 22060 31084
rect 22020 29646 22048 31078
rect 22112 30666 22140 31350
rect 22284 31340 22336 31346
rect 22284 31282 22336 31288
rect 22100 30660 22152 30666
rect 22100 30602 22152 30608
rect 22296 30394 22324 31282
rect 22388 30938 22416 31826
rect 22572 31414 22600 31878
rect 22756 31804 22784 34156
rect 24228 34134 24256 34546
rect 24216 34128 24268 34134
rect 24216 34070 24268 34076
rect 22928 34060 22980 34066
rect 22928 34002 22980 34008
rect 22836 33992 22888 33998
rect 22836 33934 22888 33940
rect 22848 33522 22876 33934
rect 22836 33516 22888 33522
rect 22836 33458 22888 33464
rect 22848 33114 22876 33458
rect 22940 33114 22968 34002
rect 24124 33652 24176 33658
rect 24124 33594 24176 33600
rect 23112 33516 23164 33522
rect 23112 33458 23164 33464
rect 23480 33516 23532 33522
rect 23480 33458 23532 33464
rect 22836 33108 22888 33114
rect 22836 33050 22888 33056
rect 22928 33108 22980 33114
rect 22928 33050 22980 33056
rect 23124 32910 23152 33458
rect 23296 33448 23348 33454
rect 23296 33390 23348 33396
rect 23308 33046 23336 33390
rect 23388 33108 23440 33114
rect 23388 33050 23440 33056
rect 23296 33040 23348 33046
rect 23296 32982 23348 32988
rect 23112 32904 23164 32910
rect 23112 32846 23164 32852
rect 23124 31890 23152 32846
rect 23400 32434 23428 33050
rect 23492 32910 23520 33458
rect 23480 32904 23532 32910
rect 23480 32846 23532 32852
rect 23388 32428 23440 32434
rect 23388 32370 23440 32376
rect 23296 32360 23348 32366
rect 23296 32302 23348 32308
rect 23112 31884 23164 31890
rect 23112 31826 23164 31832
rect 22664 31776 22784 31804
rect 22560 31408 22612 31414
rect 22560 31350 22612 31356
rect 22376 30932 22428 30938
rect 22376 30874 22428 30880
rect 22284 30388 22336 30394
rect 22284 30330 22336 30336
rect 22296 29714 22324 30330
rect 22284 29708 22336 29714
rect 22284 29650 22336 29656
rect 20996 29582 21048 29588
rect 21008 29306 21036 29582
rect 21836 29566 21956 29594
rect 22008 29640 22060 29646
rect 22008 29582 22060 29588
rect 22376 29572 22428 29578
rect 20996 29300 21048 29306
rect 20996 29242 21048 29248
rect 21088 29232 21140 29238
rect 21088 29174 21140 29180
rect 21100 28626 21128 29174
rect 21088 28620 21140 28626
rect 21088 28562 21140 28568
rect 20994 28112 21050 28121
rect 20994 28047 21050 28056
rect 21008 27606 21036 28047
rect 20996 27600 21048 27606
rect 20996 27542 21048 27548
rect 21548 27464 21600 27470
rect 21548 27406 21600 27412
rect 21560 27062 21588 27406
rect 21836 27130 21864 29566
rect 22376 29514 22428 29520
rect 21916 29504 21968 29510
rect 21916 29446 21968 29452
rect 21928 28558 21956 29446
rect 22008 29164 22060 29170
rect 22008 29106 22060 29112
rect 21916 28552 21968 28558
rect 21916 28494 21968 28500
rect 22020 27130 22048 29106
rect 22100 29096 22152 29102
rect 22100 29038 22152 29044
rect 22112 28490 22140 29038
rect 22388 28966 22416 29514
rect 22560 29504 22612 29510
rect 22560 29446 22612 29452
rect 22572 29306 22600 29446
rect 22560 29300 22612 29306
rect 22560 29242 22612 29248
rect 22376 28960 22428 28966
rect 22376 28902 22428 28908
rect 22100 28484 22152 28490
rect 22100 28426 22152 28432
rect 22112 27674 22140 28426
rect 22282 28112 22338 28121
rect 22282 28047 22284 28056
rect 22336 28047 22338 28056
rect 22284 28018 22336 28024
rect 22100 27668 22152 27674
rect 22100 27610 22152 27616
rect 22192 27600 22244 27606
rect 22192 27542 22244 27548
rect 21824 27124 21876 27130
rect 21824 27066 21876 27072
rect 22008 27124 22060 27130
rect 22008 27066 22060 27072
rect 21548 27056 21600 27062
rect 21548 26998 21600 27004
rect 21088 26988 21140 26994
rect 21088 26930 21140 26936
rect 21100 26586 21128 26930
rect 21088 26580 21140 26586
rect 21088 26522 21140 26528
rect 21836 26382 21864 27066
rect 22204 26586 22232 27542
rect 22284 27464 22336 27470
rect 22284 27406 22336 27412
rect 22296 26926 22324 27406
rect 22284 26920 22336 26926
rect 22284 26862 22336 26868
rect 22192 26580 22244 26586
rect 22192 26522 22244 26528
rect 22296 26450 22324 26862
rect 22468 26852 22520 26858
rect 22468 26794 22520 26800
rect 22284 26444 22336 26450
rect 22284 26386 22336 26392
rect 21824 26376 21876 26382
rect 21824 26318 21876 26324
rect 21836 26042 21864 26318
rect 22480 26314 22508 26794
rect 22468 26308 22520 26314
rect 22468 26250 22520 26256
rect 21824 26036 21876 26042
rect 21824 25978 21876 25984
rect 22480 25702 22508 26250
rect 22468 25696 22520 25702
rect 22468 25638 22520 25644
rect 22480 5574 22508 25638
rect 22664 22094 22692 31776
rect 23308 31482 23336 32302
rect 23492 32298 23520 32846
rect 23572 32496 23624 32502
rect 23572 32438 23624 32444
rect 23480 32292 23532 32298
rect 23480 32234 23532 32240
rect 23492 31822 23520 32234
rect 23584 31890 23612 32438
rect 23572 31884 23624 31890
rect 23572 31826 23624 31832
rect 23480 31816 23532 31822
rect 23480 31758 23532 31764
rect 23296 31476 23348 31482
rect 23296 31418 23348 31424
rect 23018 31240 23074 31249
rect 23018 31175 23074 31184
rect 23032 30258 23060 31175
rect 24136 30734 24164 33594
rect 24216 33380 24268 33386
rect 24216 33322 24268 33328
rect 24228 31482 24256 33322
rect 24308 31748 24360 31754
rect 24308 31690 24360 31696
rect 24216 31476 24268 31482
rect 24216 31418 24268 31424
rect 24124 30728 24176 30734
rect 24124 30670 24176 30676
rect 23756 30592 23808 30598
rect 23756 30534 23808 30540
rect 24032 30592 24084 30598
rect 24032 30534 24084 30540
rect 23020 30252 23072 30258
rect 23020 30194 23072 30200
rect 22836 29844 22888 29850
rect 22836 29786 22888 29792
rect 22848 29714 22876 29786
rect 22744 29708 22796 29714
rect 22744 29650 22796 29656
rect 22836 29708 22888 29714
rect 22836 29650 22888 29656
rect 22756 28626 22784 29650
rect 23032 29322 23060 30194
rect 23296 29708 23348 29714
rect 23296 29650 23348 29656
rect 23032 29294 23152 29322
rect 23308 29306 23336 29650
rect 23768 29646 23796 30534
rect 24044 30258 24072 30534
rect 24032 30252 24084 30258
rect 24032 30194 24084 30200
rect 23940 30184 23992 30190
rect 23940 30126 23992 30132
rect 23756 29640 23808 29646
rect 23756 29582 23808 29588
rect 23664 29504 23716 29510
rect 23664 29446 23716 29452
rect 23020 29164 23072 29170
rect 23020 29106 23072 29112
rect 22928 28960 22980 28966
rect 22928 28902 22980 28908
rect 22940 28694 22968 28902
rect 22928 28688 22980 28694
rect 22928 28630 22980 28636
rect 22744 28620 22796 28626
rect 22744 28562 22796 28568
rect 22940 27470 22968 28630
rect 23032 28490 23060 29106
rect 23124 28558 23152 29294
rect 23296 29300 23348 29306
rect 23296 29242 23348 29248
rect 23676 29170 23704 29446
rect 23952 29306 23980 30126
rect 23940 29300 23992 29306
rect 23940 29242 23992 29248
rect 23664 29164 23716 29170
rect 23664 29106 23716 29112
rect 24228 28762 24256 31418
rect 24320 30802 24348 31690
rect 24308 30796 24360 30802
rect 24308 30738 24360 30744
rect 24412 30190 24440 35498
rect 24504 35086 24532 35527
rect 24492 35080 24544 35086
rect 24492 35022 24544 35028
rect 24688 34746 24716 35634
rect 24780 35290 24808 35974
rect 24768 35284 24820 35290
rect 24768 35226 24820 35232
rect 24676 34740 24728 34746
rect 24676 34682 24728 34688
rect 24780 34610 24808 35226
rect 24872 35018 24900 37674
rect 24964 35698 24992 38286
rect 24952 35692 25004 35698
rect 24952 35634 25004 35640
rect 24964 35086 24992 35634
rect 24952 35080 25004 35086
rect 24952 35022 25004 35028
rect 24860 35012 24912 35018
rect 24860 34954 24912 34960
rect 25056 34746 25084 39238
rect 25148 38196 25176 45834
rect 25240 45665 25268 46514
rect 25976 46170 26004 46582
rect 25964 46164 26016 46170
rect 25964 46106 26016 46112
rect 25226 45656 25282 45665
rect 25976 45642 26004 46106
rect 26160 45830 26188 46854
rect 26608 46572 26660 46578
rect 26608 46514 26660 46520
rect 26424 46368 26476 46374
rect 26424 46310 26476 46316
rect 26238 45928 26294 45937
rect 26238 45863 26294 45872
rect 26148 45824 26200 45830
rect 26148 45766 26200 45772
rect 25976 45614 26096 45642
rect 26160 45626 26188 45766
rect 25226 45591 25282 45600
rect 25964 45484 26016 45490
rect 25964 45426 26016 45432
rect 25502 45384 25558 45393
rect 25502 45319 25558 45328
rect 25320 44464 25372 44470
rect 25320 44406 25372 44412
rect 25332 41562 25360 44406
rect 25516 44266 25544 45319
rect 25976 45082 26004 45426
rect 25964 45076 26016 45082
rect 25964 45018 26016 45024
rect 25780 45008 25832 45014
rect 25780 44950 25832 44956
rect 25792 44742 25820 44950
rect 26068 44878 26096 45614
rect 26148 45620 26200 45626
rect 26148 45562 26200 45568
rect 26252 45490 26280 45863
rect 26240 45484 26292 45490
rect 26240 45426 26292 45432
rect 26056 44872 26108 44878
rect 26056 44814 26108 44820
rect 25780 44736 25832 44742
rect 25780 44678 25832 44684
rect 25504 44260 25556 44266
rect 25504 44202 25556 44208
rect 25596 44260 25648 44266
rect 25596 44202 25648 44208
rect 25504 43988 25556 43994
rect 25504 43930 25556 43936
rect 25412 43104 25464 43110
rect 25412 43046 25464 43052
rect 25424 41750 25452 43046
rect 25516 42226 25544 43930
rect 25504 42220 25556 42226
rect 25504 42162 25556 42168
rect 25412 41744 25464 41750
rect 25412 41686 25464 41692
rect 25332 41534 25452 41562
rect 25320 41472 25372 41478
rect 25320 41414 25372 41420
rect 25228 41132 25280 41138
rect 25228 41074 25280 41080
rect 25240 39370 25268 41074
rect 25228 39364 25280 39370
rect 25228 39306 25280 39312
rect 25332 38554 25360 41414
rect 25424 41002 25452 41534
rect 25504 41064 25556 41070
rect 25504 41006 25556 41012
rect 25412 40996 25464 41002
rect 25412 40938 25464 40944
rect 25516 40186 25544 41006
rect 25608 40610 25636 44202
rect 25792 42770 25820 44678
rect 26056 44192 26108 44198
rect 26056 44134 26108 44140
rect 25780 42764 25832 42770
rect 25780 42706 25832 42712
rect 25688 42696 25740 42702
rect 25688 42638 25740 42644
rect 25700 40730 25728 42638
rect 26068 42566 26096 44134
rect 26332 43308 26384 43314
rect 26332 43250 26384 43256
rect 26344 42838 26372 43250
rect 26332 42832 26384 42838
rect 26332 42774 26384 42780
rect 26056 42560 26108 42566
rect 26056 42502 26108 42508
rect 25964 42016 26016 42022
rect 25964 41958 26016 41964
rect 25976 41818 26004 41958
rect 25964 41812 26016 41818
rect 25964 41754 26016 41760
rect 25780 41472 25832 41478
rect 25780 41414 25832 41420
rect 25792 41138 25820 41414
rect 25976 41206 26004 41754
rect 25964 41200 26016 41206
rect 25884 41160 25964 41188
rect 25780 41132 25832 41138
rect 25780 41074 25832 41080
rect 25884 40746 25912 41160
rect 25964 41142 26016 41148
rect 25688 40724 25740 40730
rect 25688 40666 25740 40672
rect 25792 40718 25912 40746
rect 25964 40724 26016 40730
rect 25608 40582 25728 40610
rect 25596 40452 25648 40458
rect 25596 40394 25648 40400
rect 25504 40180 25556 40186
rect 25504 40122 25556 40128
rect 25608 40118 25636 40394
rect 25596 40112 25648 40118
rect 25596 40054 25648 40060
rect 25504 40044 25556 40050
rect 25504 39986 25556 39992
rect 25516 39574 25544 39986
rect 25504 39568 25556 39574
rect 25504 39510 25556 39516
rect 25516 39438 25544 39510
rect 25504 39432 25556 39438
rect 25504 39374 25556 39380
rect 25596 39432 25648 39438
rect 25596 39374 25648 39380
rect 25516 39030 25544 39374
rect 25608 39098 25636 39374
rect 25596 39092 25648 39098
rect 25596 39034 25648 39040
rect 25504 39024 25556 39030
rect 25504 38966 25556 38972
rect 25320 38548 25372 38554
rect 25320 38490 25372 38496
rect 25412 38548 25464 38554
rect 25412 38490 25464 38496
rect 25424 38350 25452 38490
rect 25412 38344 25464 38350
rect 25412 38286 25464 38292
rect 25148 38168 25544 38196
rect 25136 37392 25188 37398
rect 25136 37334 25188 37340
rect 25412 37392 25464 37398
rect 25412 37334 25464 37340
rect 25148 36854 25176 37334
rect 25136 36848 25188 36854
rect 25136 36790 25188 36796
rect 25228 36848 25280 36854
rect 25228 36790 25280 36796
rect 25136 36644 25188 36650
rect 25136 36586 25188 36592
rect 25148 35494 25176 36586
rect 25240 36174 25268 36790
rect 25320 36576 25372 36582
rect 25320 36518 25372 36524
rect 25228 36168 25280 36174
rect 25228 36110 25280 36116
rect 25332 36106 25360 36518
rect 25424 36378 25452 37334
rect 25412 36372 25464 36378
rect 25412 36314 25464 36320
rect 25320 36100 25372 36106
rect 25320 36042 25372 36048
rect 25424 36038 25452 36314
rect 25412 36032 25464 36038
rect 25412 35974 25464 35980
rect 25410 35864 25466 35873
rect 25516 35834 25544 38168
rect 25700 38010 25728 40582
rect 25792 40118 25820 40718
rect 25964 40666 26016 40672
rect 25872 40656 25924 40662
rect 25872 40598 25924 40604
rect 25780 40112 25832 40118
rect 25780 40054 25832 40060
rect 25884 39846 25912 40598
rect 25976 40118 26004 40666
rect 25964 40112 26016 40118
rect 25964 40054 26016 40060
rect 26068 39914 26096 42502
rect 26344 40594 26372 42774
rect 26332 40588 26384 40594
rect 26332 40530 26384 40536
rect 26160 40458 26280 40474
rect 26160 40452 26292 40458
rect 26160 40446 26240 40452
rect 26160 40186 26188 40446
rect 26240 40394 26292 40400
rect 26148 40180 26200 40186
rect 26148 40122 26200 40128
rect 26240 40112 26292 40118
rect 26238 40080 26240 40089
rect 26292 40080 26294 40089
rect 26238 40015 26294 40024
rect 26056 39908 26108 39914
rect 26056 39850 26108 39856
rect 25872 39840 25924 39846
rect 25872 39782 25924 39788
rect 26068 39506 26096 39850
rect 26436 39522 26464 46310
rect 26056 39500 26108 39506
rect 26056 39442 26108 39448
rect 26148 39500 26200 39506
rect 26148 39442 26200 39448
rect 26344 39494 26464 39522
rect 25964 38208 26016 38214
rect 25964 38150 26016 38156
rect 25688 38004 25740 38010
rect 25688 37946 25740 37952
rect 25700 37466 25728 37946
rect 25976 37874 26004 38150
rect 25964 37868 26016 37874
rect 25964 37810 26016 37816
rect 26068 37670 26096 39442
rect 26160 39302 26188 39442
rect 26148 39296 26200 39302
rect 26148 39238 26200 39244
rect 26240 38752 26292 38758
rect 26240 38694 26292 38700
rect 26252 38214 26280 38694
rect 26344 38418 26372 39494
rect 26424 39432 26476 39438
rect 26424 39374 26476 39380
rect 26332 38412 26384 38418
rect 26332 38354 26384 38360
rect 26240 38208 26292 38214
rect 26240 38150 26292 38156
rect 25780 37664 25832 37670
rect 25780 37606 25832 37612
rect 26056 37664 26108 37670
rect 26056 37606 26108 37612
rect 25688 37460 25740 37466
rect 25688 37402 25740 37408
rect 25700 36582 25728 37402
rect 25688 36576 25740 36582
rect 25688 36518 25740 36524
rect 25792 36038 25820 37606
rect 26068 37330 26096 37606
rect 26056 37324 26108 37330
rect 26056 37266 26108 37272
rect 25964 37256 26016 37262
rect 25964 37198 26016 37204
rect 25872 36848 25924 36854
rect 25872 36790 25924 36796
rect 25780 36032 25832 36038
rect 25780 35974 25832 35980
rect 25410 35799 25412 35808
rect 25464 35799 25466 35808
rect 25504 35828 25556 35834
rect 25412 35770 25464 35776
rect 25504 35770 25556 35776
rect 25136 35488 25188 35494
rect 25136 35430 25188 35436
rect 25148 35154 25176 35430
rect 25136 35148 25188 35154
rect 25136 35090 25188 35096
rect 25044 34740 25096 34746
rect 25044 34682 25096 34688
rect 25042 34640 25098 34649
rect 24768 34604 24820 34610
rect 25792 34610 25820 35974
rect 25884 35698 25912 36790
rect 25976 36582 26004 37198
rect 26252 36922 26280 38150
rect 26344 37466 26372 38354
rect 26436 37874 26464 39374
rect 26424 37868 26476 37874
rect 26424 37810 26476 37816
rect 26332 37460 26384 37466
rect 26332 37402 26384 37408
rect 26240 36916 26292 36922
rect 26240 36858 26292 36864
rect 26148 36644 26200 36650
rect 26148 36586 26200 36592
rect 25964 36576 26016 36582
rect 25964 36518 26016 36524
rect 25976 35766 26004 36518
rect 26160 36174 26188 36586
rect 26148 36168 26200 36174
rect 26148 36110 26200 36116
rect 26056 36032 26108 36038
rect 26056 35974 26108 35980
rect 25964 35760 26016 35766
rect 25964 35702 26016 35708
rect 25872 35692 25924 35698
rect 25872 35634 25924 35640
rect 25884 35601 25912 35634
rect 26068 35630 26096 35974
rect 26056 35624 26108 35630
rect 25870 35592 25926 35601
rect 26056 35566 26108 35572
rect 25870 35527 25926 35536
rect 26160 35086 26188 36110
rect 26148 35080 26200 35086
rect 26148 35022 26200 35028
rect 26240 35080 26292 35086
rect 26240 35022 26292 35028
rect 25872 35012 25924 35018
rect 25872 34954 25924 34960
rect 25042 34575 25098 34584
rect 25228 34604 25280 34610
rect 24768 34546 24820 34552
rect 25056 34406 25084 34575
rect 25228 34546 25280 34552
rect 25780 34604 25832 34610
rect 25780 34546 25832 34552
rect 25044 34400 25096 34406
rect 25044 34342 25096 34348
rect 25240 34202 25268 34546
rect 25412 34536 25464 34542
rect 25412 34478 25464 34484
rect 25688 34536 25740 34542
rect 25688 34478 25740 34484
rect 25136 34196 25188 34202
rect 25136 34138 25188 34144
rect 25228 34196 25280 34202
rect 25228 34138 25280 34144
rect 24768 33992 24820 33998
rect 24768 33934 24820 33940
rect 24780 33658 24808 33934
rect 24768 33652 24820 33658
rect 24768 33594 24820 33600
rect 24780 33522 25084 33538
rect 24768 33516 25096 33522
rect 24820 33510 25044 33516
rect 24768 33458 24820 33464
rect 25044 33458 25096 33464
rect 25148 33386 25176 34138
rect 25424 33930 25452 34478
rect 25504 34196 25556 34202
rect 25504 34138 25556 34144
rect 25412 33924 25464 33930
rect 25412 33866 25464 33872
rect 25228 33516 25280 33522
rect 25228 33458 25280 33464
rect 24768 33380 24820 33386
rect 24768 33322 24820 33328
rect 25136 33380 25188 33386
rect 25136 33322 25188 33328
rect 24780 32910 24808 33322
rect 24768 32904 24820 32910
rect 24768 32846 24820 32852
rect 24860 32904 24912 32910
rect 24860 32846 24912 32852
rect 24676 32292 24728 32298
rect 24676 32234 24728 32240
rect 24688 31754 24716 32234
rect 24676 31748 24728 31754
rect 24676 31690 24728 31696
rect 24872 31482 24900 32846
rect 24952 32496 25004 32502
rect 24952 32438 25004 32444
rect 24964 31822 24992 32438
rect 25240 32298 25268 33458
rect 25516 32910 25544 34138
rect 25700 33674 25728 34478
rect 25792 34082 25820 34546
rect 25884 34202 25912 34954
rect 26056 34944 26108 34950
rect 26056 34886 26108 34892
rect 26068 34610 26096 34886
rect 26160 34746 26188 35022
rect 26148 34740 26200 34746
rect 26148 34682 26200 34688
rect 26252 34610 26280 35022
rect 26056 34604 26108 34610
rect 26056 34546 26108 34552
rect 26240 34604 26292 34610
rect 26240 34546 26292 34552
rect 25872 34196 25924 34202
rect 25872 34138 25924 34144
rect 25792 34054 26096 34082
rect 25700 33646 25912 33674
rect 25780 33516 25832 33522
rect 25780 33458 25832 33464
rect 25688 33312 25740 33318
rect 25688 33254 25740 33260
rect 25700 32978 25728 33254
rect 25792 33114 25820 33458
rect 25780 33108 25832 33114
rect 25780 33050 25832 33056
rect 25688 32972 25740 32978
rect 25688 32914 25740 32920
rect 25504 32904 25556 32910
rect 25504 32846 25556 32852
rect 25504 32428 25556 32434
rect 25504 32370 25556 32376
rect 25228 32292 25280 32298
rect 25228 32234 25280 32240
rect 25516 32026 25544 32370
rect 25596 32292 25648 32298
rect 25596 32234 25648 32240
rect 25608 32026 25636 32234
rect 25504 32020 25556 32026
rect 25504 31962 25556 31968
rect 25596 32020 25648 32026
rect 25596 31962 25648 31968
rect 24952 31816 25004 31822
rect 24952 31758 25004 31764
rect 24964 31482 24992 31758
rect 24860 31476 24912 31482
rect 24860 31418 24912 31424
rect 24952 31476 25004 31482
rect 24952 31418 25004 31424
rect 24492 30728 24544 30734
rect 24492 30670 24544 30676
rect 24400 30184 24452 30190
rect 24400 30126 24452 30132
rect 24504 29578 24532 30670
rect 24872 30598 24900 31418
rect 25516 31142 25544 31962
rect 25792 31906 25820 33050
rect 25700 31890 25820 31906
rect 25688 31884 25820 31890
rect 25740 31878 25820 31884
rect 25688 31826 25740 31832
rect 25780 31816 25832 31822
rect 25780 31758 25832 31764
rect 25792 31414 25820 31758
rect 25780 31408 25832 31414
rect 25780 31350 25832 31356
rect 25504 31136 25556 31142
rect 25504 31078 25556 31084
rect 24768 30592 24820 30598
rect 24768 30534 24820 30540
rect 24860 30592 24912 30598
rect 24860 30534 24912 30540
rect 24780 30394 24808 30534
rect 24768 30388 24820 30394
rect 24768 30330 24820 30336
rect 24492 29572 24544 29578
rect 24492 29514 24544 29520
rect 24780 29306 24808 30330
rect 24872 29510 24900 30534
rect 25136 30252 25188 30258
rect 25136 30194 25188 30200
rect 25780 30252 25832 30258
rect 25780 30194 25832 30200
rect 25148 29850 25176 30194
rect 25228 30048 25280 30054
rect 25228 29990 25280 29996
rect 25136 29844 25188 29850
rect 25136 29786 25188 29792
rect 25044 29640 25096 29646
rect 25044 29582 25096 29588
rect 24860 29504 24912 29510
rect 24860 29446 24912 29452
rect 24768 29300 24820 29306
rect 24768 29242 24820 29248
rect 24492 29164 24544 29170
rect 24676 29164 24728 29170
rect 24544 29124 24624 29152
rect 24492 29106 24544 29112
rect 23480 28756 23532 28762
rect 23480 28698 23532 28704
rect 24216 28756 24268 28762
rect 24216 28698 24268 28704
rect 23112 28552 23164 28558
rect 23112 28494 23164 28500
rect 23020 28484 23072 28490
rect 23020 28426 23072 28432
rect 23492 28150 23520 28698
rect 24596 28626 24624 29124
rect 24872 29152 24900 29446
rect 24728 29124 24900 29152
rect 24676 29106 24728 29112
rect 24872 28966 24900 29124
rect 24860 28960 24912 28966
rect 24860 28902 24912 28908
rect 24584 28620 24636 28626
rect 24584 28562 24636 28568
rect 23480 28144 23532 28150
rect 23480 28086 23532 28092
rect 23492 28014 23520 28086
rect 23480 28008 23532 28014
rect 23480 27950 23532 27956
rect 23572 27872 23624 27878
rect 23572 27814 23624 27820
rect 23584 27470 23612 27814
rect 22928 27464 22980 27470
rect 22928 27406 22980 27412
rect 23572 27464 23624 27470
rect 23572 27406 23624 27412
rect 22940 26382 22968 27406
rect 23020 27396 23072 27402
rect 23020 27338 23072 27344
rect 23032 26994 23060 27338
rect 24596 27130 24624 28562
rect 24872 28558 24900 28902
rect 25056 28762 25084 29582
rect 25148 29170 25176 29786
rect 25240 29714 25268 29990
rect 25228 29708 25280 29714
rect 25228 29650 25280 29656
rect 25792 29646 25820 30194
rect 25884 29782 25912 33646
rect 25964 32904 26016 32910
rect 25964 32846 26016 32852
rect 25976 32570 26004 32846
rect 25964 32564 26016 32570
rect 25964 32506 26016 32512
rect 26068 31414 26096 34054
rect 26620 32842 26648 46514
rect 26792 45620 26844 45626
rect 26792 45562 26844 45568
rect 26700 42560 26752 42566
rect 26700 42502 26752 42508
rect 26712 39982 26740 42502
rect 26700 39976 26752 39982
rect 26700 39918 26752 39924
rect 26700 39840 26752 39846
rect 26700 39782 26752 39788
rect 26712 38350 26740 39782
rect 26700 38344 26752 38350
rect 26700 38286 26752 38292
rect 26712 37369 26740 38286
rect 26698 37360 26754 37369
rect 26698 37295 26754 37304
rect 26804 36378 26832 45562
rect 26896 41414 26924 47466
rect 27080 46050 27108 49200
rect 28356 47116 28408 47122
rect 28356 47058 28408 47064
rect 28368 46578 28396 47058
rect 28816 46980 28868 46986
rect 28816 46922 28868 46928
rect 28356 46572 28408 46578
rect 28356 46514 28408 46520
rect 27988 46504 28040 46510
rect 27988 46446 28040 46452
rect 27436 46368 27488 46374
rect 27436 46310 27488 46316
rect 27080 46022 27200 46050
rect 27068 45960 27120 45966
rect 27068 45902 27120 45908
rect 26976 45824 27028 45830
rect 26976 45766 27028 45772
rect 26988 45490 27016 45766
rect 26976 45484 27028 45490
rect 26976 45426 27028 45432
rect 26988 43926 27016 45426
rect 27080 44946 27108 45902
rect 27172 45354 27200 46022
rect 27160 45348 27212 45354
rect 27160 45290 27212 45296
rect 27068 44940 27120 44946
rect 27068 44882 27120 44888
rect 26976 43920 27028 43926
rect 26976 43862 27028 43868
rect 27080 43858 27108 44882
rect 27068 43852 27120 43858
rect 27068 43794 27120 43800
rect 26976 43784 27028 43790
rect 26976 43726 27028 43732
rect 26988 43246 27016 43726
rect 27080 43314 27108 43794
rect 27252 43376 27304 43382
rect 27252 43318 27304 43324
rect 27068 43308 27120 43314
rect 27068 43250 27120 43256
rect 26976 43240 27028 43246
rect 26976 43182 27028 43188
rect 27080 42770 27108 43250
rect 27068 42764 27120 42770
rect 27068 42706 27120 42712
rect 27080 41818 27108 42706
rect 27160 42016 27212 42022
rect 27160 41958 27212 41964
rect 27172 41857 27200 41958
rect 27158 41848 27214 41857
rect 27068 41812 27120 41818
rect 27158 41783 27214 41792
rect 27068 41754 27120 41760
rect 27080 41698 27108 41754
rect 27080 41670 27200 41698
rect 26896 41386 27108 41414
rect 27080 41018 27108 41386
rect 26896 40990 27108 41018
rect 26896 36825 26924 40990
rect 27068 40928 27120 40934
rect 27068 40870 27120 40876
rect 27080 40730 27108 40870
rect 27068 40724 27120 40730
rect 27068 40666 27120 40672
rect 27172 40594 27200 41670
rect 27160 40588 27212 40594
rect 27160 40530 27212 40536
rect 27264 40186 27292 43318
rect 27344 41744 27396 41750
rect 27344 41686 27396 41692
rect 27356 41313 27384 41686
rect 27342 41304 27398 41313
rect 27448 41274 27476 46310
rect 27528 44804 27580 44810
rect 27528 44746 27580 44752
rect 27540 41449 27568 44746
rect 27896 44396 27948 44402
rect 27896 44338 27948 44344
rect 27620 43648 27672 43654
rect 27620 43590 27672 43596
rect 27632 43110 27660 43590
rect 27620 43104 27672 43110
rect 27620 43046 27672 43052
rect 27632 41721 27660 43046
rect 27712 41812 27764 41818
rect 27712 41754 27764 41760
rect 27618 41712 27674 41721
rect 27618 41647 27674 41656
rect 27526 41440 27582 41449
rect 27526 41375 27582 41384
rect 27342 41239 27398 41248
rect 27436 41268 27488 41274
rect 27252 40180 27304 40186
rect 27252 40122 27304 40128
rect 27068 40044 27120 40050
rect 27068 39986 27120 39992
rect 27080 39642 27108 39986
rect 27160 39976 27212 39982
rect 27160 39918 27212 39924
rect 27068 39636 27120 39642
rect 27068 39578 27120 39584
rect 27172 39506 27200 39918
rect 27160 39500 27212 39506
rect 27160 39442 27212 39448
rect 27356 39438 27384 41239
rect 27436 41210 27488 41216
rect 27632 40458 27660 41647
rect 27724 41478 27752 41754
rect 27802 41576 27858 41585
rect 27802 41511 27858 41520
rect 27712 41472 27764 41478
rect 27712 41414 27764 41420
rect 27620 40452 27672 40458
rect 27620 40394 27672 40400
rect 27528 40044 27580 40050
rect 27528 39986 27580 39992
rect 27344 39432 27396 39438
rect 27344 39374 27396 39380
rect 27540 38894 27568 39986
rect 27528 38888 27580 38894
rect 27528 38830 27580 38836
rect 27252 38752 27304 38758
rect 27252 38694 27304 38700
rect 27068 38412 27120 38418
rect 27068 38354 27120 38360
rect 27080 37330 27108 38354
rect 27264 38350 27292 38694
rect 27724 38486 27752 41414
rect 27816 41274 27844 41511
rect 27804 41268 27856 41274
rect 27804 41210 27856 41216
rect 27804 38548 27856 38554
rect 27804 38490 27856 38496
rect 27712 38480 27764 38486
rect 27712 38422 27764 38428
rect 27816 38350 27844 38490
rect 27252 38344 27304 38350
rect 27436 38344 27488 38350
rect 27252 38286 27304 38292
rect 27434 38312 27436 38321
rect 27620 38344 27672 38350
rect 27488 38312 27490 38321
rect 27620 38286 27672 38292
rect 27804 38344 27856 38350
rect 27804 38286 27856 38292
rect 27434 38247 27490 38256
rect 27160 37936 27212 37942
rect 27160 37878 27212 37884
rect 27172 37466 27200 37878
rect 27160 37460 27212 37466
rect 27160 37402 27212 37408
rect 27068 37324 27120 37330
rect 27068 37266 27120 37272
rect 26976 37256 27028 37262
rect 26974 37224 26976 37233
rect 27028 37224 27030 37233
rect 26974 37159 27030 37168
rect 26882 36816 26938 36825
rect 26882 36751 26938 36760
rect 27528 36712 27580 36718
rect 27528 36654 27580 36660
rect 27540 36378 27568 36654
rect 27632 36378 27660 38286
rect 27802 37496 27858 37505
rect 27802 37431 27858 37440
rect 27816 37398 27844 37431
rect 27804 37392 27856 37398
rect 27804 37334 27856 37340
rect 27712 37324 27764 37330
rect 27712 37266 27764 37272
rect 26792 36372 26844 36378
rect 26792 36314 26844 36320
rect 27528 36372 27580 36378
rect 27528 36314 27580 36320
rect 27620 36372 27672 36378
rect 27620 36314 27672 36320
rect 26804 35766 26832 36314
rect 27724 36174 27752 37266
rect 27816 36786 27844 37334
rect 27804 36780 27856 36786
rect 27804 36722 27856 36728
rect 27712 36168 27764 36174
rect 27712 36110 27764 36116
rect 26792 35760 26844 35766
rect 26792 35702 26844 35708
rect 27160 35760 27212 35766
rect 27160 35702 27212 35708
rect 26804 35018 26832 35702
rect 26976 35556 27028 35562
rect 26976 35498 27028 35504
rect 26988 35290 27016 35498
rect 27068 35488 27120 35494
rect 27068 35430 27120 35436
rect 26976 35284 27028 35290
rect 26976 35226 27028 35232
rect 26792 35012 26844 35018
rect 26792 34954 26844 34960
rect 26988 33998 27016 35226
rect 27080 35086 27108 35430
rect 27068 35080 27120 35086
rect 27068 35022 27120 35028
rect 27066 34912 27122 34921
rect 27066 34847 27122 34856
rect 27080 34542 27108 34847
rect 27172 34610 27200 35702
rect 27620 35692 27672 35698
rect 27620 35634 27672 35640
rect 27252 35488 27304 35494
rect 27252 35430 27304 35436
rect 27264 35086 27292 35430
rect 27252 35080 27304 35086
rect 27252 35022 27304 35028
rect 27632 35018 27660 35634
rect 27712 35624 27764 35630
rect 27712 35566 27764 35572
rect 27724 35222 27752 35566
rect 27712 35216 27764 35222
rect 27712 35158 27764 35164
rect 27620 35012 27672 35018
rect 27620 34954 27672 34960
rect 27252 34944 27304 34950
rect 27252 34886 27304 34892
rect 27344 34944 27396 34950
rect 27344 34886 27396 34892
rect 27160 34604 27212 34610
rect 27160 34546 27212 34552
rect 27264 34542 27292 34886
rect 27068 34536 27120 34542
rect 27068 34478 27120 34484
rect 27252 34536 27304 34542
rect 27252 34478 27304 34484
rect 26792 33992 26844 33998
rect 26792 33934 26844 33940
rect 26976 33992 27028 33998
rect 26976 33934 27028 33940
rect 26804 33046 26832 33934
rect 26976 33856 27028 33862
rect 26976 33798 27028 33804
rect 26988 33454 27016 33798
rect 26976 33448 27028 33454
rect 26976 33390 27028 33396
rect 27160 33312 27212 33318
rect 27160 33254 27212 33260
rect 26792 33040 26844 33046
rect 26792 32982 26844 32988
rect 26700 32904 26752 32910
rect 27068 32904 27120 32910
rect 26752 32864 27068 32892
rect 26700 32846 26752 32852
rect 27068 32846 27120 32852
rect 26608 32836 26660 32842
rect 26608 32778 26660 32784
rect 26712 31958 26740 32846
rect 27172 32434 27200 33254
rect 26792 32428 26844 32434
rect 26792 32370 26844 32376
rect 27160 32428 27212 32434
rect 27160 32370 27212 32376
rect 26700 31952 26752 31958
rect 26700 31894 26752 31900
rect 26608 31816 26660 31822
rect 26608 31758 26660 31764
rect 26240 31476 26292 31482
rect 26240 31418 26292 31424
rect 26056 31408 26108 31414
rect 26056 31350 26108 31356
rect 26252 31346 26280 31418
rect 26240 31340 26292 31346
rect 26240 31282 26292 31288
rect 25964 30728 26016 30734
rect 25964 30670 26016 30676
rect 25872 29776 25924 29782
rect 25872 29718 25924 29724
rect 25976 29646 26004 30670
rect 26252 30598 26280 31282
rect 26240 30592 26292 30598
rect 26240 30534 26292 30540
rect 26516 30592 26568 30598
rect 26516 30534 26568 30540
rect 26240 30048 26292 30054
rect 26240 29990 26292 29996
rect 25780 29640 25832 29646
rect 25780 29582 25832 29588
rect 25964 29640 26016 29646
rect 25964 29582 26016 29588
rect 25688 29504 25740 29510
rect 25688 29446 25740 29452
rect 25700 29170 25728 29446
rect 25136 29164 25188 29170
rect 25136 29106 25188 29112
rect 25688 29164 25740 29170
rect 25688 29106 25740 29112
rect 25700 28966 25728 29106
rect 25688 28960 25740 28966
rect 25688 28902 25740 28908
rect 25044 28756 25096 28762
rect 25044 28698 25096 28704
rect 24860 28552 24912 28558
rect 24860 28494 24912 28500
rect 24768 28076 24820 28082
rect 24768 28018 24820 28024
rect 24780 27470 24808 28018
rect 24872 27946 24900 28494
rect 26056 28144 26108 28150
rect 26056 28086 26108 28092
rect 25964 28076 26016 28082
rect 25964 28018 26016 28024
rect 25228 28008 25280 28014
rect 25228 27950 25280 27956
rect 24860 27940 24912 27946
rect 24860 27882 24912 27888
rect 24952 27872 25004 27878
rect 24952 27814 25004 27820
rect 24964 27606 24992 27814
rect 24952 27600 25004 27606
rect 24952 27542 25004 27548
rect 24768 27464 24820 27470
rect 24964 27418 24992 27542
rect 24768 27406 24820 27412
rect 24780 27130 24808 27406
rect 24872 27390 24992 27418
rect 25136 27464 25188 27470
rect 25136 27406 25188 27412
rect 24584 27124 24636 27130
rect 24584 27066 24636 27072
rect 24768 27124 24820 27130
rect 24768 27066 24820 27072
rect 24780 26994 24808 27066
rect 23020 26988 23072 26994
rect 23020 26930 23072 26936
rect 24032 26988 24084 26994
rect 24032 26930 24084 26936
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 23112 26920 23164 26926
rect 23112 26862 23164 26868
rect 23124 26586 23152 26862
rect 23112 26580 23164 26586
rect 23112 26522 23164 26528
rect 24044 26518 24072 26930
rect 24872 26874 24900 27390
rect 24952 27328 25004 27334
rect 24952 27270 25004 27276
rect 24964 26994 24992 27270
rect 24952 26988 25004 26994
rect 24952 26930 25004 26936
rect 25044 26988 25096 26994
rect 25044 26930 25096 26936
rect 24872 26858 24992 26874
rect 24872 26852 25004 26858
rect 24872 26846 24952 26852
rect 24952 26794 25004 26800
rect 24860 26784 24912 26790
rect 24860 26726 24912 26732
rect 24032 26512 24084 26518
rect 24032 26454 24084 26460
rect 22928 26376 22980 26382
rect 22928 26318 22980 26324
rect 24584 25900 24636 25906
rect 24584 25842 24636 25848
rect 24768 25900 24820 25906
rect 24768 25842 24820 25848
rect 23756 25152 23808 25158
rect 23756 25094 23808 25100
rect 23768 24818 23796 25094
rect 24596 24818 24624 25842
rect 23756 24812 23808 24818
rect 23756 24754 23808 24760
rect 23940 24812 23992 24818
rect 23940 24754 23992 24760
rect 24584 24812 24636 24818
rect 24584 24754 24636 24760
rect 23204 24744 23256 24750
rect 23204 24686 23256 24692
rect 22572 22066 22692 22094
rect 22468 5568 22520 5574
rect 22468 5510 22520 5516
rect 20904 2644 20956 2650
rect 20904 2586 20956 2592
rect 22572 2582 22600 22066
rect 23216 2650 23244 24686
rect 23768 24206 23796 24754
rect 23952 24274 23980 24754
rect 24596 24410 24624 24754
rect 24780 24750 24808 25842
rect 24872 25786 24900 26726
rect 25056 26586 25084 26930
rect 25044 26580 25096 26586
rect 25044 26522 25096 26528
rect 25148 26382 25176 27406
rect 25240 27062 25268 27950
rect 25504 27940 25556 27946
rect 25504 27882 25556 27888
rect 25228 27056 25280 27062
rect 25228 26998 25280 27004
rect 25136 26376 25188 26382
rect 25136 26318 25188 26324
rect 24872 25758 24992 25786
rect 24860 25696 24912 25702
rect 24860 25638 24912 25644
rect 24872 25294 24900 25638
rect 24964 25362 24992 25758
rect 24952 25356 25004 25362
rect 24952 25298 25004 25304
rect 24860 25288 24912 25294
rect 24860 25230 24912 25236
rect 24964 25242 24992 25298
rect 24964 25214 25084 25242
rect 25056 24818 25084 25214
rect 25044 24812 25096 24818
rect 25044 24754 25096 24760
rect 24768 24744 24820 24750
rect 24768 24686 24820 24692
rect 24584 24404 24636 24410
rect 24584 24346 24636 24352
rect 23940 24268 23992 24274
rect 23940 24210 23992 24216
rect 23756 24200 23808 24206
rect 23756 24142 23808 24148
rect 23768 24070 23796 24142
rect 23756 24064 23808 24070
rect 23756 24006 23808 24012
rect 23204 2644 23256 2650
rect 23204 2586 23256 2592
rect 22560 2576 22612 2582
rect 22560 2518 22612 2524
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 22560 2440 22612 2446
rect 22560 2382 22612 2388
rect 20732 2292 20760 2382
rect 20640 2264 20760 2292
rect 20352 1828 20404 1834
rect 20352 1770 20404 1776
rect 20640 800 20668 2264
rect 22572 800 22600 2382
rect 23768 2378 23796 24006
rect 24492 2848 24544 2854
rect 24492 2790 24544 2796
rect 24504 2378 24532 2790
rect 25516 2582 25544 27882
rect 25976 27334 26004 28018
rect 26068 27674 26096 28086
rect 26056 27668 26108 27674
rect 26056 27610 26108 27616
rect 26252 27470 26280 29990
rect 26424 29708 26476 29714
rect 26424 29650 26476 29656
rect 26332 29096 26384 29102
rect 26332 29038 26384 29044
rect 26344 28762 26372 29038
rect 26332 28756 26384 28762
rect 26332 28698 26384 28704
rect 26332 28552 26384 28558
rect 26436 28540 26464 29650
rect 26528 28966 26556 30534
rect 26516 28960 26568 28966
rect 26516 28902 26568 28908
rect 26384 28512 26464 28540
rect 26332 28494 26384 28500
rect 26240 27464 26292 27470
rect 26240 27406 26292 27412
rect 25964 27328 26016 27334
rect 25964 27270 26016 27276
rect 25976 27130 26004 27270
rect 25964 27124 26016 27130
rect 25964 27066 26016 27072
rect 26252 26382 26280 27406
rect 26344 27130 26372 28494
rect 26528 28082 26556 28902
rect 26516 28076 26568 28082
rect 26516 28018 26568 28024
rect 26528 27402 26556 28018
rect 26516 27396 26568 27402
rect 26516 27338 26568 27344
rect 26332 27124 26384 27130
rect 26332 27066 26384 27072
rect 26528 26586 26556 27338
rect 26516 26580 26568 26586
rect 26516 26522 26568 26528
rect 25780 26376 25832 26382
rect 25780 26318 25832 26324
rect 26240 26376 26292 26382
rect 26240 26318 26292 26324
rect 25792 25430 25820 26318
rect 26148 25832 26200 25838
rect 26148 25774 26200 25780
rect 26160 25430 26188 25774
rect 26252 25702 26280 26318
rect 26240 25696 26292 25702
rect 26240 25638 26292 25644
rect 25780 25424 25832 25430
rect 25780 25366 25832 25372
rect 26148 25424 26200 25430
rect 26148 25366 26200 25372
rect 26160 24954 26188 25366
rect 26148 24948 26200 24954
rect 26148 24890 26200 24896
rect 26252 2650 26280 25638
rect 26620 24410 26648 31758
rect 26804 31754 26832 32370
rect 27172 31906 27200 32370
rect 27080 31878 27200 31906
rect 27080 31822 27108 31878
rect 27068 31816 27120 31822
rect 27068 31758 27120 31764
rect 26792 31748 26844 31754
rect 26792 31690 26844 31696
rect 27264 31482 27292 34478
rect 27356 33522 27384 34886
rect 27632 34678 27660 34954
rect 27620 34672 27672 34678
rect 27620 34614 27672 34620
rect 27620 34536 27672 34542
rect 27620 34478 27672 34484
rect 27632 34202 27660 34478
rect 27620 34196 27672 34202
rect 27620 34138 27672 34144
rect 27724 34082 27752 35158
rect 27528 34060 27580 34066
rect 27528 34002 27580 34008
rect 27632 34054 27752 34082
rect 27344 33516 27396 33522
rect 27344 33458 27396 33464
rect 27436 33516 27488 33522
rect 27436 33458 27488 33464
rect 27252 31476 27304 31482
rect 27252 31418 27304 31424
rect 27068 31340 27120 31346
rect 27068 31282 27120 31288
rect 27080 31142 27108 31282
rect 27068 31136 27120 31142
rect 27068 31078 27120 31084
rect 26792 30728 26844 30734
rect 26792 30670 26844 30676
rect 26804 30122 26832 30670
rect 26976 30592 27028 30598
rect 26976 30534 27028 30540
rect 26884 30252 26936 30258
rect 26884 30194 26936 30200
rect 26792 30116 26844 30122
rect 26792 30058 26844 30064
rect 26804 29850 26832 30058
rect 26792 29844 26844 29850
rect 26792 29786 26844 29792
rect 26896 29646 26924 30194
rect 26884 29640 26936 29646
rect 26884 29582 26936 29588
rect 26792 28484 26844 28490
rect 26792 28426 26844 28432
rect 26804 27946 26832 28426
rect 26896 28422 26924 29582
rect 26988 29170 27016 30534
rect 27080 30054 27108 31078
rect 27264 30870 27292 31418
rect 27252 30864 27304 30870
rect 27252 30806 27304 30812
rect 27448 30326 27476 33458
rect 27540 33114 27568 34002
rect 27632 33862 27660 34054
rect 27712 33924 27764 33930
rect 27712 33866 27764 33872
rect 27620 33856 27672 33862
rect 27620 33798 27672 33804
rect 27620 33652 27672 33658
rect 27620 33594 27672 33600
rect 27528 33108 27580 33114
rect 27528 33050 27580 33056
rect 27632 32994 27660 33594
rect 27724 33522 27752 33866
rect 27712 33516 27764 33522
rect 27712 33458 27764 33464
rect 27540 32966 27660 32994
rect 27540 32502 27568 32966
rect 27816 32858 27844 36722
rect 27908 35873 27936 44338
rect 28000 38554 28028 46446
rect 28632 46028 28684 46034
rect 28632 45970 28684 45976
rect 28540 45824 28592 45830
rect 28540 45766 28592 45772
rect 28356 45280 28408 45286
rect 28356 45222 28408 45228
rect 28080 44736 28132 44742
rect 28080 44678 28132 44684
rect 28092 43450 28120 44678
rect 28368 44577 28396 45222
rect 28354 44568 28410 44577
rect 28354 44503 28410 44512
rect 28080 43444 28132 43450
rect 28080 43386 28132 43392
rect 28092 41818 28120 43386
rect 28080 41812 28132 41818
rect 28080 41754 28132 41760
rect 28356 39840 28408 39846
rect 28408 39800 28488 39828
rect 28356 39782 28408 39788
rect 28080 39432 28132 39438
rect 28080 39374 28132 39380
rect 28356 39432 28408 39438
rect 28356 39374 28408 39380
rect 27988 38548 28040 38554
rect 27988 38490 28040 38496
rect 27988 37256 28040 37262
rect 27988 37198 28040 37204
rect 28000 36174 28028 37198
rect 27988 36168 28040 36174
rect 27988 36110 28040 36116
rect 27894 35864 27950 35873
rect 27894 35799 27950 35808
rect 27894 34912 27950 34921
rect 27894 34847 27950 34856
rect 27908 33658 27936 34847
rect 27988 34128 28040 34134
rect 27988 34070 28040 34076
rect 27896 33652 27948 33658
rect 27896 33594 27948 33600
rect 27724 32830 27844 32858
rect 27896 32836 27948 32842
rect 27620 32768 27672 32774
rect 27620 32710 27672 32716
rect 27528 32496 27580 32502
rect 27528 32438 27580 32444
rect 27632 32434 27660 32710
rect 27620 32428 27672 32434
rect 27620 32370 27672 32376
rect 27620 31816 27672 31822
rect 27620 31758 27672 31764
rect 27632 31482 27660 31758
rect 27724 31754 27752 32830
rect 27896 32778 27948 32784
rect 27804 32768 27856 32774
rect 27804 32710 27856 32716
rect 27816 32570 27844 32710
rect 27804 32564 27856 32570
rect 27804 32506 27856 32512
rect 27816 32366 27844 32506
rect 27804 32360 27856 32366
rect 27804 32302 27856 32308
rect 27908 32314 27936 32778
rect 28000 32502 28028 34070
rect 27988 32496 28040 32502
rect 27988 32438 28040 32444
rect 27816 31958 27844 32302
rect 27908 32286 28028 32314
rect 27896 32224 27948 32230
rect 27896 32166 27948 32172
rect 27804 31952 27856 31958
rect 27804 31894 27856 31900
rect 27908 31822 27936 32166
rect 27896 31816 27948 31822
rect 27896 31758 27948 31764
rect 27724 31726 27844 31754
rect 27712 31680 27764 31686
rect 27712 31622 27764 31628
rect 27528 31476 27580 31482
rect 27528 31418 27580 31424
rect 27620 31476 27672 31482
rect 27620 31418 27672 31424
rect 27540 30666 27568 31418
rect 27724 30938 27752 31622
rect 27712 30932 27764 30938
rect 27712 30874 27764 30880
rect 27528 30660 27580 30666
rect 27528 30602 27580 30608
rect 27436 30320 27488 30326
rect 27436 30262 27488 30268
rect 27068 30048 27120 30054
rect 27068 29990 27120 29996
rect 27540 29714 27568 30602
rect 27816 30054 27844 31726
rect 28000 31482 28028 32286
rect 28092 32026 28120 39374
rect 28368 39098 28396 39374
rect 28460 39098 28488 39800
rect 28356 39092 28408 39098
rect 28356 39034 28408 39040
rect 28448 39092 28500 39098
rect 28448 39034 28500 39040
rect 28460 38978 28488 39034
rect 28264 38956 28316 38962
rect 28264 38898 28316 38904
rect 28368 38950 28488 38978
rect 28172 38820 28224 38826
rect 28172 38762 28224 38768
rect 28184 37466 28212 38762
rect 28172 37460 28224 37466
rect 28172 37402 28224 37408
rect 28184 36802 28212 37402
rect 28276 36922 28304 38898
rect 28368 37874 28396 38950
rect 28448 38888 28500 38894
rect 28448 38830 28500 38836
rect 28460 38486 28488 38830
rect 28448 38480 28500 38486
rect 28448 38422 28500 38428
rect 28460 38282 28488 38422
rect 28448 38276 28500 38282
rect 28448 38218 28500 38224
rect 28356 37868 28408 37874
rect 28356 37810 28408 37816
rect 28448 37800 28500 37806
rect 28446 37768 28448 37777
rect 28500 37768 28502 37777
rect 28356 37732 28408 37738
rect 28446 37703 28502 37712
rect 28356 37674 28408 37680
rect 28368 37398 28396 37674
rect 28448 37664 28500 37670
rect 28448 37606 28500 37612
rect 28356 37392 28408 37398
rect 28356 37334 28408 37340
rect 28460 37262 28488 37606
rect 28552 37466 28580 45766
rect 28644 45626 28672 45970
rect 28632 45620 28684 45626
rect 28632 45562 28684 45568
rect 28724 43648 28776 43654
rect 28724 43590 28776 43596
rect 28632 42560 28684 42566
rect 28632 42502 28684 42508
rect 28644 41721 28672 42502
rect 28630 41712 28686 41721
rect 28630 41647 28686 41656
rect 28632 38956 28684 38962
rect 28632 38898 28684 38904
rect 28644 38350 28672 38898
rect 28736 38468 28764 43590
rect 28828 39642 28856 46922
rect 29012 45626 29040 49200
rect 30840 47796 30892 47802
rect 30840 47738 30892 47744
rect 29828 47728 29880 47734
rect 29828 47670 29880 47676
rect 29840 47054 29868 47670
rect 30852 47190 30880 47738
rect 30840 47184 30892 47190
rect 30840 47126 30892 47132
rect 29828 47048 29880 47054
rect 30852 47025 30880 47126
rect 29828 46990 29880 46996
rect 30838 47016 30894 47025
rect 29184 46980 29236 46986
rect 30838 46951 30894 46960
rect 29184 46922 29236 46928
rect 29092 45960 29144 45966
rect 29092 45902 29144 45908
rect 29000 45620 29052 45626
rect 29000 45562 29052 45568
rect 29104 44520 29132 45902
rect 29012 44492 29132 44520
rect 29012 44334 29040 44492
rect 29000 44328 29052 44334
rect 29000 44270 29052 44276
rect 29000 44192 29052 44198
rect 29052 44152 29132 44180
rect 29000 44134 29052 44140
rect 29000 43444 29052 43450
rect 29000 43386 29052 43392
rect 28908 42560 28960 42566
rect 28908 42502 28960 42508
rect 28920 41993 28948 42502
rect 28906 41984 28962 41993
rect 28906 41919 28962 41928
rect 29012 41614 29040 43386
rect 29104 42226 29132 44152
rect 29196 43722 29224 46922
rect 30944 46578 30972 49200
rect 32496 47660 32548 47666
rect 32496 47602 32548 47608
rect 32128 47048 32180 47054
rect 32128 46990 32180 46996
rect 31944 46980 31996 46986
rect 31944 46922 31996 46928
rect 30932 46572 30984 46578
rect 30932 46514 30984 46520
rect 31484 46572 31536 46578
rect 31484 46514 31536 46520
rect 29642 46472 29698 46481
rect 29642 46407 29698 46416
rect 31024 46436 31076 46442
rect 29656 45490 29684 46407
rect 31024 46378 31076 46384
rect 31036 46102 31064 46378
rect 31300 46368 31352 46374
rect 31300 46310 31352 46316
rect 31024 46096 31076 46102
rect 31024 46038 31076 46044
rect 30288 45960 30340 45966
rect 30288 45902 30340 45908
rect 30012 45824 30064 45830
rect 30012 45766 30064 45772
rect 29644 45484 29696 45490
rect 29644 45426 29696 45432
rect 29276 44804 29328 44810
rect 29276 44746 29328 44752
rect 29184 43716 29236 43722
rect 29184 43658 29236 43664
rect 29196 43450 29224 43658
rect 29184 43444 29236 43450
rect 29184 43386 29236 43392
rect 29288 43058 29316 44746
rect 29368 43784 29420 43790
rect 29368 43726 29420 43732
rect 29196 43030 29316 43058
rect 29092 42220 29144 42226
rect 29092 42162 29144 42168
rect 29104 41682 29132 42162
rect 29092 41676 29144 41682
rect 29092 41618 29144 41624
rect 29000 41608 29052 41614
rect 29000 41550 29052 41556
rect 28908 41472 28960 41478
rect 28908 41414 28960 41420
rect 28920 41313 28948 41414
rect 28906 41304 28962 41313
rect 28906 41239 28962 41248
rect 28920 40497 28948 41239
rect 29012 41206 29040 41550
rect 29104 41274 29132 41618
rect 29092 41268 29144 41274
rect 29092 41210 29144 41216
rect 29000 41200 29052 41206
rect 29000 41142 29052 41148
rect 29104 41138 29132 41210
rect 29092 41132 29144 41138
rect 29092 41074 29144 41080
rect 29000 40996 29052 41002
rect 29000 40938 29052 40944
rect 28906 40488 28962 40497
rect 28906 40423 28962 40432
rect 28816 39636 28868 39642
rect 28816 39578 28868 39584
rect 29012 39438 29040 40938
rect 29104 40594 29132 41074
rect 29092 40588 29144 40594
rect 29092 40530 29144 40536
rect 29000 39432 29052 39438
rect 29000 39374 29052 39380
rect 29092 39364 29144 39370
rect 29092 39306 29144 39312
rect 28816 38956 28868 38962
rect 28868 38916 28948 38944
rect 28816 38898 28868 38904
rect 28736 38440 28856 38468
rect 28632 38344 28684 38350
rect 28632 38286 28684 38292
rect 28632 37868 28684 37874
rect 28632 37810 28684 37816
rect 28644 37505 28672 37810
rect 28630 37496 28686 37505
rect 28540 37460 28592 37466
rect 28630 37431 28686 37440
rect 28540 37402 28592 37408
rect 28448 37256 28500 37262
rect 28448 37198 28500 37204
rect 28632 37256 28684 37262
rect 28632 37198 28684 37204
rect 28724 37256 28776 37262
rect 28724 37198 28776 37204
rect 28540 37120 28592 37126
rect 28540 37062 28592 37068
rect 28264 36916 28316 36922
rect 28264 36858 28316 36864
rect 28184 36774 28304 36802
rect 28552 36786 28580 37062
rect 28644 36922 28672 37198
rect 28632 36916 28684 36922
rect 28632 36858 28684 36864
rect 28736 36786 28764 37198
rect 28172 36576 28224 36582
rect 28172 36518 28224 36524
rect 28184 36174 28212 36518
rect 28172 36168 28224 36174
rect 28172 36110 28224 36116
rect 28276 35290 28304 36774
rect 28448 36780 28500 36786
rect 28448 36722 28500 36728
rect 28540 36780 28592 36786
rect 28540 36722 28592 36728
rect 28724 36780 28776 36786
rect 28724 36722 28776 36728
rect 28460 36650 28488 36722
rect 28448 36644 28500 36650
rect 28448 36586 28500 36592
rect 28460 36242 28488 36586
rect 28632 36304 28684 36310
rect 28632 36246 28684 36252
rect 28448 36236 28500 36242
rect 28448 36178 28500 36184
rect 28172 35284 28224 35290
rect 28172 35226 28224 35232
rect 28264 35284 28316 35290
rect 28264 35226 28316 35232
rect 28184 34921 28212 35226
rect 28276 35086 28304 35226
rect 28264 35080 28316 35086
rect 28264 35022 28316 35028
rect 28264 34944 28316 34950
rect 28170 34912 28226 34921
rect 28264 34886 28316 34892
rect 28170 34847 28226 34856
rect 28276 34678 28304 34886
rect 28264 34672 28316 34678
rect 28264 34614 28316 34620
rect 28172 34604 28224 34610
rect 28172 34546 28224 34552
rect 28080 32020 28132 32026
rect 28080 31962 28132 31968
rect 27988 31476 28040 31482
rect 27988 31418 28040 31424
rect 27896 31340 27948 31346
rect 27896 31282 27948 31288
rect 27908 30666 27936 31282
rect 28184 31278 28212 34546
rect 28276 33998 28304 34614
rect 28356 34468 28408 34474
rect 28356 34410 28408 34416
rect 28264 33992 28316 33998
rect 28264 33934 28316 33940
rect 28368 33658 28396 34410
rect 28448 34400 28500 34406
rect 28448 34342 28500 34348
rect 28460 33998 28488 34342
rect 28448 33992 28500 33998
rect 28448 33934 28500 33940
rect 28540 33856 28592 33862
rect 28540 33798 28592 33804
rect 28356 33652 28408 33658
rect 28356 33594 28408 33600
rect 28368 32994 28396 33594
rect 28448 33108 28500 33114
rect 28448 33050 28500 33056
rect 28276 32966 28396 32994
rect 28276 32366 28304 32966
rect 28356 32904 28408 32910
rect 28356 32846 28408 32852
rect 28264 32360 28316 32366
rect 28264 32302 28316 32308
rect 28368 32298 28396 32846
rect 28356 32292 28408 32298
rect 28356 32234 28408 32240
rect 28368 32026 28396 32234
rect 28356 32020 28408 32026
rect 28356 31962 28408 31968
rect 28368 31890 28396 31962
rect 28264 31884 28316 31890
rect 28264 31826 28316 31832
rect 28356 31884 28408 31890
rect 28356 31826 28408 31832
rect 28276 31346 28304 31826
rect 28368 31346 28396 31826
rect 28460 31804 28488 33050
rect 28552 32570 28580 33798
rect 28540 32564 28592 32570
rect 28540 32506 28592 32512
rect 28644 32298 28672 36246
rect 28736 36174 28764 36722
rect 28724 36168 28776 36174
rect 28724 36110 28776 36116
rect 28828 35562 28856 38440
rect 28920 36310 28948 38916
rect 29104 38826 29132 39306
rect 29092 38820 29144 38826
rect 29092 38762 29144 38768
rect 29000 38412 29052 38418
rect 29000 38354 29052 38360
rect 29012 37942 29040 38354
rect 29000 37936 29052 37942
rect 29000 37878 29052 37884
rect 29000 36576 29052 36582
rect 29000 36518 29052 36524
rect 28908 36304 28960 36310
rect 28908 36246 28960 36252
rect 28816 35556 28868 35562
rect 28816 35498 28868 35504
rect 29012 35442 29040 36518
rect 29104 35698 29132 38762
rect 29196 38593 29224 43030
rect 29276 42152 29328 42158
rect 29276 42094 29328 42100
rect 29182 38584 29238 38593
rect 29182 38519 29238 38528
rect 29092 35692 29144 35698
rect 29092 35634 29144 35640
rect 28736 35414 29040 35442
rect 28736 34610 28764 35414
rect 28908 34944 28960 34950
rect 28908 34886 28960 34892
rect 28920 34610 28948 34886
rect 28724 34604 28776 34610
rect 28724 34546 28776 34552
rect 28908 34604 28960 34610
rect 28908 34546 28960 34552
rect 28816 34536 28868 34542
rect 28816 34478 28868 34484
rect 28724 34468 28776 34474
rect 28724 34410 28776 34416
rect 28632 32292 28684 32298
rect 28632 32234 28684 32240
rect 28540 31816 28592 31822
rect 28460 31776 28540 31804
rect 28540 31758 28592 31764
rect 28264 31340 28316 31346
rect 28264 31282 28316 31288
rect 28356 31340 28408 31346
rect 28356 31282 28408 31288
rect 28172 31272 28224 31278
rect 28172 31214 28224 31220
rect 28540 31272 28592 31278
rect 28540 31214 28592 31220
rect 27896 30660 27948 30666
rect 27896 30602 27948 30608
rect 27620 30048 27672 30054
rect 27620 29990 27672 29996
rect 27804 30048 27856 30054
rect 27804 29990 27856 29996
rect 27632 29714 27660 29990
rect 27908 29850 27936 30602
rect 28552 30258 28580 31214
rect 28356 30252 28408 30258
rect 28356 30194 28408 30200
rect 28540 30252 28592 30258
rect 28540 30194 28592 30200
rect 27896 29844 27948 29850
rect 27896 29786 27948 29792
rect 27528 29708 27580 29714
rect 27528 29650 27580 29656
rect 27620 29708 27672 29714
rect 27620 29650 27672 29656
rect 27160 29640 27212 29646
rect 27160 29582 27212 29588
rect 26976 29164 27028 29170
rect 26976 29106 27028 29112
rect 27172 28558 27200 29582
rect 27632 29306 27660 29650
rect 28368 29646 28396 30194
rect 28356 29640 28408 29646
rect 28356 29582 28408 29588
rect 28264 29504 28316 29510
rect 28264 29446 28316 29452
rect 28276 29306 28304 29446
rect 28736 29306 28764 34410
rect 28828 33130 28856 34478
rect 29288 34202 29316 42094
rect 29380 39914 29408 43726
rect 29828 42696 29880 42702
rect 29828 42638 29880 42644
rect 29368 39908 29420 39914
rect 29368 39850 29420 39856
rect 29840 39642 29868 42638
rect 29920 41608 29972 41614
rect 29920 41550 29972 41556
rect 29828 39636 29880 39642
rect 29828 39578 29880 39584
rect 29736 38956 29788 38962
rect 29736 38898 29788 38904
rect 29644 38888 29696 38894
rect 29644 38830 29696 38836
rect 29460 38820 29512 38826
rect 29460 38762 29512 38768
rect 29472 35630 29500 38762
rect 29656 38554 29684 38830
rect 29644 38548 29696 38554
rect 29644 38490 29696 38496
rect 29748 38434 29776 38898
rect 29564 38406 29776 38434
rect 29564 38214 29592 38406
rect 29748 38350 29776 38406
rect 29644 38344 29696 38350
rect 29644 38286 29696 38292
rect 29736 38344 29788 38350
rect 29736 38286 29788 38292
rect 29552 38208 29604 38214
rect 29552 38150 29604 38156
rect 29552 37868 29604 37874
rect 29552 37810 29604 37816
rect 29564 36786 29592 37810
rect 29552 36780 29604 36786
rect 29552 36722 29604 36728
rect 29564 36689 29592 36722
rect 29550 36680 29606 36689
rect 29656 36650 29684 38286
rect 29736 38208 29788 38214
rect 29736 38150 29788 38156
rect 29748 37194 29776 38150
rect 29932 38010 29960 41550
rect 29920 38004 29972 38010
rect 29920 37946 29972 37952
rect 30024 37806 30052 45766
rect 30300 45665 30328 45902
rect 30286 45656 30342 45665
rect 30286 45591 30342 45600
rect 30380 45620 30432 45626
rect 30380 45562 30432 45568
rect 30392 43382 30420 45562
rect 31024 45416 31076 45422
rect 31024 45358 31076 45364
rect 31036 45082 31064 45358
rect 30932 45076 30984 45082
rect 30932 45018 30984 45024
rect 31024 45076 31076 45082
rect 31024 45018 31076 45024
rect 30656 44872 30708 44878
rect 30656 44814 30708 44820
rect 30472 44192 30524 44198
rect 30472 44134 30524 44140
rect 30380 43376 30432 43382
rect 30484 43353 30512 44134
rect 30564 43648 30616 43654
rect 30564 43590 30616 43596
rect 30380 43318 30432 43324
rect 30470 43344 30526 43353
rect 30470 43279 30526 43288
rect 30472 42356 30524 42362
rect 30472 42298 30524 42304
rect 30380 42016 30432 42022
rect 30380 41958 30432 41964
rect 30392 41721 30420 41958
rect 30378 41712 30434 41721
rect 30378 41647 30434 41656
rect 30196 41608 30248 41614
rect 30196 41550 30248 41556
rect 30104 40044 30156 40050
rect 30104 39986 30156 39992
rect 30116 38010 30144 39986
rect 30208 39982 30236 41550
rect 30484 41478 30512 42298
rect 30472 41472 30524 41478
rect 30472 41414 30524 41420
rect 30576 40934 30604 43590
rect 30668 42362 30696 44814
rect 30840 43104 30892 43110
rect 30840 43046 30892 43052
rect 30656 42356 30708 42362
rect 30656 42298 30708 42304
rect 30656 42220 30708 42226
rect 30656 42162 30708 42168
rect 30564 40928 30616 40934
rect 30564 40870 30616 40876
rect 30288 40044 30340 40050
rect 30288 39986 30340 39992
rect 30380 40044 30432 40050
rect 30380 39986 30432 39992
rect 30472 40044 30524 40050
rect 30472 39986 30524 39992
rect 30196 39976 30248 39982
rect 30196 39918 30248 39924
rect 30196 39840 30248 39846
rect 30196 39782 30248 39788
rect 30208 38350 30236 39782
rect 30196 38344 30248 38350
rect 30196 38286 30248 38292
rect 30300 38010 30328 39986
rect 30392 38554 30420 39986
rect 30484 39914 30512 39986
rect 30472 39908 30524 39914
rect 30472 39850 30524 39856
rect 30576 39438 30604 40870
rect 30564 39432 30616 39438
rect 30564 39374 30616 39380
rect 30472 39296 30524 39302
rect 30472 39238 30524 39244
rect 30380 38548 30432 38554
rect 30380 38490 30432 38496
rect 30104 38004 30156 38010
rect 30104 37946 30156 37952
rect 30288 38004 30340 38010
rect 30288 37946 30340 37952
rect 30288 37868 30340 37874
rect 30288 37810 30340 37816
rect 30012 37800 30064 37806
rect 30300 37777 30328 37810
rect 30012 37742 30064 37748
rect 30286 37768 30342 37777
rect 30196 37732 30248 37738
rect 30286 37703 30342 37712
rect 30196 37674 30248 37680
rect 30208 37398 30236 37674
rect 30196 37392 30248 37398
rect 30196 37334 30248 37340
rect 30104 37324 30156 37330
rect 30104 37266 30156 37272
rect 30116 37233 30144 37266
rect 30102 37224 30158 37233
rect 29736 37188 29788 37194
rect 30102 37159 30158 37168
rect 29736 37130 29788 37136
rect 29828 37120 29880 37126
rect 29828 37062 29880 37068
rect 29840 36854 29868 37062
rect 29828 36848 29880 36854
rect 29828 36790 29880 36796
rect 30116 36786 30144 37159
rect 30104 36780 30156 36786
rect 30104 36722 30156 36728
rect 29550 36615 29606 36624
rect 29644 36644 29696 36650
rect 29644 36586 29696 36592
rect 30102 36544 30158 36553
rect 30102 36479 30158 36488
rect 30012 35828 30064 35834
rect 30012 35770 30064 35776
rect 29460 35624 29512 35630
rect 29460 35566 29512 35572
rect 29828 35624 29880 35630
rect 29828 35566 29880 35572
rect 29552 35488 29604 35494
rect 29552 35430 29604 35436
rect 29564 34202 29592 35430
rect 29276 34196 29328 34202
rect 29276 34138 29328 34144
rect 29552 34196 29604 34202
rect 29552 34138 29604 34144
rect 29184 33516 29236 33522
rect 29184 33458 29236 33464
rect 28828 33102 28948 33130
rect 28816 32768 28868 32774
rect 28816 32710 28868 32716
rect 28828 32434 28856 32710
rect 28816 32428 28868 32434
rect 28816 32370 28868 32376
rect 28816 30320 28868 30326
rect 28816 30262 28868 30268
rect 28828 30054 28856 30262
rect 28816 30048 28868 30054
rect 28816 29990 28868 29996
rect 28920 29850 28948 33102
rect 29000 32224 29052 32230
rect 29000 32166 29052 32172
rect 29012 32026 29040 32166
rect 29000 32020 29052 32026
rect 29000 31962 29052 31968
rect 29000 31748 29052 31754
rect 29000 31690 29052 31696
rect 29012 31482 29040 31690
rect 29000 31476 29052 31482
rect 29000 31418 29052 31424
rect 29092 31408 29144 31414
rect 29092 31350 29144 31356
rect 29000 30592 29052 30598
rect 29000 30534 29052 30540
rect 28908 29844 28960 29850
rect 28908 29786 28960 29792
rect 27620 29300 27672 29306
rect 27620 29242 27672 29248
rect 28264 29300 28316 29306
rect 28264 29242 28316 29248
rect 28724 29300 28776 29306
rect 28724 29242 28776 29248
rect 27988 29164 28040 29170
rect 27988 29106 28040 29112
rect 28172 29164 28224 29170
rect 28172 29106 28224 29112
rect 27896 29028 27948 29034
rect 27896 28970 27948 28976
rect 27908 28626 27936 28970
rect 27896 28620 27948 28626
rect 27896 28562 27948 28568
rect 27160 28552 27212 28558
rect 27160 28494 27212 28500
rect 27068 28484 27120 28490
rect 27068 28426 27120 28432
rect 26884 28416 26936 28422
rect 26884 28358 26936 28364
rect 27080 28218 27108 28426
rect 27068 28212 27120 28218
rect 27068 28154 27120 28160
rect 26792 27940 26844 27946
rect 26792 27882 26844 27888
rect 27172 27674 27200 28494
rect 27908 28218 27936 28562
rect 28000 28558 28028 29106
rect 28184 28762 28212 29106
rect 28172 28756 28224 28762
rect 28172 28698 28224 28704
rect 28276 28626 28304 29242
rect 28264 28620 28316 28626
rect 28264 28562 28316 28568
rect 27988 28552 28040 28558
rect 27988 28494 28040 28500
rect 27896 28212 27948 28218
rect 27896 28154 27948 28160
rect 27712 28008 27764 28014
rect 27712 27950 27764 27956
rect 27160 27668 27212 27674
rect 27160 27610 27212 27616
rect 27172 27470 27200 27610
rect 27160 27464 27212 27470
rect 27160 27406 27212 27412
rect 27160 27328 27212 27334
rect 27160 27270 27212 27276
rect 27344 27328 27396 27334
rect 27344 27270 27396 27276
rect 27436 27328 27488 27334
rect 27436 27270 27488 27276
rect 27172 26994 27200 27270
rect 27160 26988 27212 26994
rect 27160 26930 27212 26936
rect 27356 26926 27384 27270
rect 27448 26994 27476 27270
rect 27436 26988 27488 26994
rect 27436 26930 27488 26936
rect 27344 26920 27396 26926
rect 27344 26862 27396 26868
rect 27356 25498 27384 26862
rect 27448 26314 27476 26930
rect 27436 26308 27488 26314
rect 27436 26250 27488 26256
rect 27344 25492 27396 25498
rect 27344 25434 27396 25440
rect 26700 25288 26752 25294
rect 26700 25230 26752 25236
rect 26712 24818 26740 25230
rect 26700 24812 26752 24818
rect 26700 24754 26752 24760
rect 27160 24812 27212 24818
rect 27160 24754 27212 24760
rect 26608 24404 26660 24410
rect 26608 24346 26660 24352
rect 27172 24070 27200 24754
rect 27160 24064 27212 24070
rect 27160 24006 27212 24012
rect 26240 2644 26292 2650
rect 26240 2586 26292 2592
rect 25504 2576 25556 2582
rect 25504 2518 25556 2524
rect 23756 2372 23808 2378
rect 23756 2314 23808 2320
rect 24492 2372 24544 2378
rect 24492 2314 24544 2320
rect 24504 800 24532 2314
rect 24952 2304 25004 2310
rect 24952 2246 25004 2252
rect 26424 2304 26476 2310
rect 26424 2246 26476 2252
rect 24964 1970 24992 2246
rect 24952 1964 25004 1970
rect 24952 1906 25004 1912
rect 26436 800 26464 2246
rect 27172 2038 27200 24006
rect 27448 11626 27476 26250
rect 27724 25838 27752 27950
rect 28000 27674 28028 28494
rect 28816 28416 28868 28422
rect 28816 28358 28868 28364
rect 28828 28082 28856 28358
rect 28816 28076 28868 28082
rect 28816 28018 28868 28024
rect 28828 27878 28856 28018
rect 28816 27872 28868 27878
rect 28816 27814 28868 27820
rect 27988 27668 28040 27674
rect 27988 27610 28040 27616
rect 28448 26988 28500 26994
rect 28448 26930 28500 26936
rect 28460 26314 28488 26930
rect 28448 26308 28500 26314
rect 28448 26250 28500 26256
rect 28172 25900 28224 25906
rect 28172 25842 28224 25848
rect 27712 25832 27764 25838
rect 27712 25774 27764 25780
rect 28184 25498 28212 25842
rect 28172 25492 28224 25498
rect 28172 25434 28224 25440
rect 28264 25492 28316 25498
rect 28264 25434 28316 25440
rect 28276 25378 28304 25434
rect 28000 25350 28304 25378
rect 28000 25226 28028 25350
rect 28080 25288 28132 25294
rect 28080 25230 28132 25236
rect 28264 25288 28316 25294
rect 28264 25230 28316 25236
rect 27988 25220 28040 25226
rect 27988 25162 28040 25168
rect 28000 24818 28028 25162
rect 28092 24954 28120 25230
rect 28080 24948 28132 24954
rect 28080 24890 28132 24896
rect 27988 24812 28040 24818
rect 27988 24754 28040 24760
rect 28000 24410 28028 24754
rect 28276 24750 28304 25230
rect 28264 24744 28316 24750
rect 28264 24686 28316 24692
rect 27988 24404 28040 24410
rect 27988 24346 28040 24352
rect 27436 11620 27488 11626
rect 27436 11562 27488 11568
rect 28356 2848 28408 2854
rect 28356 2790 28408 2796
rect 28368 2378 28396 2790
rect 28460 2514 28488 26250
rect 28828 2990 28856 27814
rect 29012 27470 29040 30534
rect 29104 30394 29132 31350
rect 29196 30598 29224 33458
rect 29644 33108 29696 33114
rect 29644 33050 29696 33056
rect 29552 32904 29604 32910
rect 29552 32846 29604 32852
rect 29564 32570 29592 32846
rect 29656 32774 29684 33050
rect 29644 32768 29696 32774
rect 29644 32710 29696 32716
rect 29552 32564 29604 32570
rect 29552 32506 29604 32512
rect 29736 32428 29788 32434
rect 29736 32370 29788 32376
rect 29368 32360 29420 32366
rect 29368 32302 29420 32308
rect 29644 32360 29696 32366
rect 29644 32302 29696 32308
rect 29380 31822 29408 32302
rect 29656 31890 29684 32302
rect 29748 32230 29776 32370
rect 29736 32224 29788 32230
rect 29736 32166 29788 32172
rect 29644 31884 29696 31890
rect 29644 31826 29696 31832
rect 29368 31816 29420 31822
rect 29420 31776 29500 31804
rect 29368 31758 29420 31764
rect 29472 31482 29500 31776
rect 29460 31476 29512 31482
rect 29460 31418 29512 31424
rect 29460 31340 29512 31346
rect 29460 31282 29512 31288
rect 29472 30734 29500 31282
rect 29656 31142 29684 31826
rect 29840 31754 29868 35566
rect 30024 35193 30052 35770
rect 30116 35698 30144 36479
rect 30104 35692 30156 35698
rect 30104 35634 30156 35640
rect 30010 35184 30066 35193
rect 30010 35119 30066 35128
rect 29920 35080 29972 35086
rect 29920 35022 29972 35028
rect 29932 34785 29960 35022
rect 29918 34776 29974 34785
rect 29918 34711 29974 34720
rect 29932 34610 29960 34711
rect 29920 34604 29972 34610
rect 29920 34546 29972 34552
rect 29932 33658 29960 34546
rect 30104 34468 30156 34474
rect 30104 34410 30156 34416
rect 29920 33652 29972 33658
rect 29920 33594 29972 33600
rect 29932 33318 29960 33594
rect 29920 33312 29972 33318
rect 29920 33254 29972 33260
rect 29920 32428 29972 32434
rect 29920 32370 29972 32376
rect 29932 32026 29960 32370
rect 30012 32224 30064 32230
rect 30012 32166 30064 32172
rect 29920 32020 29972 32026
rect 29920 31962 29972 31968
rect 30024 31890 30052 32166
rect 30012 31884 30064 31890
rect 30012 31826 30064 31832
rect 29748 31726 29868 31754
rect 29644 31136 29696 31142
rect 29644 31078 29696 31084
rect 29460 30728 29512 30734
rect 29460 30670 29512 30676
rect 29276 30660 29328 30666
rect 29276 30602 29328 30608
rect 29184 30592 29236 30598
rect 29184 30534 29236 30540
rect 29092 30388 29144 30394
rect 29092 30330 29144 30336
rect 29104 30258 29132 30330
rect 29092 30252 29144 30258
rect 29092 30194 29144 30200
rect 29000 27464 29052 27470
rect 29000 27406 29052 27412
rect 29288 25498 29316 30602
rect 29368 29640 29420 29646
rect 29368 29582 29420 29588
rect 29380 29170 29408 29582
rect 29368 29164 29420 29170
rect 29368 29106 29420 29112
rect 29380 28626 29408 29106
rect 29368 28620 29420 28626
rect 29368 28562 29420 28568
rect 29472 28422 29500 30670
rect 29552 30592 29604 30598
rect 29552 30534 29604 30540
rect 29564 30190 29592 30534
rect 29644 30252 29696 30258
rect 29644 30194 29696 30200
rect 29552 30184 29604 30190
rect 29552 30126 29604 30132
rect 29552 30048 29604 30054
rect 29552 29990 29604 29996
rect 29564 29646 29592 29990
rect 29552 29640 29604 29646
rect 29552 29582 29604 29588
rect 29656 29510 29684 30194
rect 29748 29850 29776 31726
rect 30024 31346 30052 31826
rect 30012 31340 30064 31346
rect 30012 31282 30064 31288
rect 30024 30938 30052 31282
rect 30012 30932 30064 30938
rect 30012 30874 30064 30880
rect 30116 30598 30144 34410
rect 30208 31754 30236 37334
rect 30300 37244 30328 37703
rect 30380 37256 30432 37262
rect 30300 37216 30380 37244
rect 30380 37198 30432 37204
rect 30378 36816 30434 36825
rect 30378 36751 30380 36760
rect 30432 36751 30434 36760
rect 30380 36722 30432 36728
rect 30300 36378 30420 36394
rect 30300 36372 30432 36378
rect 30300 36366 30380 36372
rect 30300 35766 30328 36366
rect 30380 36314 30432 36320
rect 30484 36224 30512 39238
rect 30576 39098 30604 39374
rect 30564 39092 30616 39098
rect 30564 39034 30616 39040
rect 30564 38956 30616 38962
rect 30564 38898 30616 38904
rect 30576 38758 30604 38898
rect 30564 38752 30616 38758
rect 30564 38694 30616 38700
rect 30576 37874 30604 38694
rect 30564 37868 30616 37874
rect 30564 37810 30616 37816
rect 30562 37088 30618 37097
rect 30562 37023 30618 37032
rect 30576 36786 30604 37023
rect 30564 36780 30616 36786
rect 30564 36722 30616 36728
rect 30564 36576 30616 36582
rect 30564 36518 30616 36524
rect 30392 36196 30512 36224
rect 30288 35760 30340 35766
rect 30288 35702 30340 35708
rect 30288 35624 30340 35630
rect 30288 35566 30340 35572
rect 30300 35290 30328 35566
rect 30288 35284 30340 35290
rect 30288 35226 30340 35232
rect 30288 33924 30340 33930
rect 30288 33866 30340 33872
rect 30300 32910 30328 33866
rect 30392 33522 30420 36196
rect 30576 36174 30604 36518
rect 30564 36168 30616 36174
rect 30484 36128 30564 36156
rect 30484 35018 30512 36128
rect 30564 36110 30616 36116
rect 30668 35834 30696 42162
rect 30748 42152 30800 42158
rect 30748 42094 30800 42100
rect 30760 38962 30788 42094
rect 30852 41290 30880 43046
rect 30944 42158 30972 45018
rect 31024 42560 31076 42566
rect 31024 42502 31076 42508
rect 30932 42152 30984 42158
rect 30932 42094 30984 42100
rect 30852 41262 30972 41290
rect 30840 41200 30892 41206
rect 30840 41142 30892 41148
rect 30748 38956 30800 38962
rect 30748 38898 30800 38904
rect 30748 37868 30800 37874
rect 30748 37810 30800 37816
rect 30760 37262 30788 37810
rect 30748 37256 30800 37262
rect 30748 37198 30800 37204
rect 30760 36417 30788 37198
rect 30746 36408 30802 36417
rect 30852 36378 30880 41142
rect 30944 37874 30972 41262
rect 30932 37868 30984 37874
rect 30932 37810 30984 37816
rect 30944 37777 30972 37810
rect 30930 37768 30986 37777
rect 30930 37703 30986 37712
rect 31036 37448 31064 42502
rect 31206 41712 31262 41721
rect 31206 41647 31208 41656
rect 31260 41647 31262 41656
rect 31208 41618 31260 41624
rect 31312 40934 31340 46310
rect 31496 45626 31524 46514
rect 31576 46368 31628 46374
rect 31576 46310 31628 46316
rect 31484 45620 31536 45626
rect 31484 45562 31536 45568
rect 31484 44328 31536 44334
rect 31484 44270 31536 44276
rect 31496 42906 31524 44270
rect 31484 42900 31536 42906
rect 31484 42842 31536 42848
rect 31392 42628 31444 42634
rect 31392 42570 31444 42576
rect 31300 40928 31352 40934
rect 31300 40870 31352 40876
rect 31116 39840 31168 39846
rect 31116 39782 31168 39788
rect 30944 37420 31064 37448
rect 30746 36343 30802 36352
rect 30840 36372 30892 36378
rect 30840 36314 30892 36320
rect 30656 35828 30708 35834
rect 30656 35770 30708 35776
rect 30840 35692 30892 35698
rect 30840 35634 30892 35640
rect 30748 35624 30800 35630
rect 30576 35584 30748 35612
rect 30576 35086 30604 35584
rect 30748 35566 30800 35572
rect 30852 35442 30880 35634
rect 30668 35414 30880 35442
rect 30564 35080 30616 35086
rect 30564 35022 30616 35028
rect 30472 35012 30524 35018
rect 30472 34954 30524 34960
rect 30380 33516 30432 33522
rect 30380 33458 30432 33464
rect 30288 32904 30340 32910
rect 30288 32846 30340 32852
rect 30196 31748 30248 31754
rect 30196 31690 30248 31696
rect 30104 30592 30156 30598
rect 30104 30534 30156 30540
rect 29920 30252 29972 30258
rect 29920 30194 29972 30200
rect 29828 30048 29880 30054
rect 29828 29990 29880 29996
rect 29736 29844 29788 29850
rect 29736 29786 29788 29792
rect 29840 29646 29868 29990
rect 29828 29640 29880 29646
rect 29828 29582 29880 29588
rect 29644 29504 29696 29510
rect 29644 29446 29696 29452
rect 29656 28762 29684 29446
rect 29736 29232 29788 29238
rect 29736 29174 29788 29180
rect 29644 28756 29696 28762
rect 29644 28698 29696 28704
rect 29748 28558 29776 29174
rect 29932 29170 29960 30194
rect 30196 30184 30248 30190
rect 30196 30126 30248 30132
rect 30208 29170 30236 30126
rect 29920 29164 29972 29170
rect 29920 29106 29972 29112
rect 30104 29164 30156 29170
rect 30104 29106 30156 29112
rect 30196 29164 30248 29170
rect 30196 29106 30248 29112
rect 29736 28552 29788 28558
rect 29736 28494 29788 28500
rect 29460 28416 29512 28422
rect 29460 28358 29512 28364
rect 29748 28218 29776 28494
rect 29932 28218 29960 29106
rect 29736 28212 29788 28218
rect 29736 28154 29788 28160
rect 29920 28212 29972 28218
rect 29920 28154 29972 28160
rect 29828 26988 29880 26994
rect 29828 26930 29880 26936
rect 29840 26586 29868 26930
rect 30116 26858 30144 29106
rect 30208 28762 30236 29106
rect 30392 28778 30420 33458
rect 30576 33454 30604 35022
rect 30472 33448 30524 33454
rect 30472 33390 30524 33396
rect 30564 33448 30616 33454
rect 30564 33390 30616 33396
rect 30484 33114 30512 33390
rect 30472 33108 30524 33114
rect 30472 33050 30524 33056
rect 30564 32904 30616 32910
rect 30484 32864 30564 32892
rect 30484 31822 30512 32864
rect 30564 32846 30616 32852
rect 30668 32552 30696 35414
rect 30840 35284 30892 35290
rect 30840 35226 30892 35232
rect 30852 35154 30880 35226
rect 30840 35148 30892 35154
rect 30840 35090 30892 35096
rect 30748 35012 30800 35018
rect 30748 34954 30800 34960
rect 30760 34746 30788 34954
rect 30944 34921 30972 37420
rect 31128 37369 31156 39782
rect 31312 39386 31340 40870
rect 31404 39574 31432 42570
rect 31392 39568 31444 39574
rect 31392 39510 31444 39516
rect 31208 39364 31260 39370
rect 31312 39358 31432 39386
rect 31208 39306 31260 39312
rect 31114 37360 31170 37369
rect 31024 37324 31076 37330
rect 31114 37295 31170 37304
rect 31024 37266 31076 37272
rect 30930 34912 30986 34921
rect 30930 34847 30986 34856
rect 30748 34740 30800 34746
rect 30748 34682 30800 34688
rect 30746 34640 30802 34649
rect 30746 34575 30748 34584
rect 30800 34575 30802 34584
rect 30748 34546 30800 34552
rect 30840 34536 30892 34542
rect 30840 34478 30892 34484
rect 30852 34134 30880 34478
rect 30840 34128 30892 34134
rect 30840 34070 30892 34076
rect 30852 33658 30880 34070
rect 30932 33992 30984 33998
rect 30932 33934 30984 33940
rect 30840 33652 30892 33658
rect 30840 33594 30892 33600
rect 30840 32768 30892 32774
rect 30840 32710 30892 32716
rect 30576 32524 30696 32552
rect 30472 31816 30524 31822
rect 30472 31758 30524 31764
rect 30484 31482 30512 31758
rect 30472 31476 30524 31482
rect 30472 31418 30524 31424
rect 30576 29850 30604 32524
rect 30852 32502 30880 32710
rect 30748 32496 30800 32502
rect 30748 32438 30800 32444
rect 30840 32496 30892 32502
rect 30840 32438 30892 32444
rect 30656 32428 30708 32434
rect 30656 32370 30708 32376
rect 30668 32026 30696 32370
rect 30656 32020 30708 32026
rect 30656 31962 30708 31968
rect 30760 31958 30788 32438
rect 30944 32298 30972 33934
rect 31036 32892 31064 37266
rect 31114 36952 31170 36961
rect 31114 36887 31170 36896
rect 31128 36854 31156 36887
rect 31116 36848 31168 36854
rect 31116 36790 31168 36796
rect 31116 36712 31168 36718
rect 31116 36654 31168 36660
rect 31128 33046 31156 36654
rect 31220 34649 31248 39306
rect 31404 38894 31432 39358
rect 31496 39284 31524 42842
rect 31588 39438 31616 46310
rect 31668 46164 31720 46170
rect 31668 46106 31720 46112
rect 31680 45626 31708 46106
rect 31760 45892 31812 45898
rect 31760 45834 31812 45840
rect 31668 45620 31720 45626
rect 31668 45562 31720 45568
rect 31772 42650 31800 45834
rect 31680 42622 31800 42650
rect 31680 42242 31708 42622
rect 31760 42560 31812 42566
rect 31760 42502 31812 42508
rect 31772 42362 31800 42502
rect 31760 42356 31812 42362
rect 31760 42298 31812 42304
rect 31852 42288 31904 42294
rect 31680 42214 31800 42242
rect 31852 42230 31904 42236
rect 31772 41041 31800 42214
rect 31864 42158 31892 42230
rect 31852 42152 31904 42158
rect 31852 42094 31904 42100
rect 31758 41032 31814 41041
rect 31758 40967 31814 40976
rect 31760 40520 31812 40526
rect 31760 40462 31812 40468
rect 31772 39574 31800 40462
rect 31760 39568 31812 39574
rect 31760 39510 31812 39516
rect 31956 39506 31984 46922
rect 32140 46578 32168 46990
rect 32508 46986 32536 47602
rect 32496 46980 32548 46986
rect 32496 46922 32548 46928
rect 32128 46572 32180 46578
rect 32128 46514 32180 46520
rect 32128 45960 32180 45966
rect 32128 45902 32180 45908
rect 32140 45490 32168 45902
rect 32128 45484 32180 45490
rect 32128 45426 32180 45432
rect 32034 45384 32090 45393
rect 32034 45319 32036 45328
rect 32088 45319 32090 45328
rect 32036 45290 32088 45296
rect 32140 45234 32168 45426
rect 32048 45206 32168 45234
rect 32048 44946 32076 45206
rect 32036 44940 32088 44946
rect 32036 44882 32088 44888
rect 32048 44470 32076 44882
rect 32312 44736 32364 44742
rect 32312 44678 32364 44684
rect 32036 44464 32088 44470
rect 32036 44406 32088 44412
rect 32048 43654 32076 44406
rect 32036 43648 32088 43654
rect 32036 43590 32088 43596
rect 32048 43382 32076 43590
rect 32036 43376 32088 43382
rect 32036 43318 32088 43324
rect 32048 42770 32076 43318
rect 32220 43104 32272 43110
rect 32220 43046 32272 43052
rect 32036 42764 32088 42770
rect 32036 42706 32088 42712
rect 32128 42152 32180 42158
rect 32128 42094 32180 42100
rect 32036 42084 32088 42090
rect 32036 42026 32088 42032
rect 32048 39982 32076 42026
rect 32140 41138 32168 42094
rect 32128 41132 32180 41138
rect 32128 41074 32180 41080
rect 32232 40633 32260 43046
rect 32324 40662 32352 44678
rect 32404 41608 32456 41614
rect 32404 41550 32456 41556
rect 32312 40656 32364 40662
rect 32218 40624 32274 40633
rect 32312 40598 32364 40604
rect 32218 40559 32274 40568
rect 32324 40390 32352 40598
rect 32416 40458 32444 41550
rect 32508 41478 32536 46922
rect 32876 46714 32904 49200
rect 34336 47252 34388 47258
rect 34336 47194 34388 47200
rect 33876 47184 33928 47190
rect 33876 47126 33928 47132
rect 32864 46708 32916 46714
rect 32864 46650 32916 46656
rect 33888 45558 33916 47126
rect 33968 46572 34020 46578
rect 33968 46514 34020 46520
rect 34060 46572 34112 46578
rect 34060 46514 34112 46520
rect 33876 45552 33928 45558
rect 33876 45494 33928 45500
rect 33232 45484 33284 45490
rect 33232 45426 33284 45432
rect 33244 43761 33272 45426
rect 33888 45286 33916 45494
rect 33876 45280 33928 45286
rect 33876 45222 33928 45228
rect 33784 44872 33836 44878
rect 33784 44814 33836 44820
rect 33324 44396 33376 44402
rect 33324 44338 33376 44344
rect 33230 43752 33286 43761
rect 33230 43687 33286 43696
rect 33140 43648 33192 43654
rect 33140 43590 33192 43596
rect 33152 42022 33180 43590
rect 33336 43450 33364 44338
rect 33600 44192 33652 44198
rect 33600 44134 33652 44140
rect 33324 43444 33376 43450
rect 33324 43386 33376 43392
rect 33324 43308 33376 43314
rect 33324 43250 33376 43256
rect 33336 43217 33364 43250
rect 33322 43208 33378 43217
rect 33322 43143 33378 43152
rect 33612 42158 33640 44134
rect 33692 43376 33744 43382
rect 33692 43318 33744 43324
rect 33600 42152 33652 42158
rect 33600 42094 33652 42100
rect 33140 42016 33192 42022
rect 33140 41958 33192 41964
rect 32496 41472 32548 41478
rect 32494 41440 32496 41449
rect 32548 41440 32550 41449
rect 32494 41375 32550 41384
rect 32680 41132 32732 41138
rect 32680 41074 32732 41080
rect 32692 40730 32720 41074
rect 32496 40724 32548 40730
rect 32496 40666 32548 40672
rect 32680 40724 32732 40730
rect 32680 40666 32732 40672
rect 32404 40452 32456 40458
rect 32404 40394 32456 40400
rect 32312 40384 32364 40390
rect 32508 40361 32536 40666
rect 32494 40352 32550 40361
rect 32312 40326 32364 40332
rect 32416 40310 32494 40338
rect 32128 40112 32180 40118
rect 32128 40054 32180 40060
rect 32036 39976 32088 39982
rect 32036 39918 32088 39924
rect 31944 39500 31996 39506
rect 31944 39442 31996 39448
rect 31576 39432 31628 39438
rect 31576 39374 31628 39380
rect 31496 39256 31708 39284
rect 31392 38888 31444 38894
rect 31392 38830 31444 38836
rect 31576 38888 31628 38894
rect 31576 38830 31628 38836
rect 31300 38752 31352 38758
rect 31300 38694 31352 38700
rect 31312 37874 31340 38694
rect 31390 38448 31446 38457
rect 31390 38383 31392 38392
rect 31444 38383 31446 38392
rect 31392 38354 31444 38360
rect 31482 38040 31538 38049
rect 31482 37975 31538 37984
rect 31300 37868 31352 37874
rect 31300 37810 31352 37816
rect 31392 37256 31444 37262
rect 31392 37198 31444 37204
rect 31404 37097 31432 37198
rect 31390 37088 31446 37097
rect 31390 37023 31446 37032
rect 31496 36938 31524 37975
rect 31404 36910 31524 36938
rect 31298 36816 31354 36825
rect 31298 36751 31300 36760
rect 31352 36751 31354 36760
rect 31300 36722 31352 36728
rect 31300 36576 31352 36582
rect 31300 36518 31352 36524
rect 31312 36310 31340 36518
rect 31404 36378 31432 36910
rect 31484 36712 31536 36718
rect 31484 36654 31536 36660
rect 31392 36372 31444 36378
rect 31392 36314 31444 36320
rect 31300 36304 31352 36310
rect 31300 36246 31352 36252
rect 31496 36174 31524 36654
rect 31484 36168 31536 36174
rect 31484 36110 31536 36116
rect 31300 36100 31352 36106
rect 31352 36060 31432 36088
rect 31300 36042 31352 36048
rect 31300 35828 31352 35834
rect 31300 35770 31352 35776
rect 31312 35290 31340 35770
rect 31300 35284 31352 35290
rect 31300 35226 31352 35232
rect 31300 34672 31352 34678
rect 31206 34640 31262 34649
rect 31300 34614 31352 34620
rect 31404 34626 31432 36060
rect 31496 35698 31524 36110
rect 31484 35692 31536 35698
rect 31484 35634 31536 35640
rect 31496 34746 31524 35634
rect 31588 35222 31616 38830
rect 31576 35216 31628 35222
rect 31576 35158 31628 35164
rect 31588 34746 31616 35158
rect 31484 34740 31536 34746
rect 31484 34682 31536 34688
rect 31576 34740 31628 34746
rect 31576 34682 31628 34688
rect 31206 34575 31262 34584
rect 31312 33998 31340 34614
rect 31404 34598 31616 34626
rect 31392 34196 31444 34202
rect 31392 34138 31444 34144
rect 31300 33992 31352 33998
rect 31300 33934 31352 33940
rect 31312 33522 31340 33934
rect 31404 33930 31432 34138
rect 31392 33924 31444 33930
rect 31392 33866 31444 33872
rect 31404 33522 31432 33866
rect 31588 33862 31616 34598
rect 31576 33856 31628 33862
rect 31576 33798 31628 33804
rect 31484 33652 31536 33658
rect 31484 33594 31536 33600
rect 31300 33516 31352 33522
rect 31300 33458 31352 33464
rect 31392 33516 31444 33522
rect 31392 33458 31444 33464
rect 31116 33040 31168 33046
rect 31116 32982 31168 32988
rect 31036 32864 31248 32892
rect 30932 32292 30984 32298
rect 30932 32234 30984 32240
rect 30840 32224 30892 32230
rect 30840 32166 30892 32172
rect 30852 32026 30880 32166
rect 30840 32020 30892 32026
rect 30840 31962 30892 31968
rect 30748 31952 30800 31958
rect 30748 31894 30800 31900
rect 30748 31816 30800 31822
rect 30748 31758 30800 31764
rect 30656 31680 30708 31686
rect 30656 31622 30708 31628
rect 30668 31346 30696 31622
rect 30656 31340 30708 31346
rect 30656 31282 30708 31288
rect 30668 30734 30696 31282
rect 30760 30938 30788 31758
rect 31024 31340 31076 31346
rect 31024 31282 31076 31288
rect 30748 30932 30800 30938
rect 30748 30874 30800 30880
rect 30656 30728 30708 30734
rect 30656 30670 30708 30676
rect 31036 30666 31064 31282
rect 31024 30660 31076 30666
rect 31024 30602 31076 30608
rect 30472 29844 30524 29850
rect 30472 29786 30524 29792
rect 30564 29844 30616 29850
rect 30564 29786 30616 29792
rect 30484 29306 30512 29786
rect 30932 29504 30984 29510
rect 30932 29446 30984 29452
rect 30944 29306 30972 29446
rect 30472 29300 30524 29306
rect 30472 29242 30524 29248
rect 30932 29300 30984 29306
rect 30932 29242 30984 29248
rect 30196 28756 30248 28762
rect 30392 28750 30512 28778
rect 30196 28698 30248 28704
rect 30380 28620 30432 28626
rect 30380 28562 30432 28568
rect 30196 28552 30248 28558
rect 30196 28494 30248 28500
rect 30208 28082 30236 28494
rect 30392 28082 30420 28562
rect 30196 28076 30248 28082
rect 30196 28018 30248 28024
rect 30380 28076 30432 28082
rect 30380 28018 30432 28024
rect 30104 26852 30156 26858
rect 30104 26794 30156 26800
rect 29828 26580 29880 26586
rect 29828 26522 29880 26528
rect 29828 26376 29880 26382
rect 29828 26318 29880 26324
rect 29840 25838 29868 26318
rect 30208 26042 30236 28018
rect 30484 27130 30512 28750
rect 31024 28416 31076 28422
rect 31024 28358 31076 28364
rect 30838 28112 30894 28121
rect 31036 28082 31064 28358
rect 30838 28047 30840 28056
rect 30892 28047 30894 28056
rect 31024 28076 31076 28082
rect 30840 28018 30892 28024
rect 31024 28018 31076 28024
rect 30852 27674 30880 28018
rect 30840 27668 30892 27674
rect 30840 27610 30892 27616
rect 30852 27470 30880 27610
rect 30840 27464 30892 27470
rect 30840 27406 30892 27412
rect 31036 27402 31064 28018
rect 31116 27464 31168 27470
rect 31116 27406 31168 27412
rect 30656 27396 30708 27402
rect 30656 27338 30708 27344
rect 31024 27396 31076 27402
rect 31024 27338 31076 27344
rect 30472 27124 30524 27130
rect 30472 27066 30524 27072
rect 30668 26994 30696 27338
rect 31128 26994 31156 27406
rect 31220 27062 31248 32864
rect 31300 31680 31352 31686
rect 31298 31648 31300 31657
rect 31352 31648 31354 31657
rect 31298 31583 31354 31592
rect 31404 31346 31432 33458
rect 31496 33318 31524 33594
rect 31484 33312 31536 33318
rect 31484 33254 31536 33260
rect 31496 32570 31524 33254
rect 31484 32564 31536 32570
rect 31484 32506 31536 32512
rect 31496 31414 31524 32506
rect 31588 32502 31616 33798
rect 31576 32496 31628 32502
rect 31576 32438 31628 32444
rect 31484 31408 31536 31414
rect 31484 31350 31536 31356
rect 31392 31340 31444 31346
rect 31392 31282 31444 31288
rect 31404 30734 31432 31282
rect 31484 31272 31536 31278
rect 31484 31214 31536 31220
rect 31496 31142 31524 31214
rect 31484 31136 31536 31142
rect 31484 31078 31536 31084
rect 31392 30728 31444 30734
rect 31392 30670 31444 30676
rect 31392 30252 31444 30258
rect 31392 30194 31444 30200
rect 31404 29782 31432 30194
rect 31484 30184 31536 30190
rect 31484 30126 31536 30132
rect 31496 30054 31524 30126
rect 31484 30048 31536 30054
rect 31484 29990 31536 29996
rect 31392 29776 31444 29782
rect 31392 29718 31444 29724
rect 31496 29646 31524 29990
rect 31484 29640 31536 29646
rect 31484 29582 31536 29588
rect 31208 27056 31260 27062
rect 31208 26998 31260 27004
rect 30288 26988 30340 26994
rect 30288 26930 30340 26936
rect 30472 26988 30524 26994
rect 30472 26930 30524 26936
rect 30656 26988 30708 26994
rect 30656 26930 30708 26936
rect 31116 26988 31168 26994
rect 31116 26930 31168 26936
rect 30300 26450 30328 26930
rect 30380 26784 30432 26790
rect 30380 26726 30432 26732
rect 30288 26444 30340 26450
rect 30288 26386 30340 26392
rect 30196 26036 30248 26042
rect 30196 25978 30248 25984
rect 30392 25906 30420 26726
rect 30484 26246 30512 26930
rect 30668 26586 30696 26930
rect 30656 26580 30708 26586
rect 30656 26522 30708 26528
rect 30472 26240 30524 26246
rect 30472 26182 30524 26188
rect 30380 25900 30432 25906
rect 30380 25842 30432 25848
rect 29828 25832 29880 25838
rect 29828 25774 29880 25780
rect 29276 25492 29328 25498
rect 29276 25434 29328 25440
rect 29840 25430 29868 25774
rect 29828 25424 29880 25430
rect 29828 25366 29880 25372
rect 28816 2984 28868 2990
rect 28816 2926 28868 2932
rect 30668 2514 30696 26522
rect 31128 26466 31156 26930
rect 31128 26438 31248 26466
rect 31116 26308 31168 26314
rect 31116 26250 31168 26256
rect 31024 26240 31076 26246
rect 31024 26182 31076 26188
rect 31036 26042 31064 26182
rect 31024 26036 31076 26042
rect 31024 25978 31076 25984
rect 31128 25906 31156 26250
rect 31116 25900 31168 25906
rect 31116 25842 31168 25848
rect 31128 25498 31156 25842
rect 31116 25492 31168 25498
rect 31116 25434 31168 25440
rect 31220 22094 31248 26438
rect 31576 26444 31628 26450
rect 31576 26386 31628 26392
rect 31588 25906 31616 26386
rect 31576 25900 31628 25906
rect 31576 25842 31628 25848
rect 31588 25498 31616 25842
rect 31576 25492 31628 25498
rect 31576 25434 31628 25440
rect 31128 22066 31248 22094
rect 31128 9926 31156 22066
rect 31680 10062 31708 39256
rect 31944 39092 31996 39098
rect 31944 39034 31996 39040
rect 31760 38956 31812 38962
rect 31760 38898 31812 38904
rect 31772 37913 31800 38898
rect 31758 37904 31814 37913
rect 31758 37839 31814 37848
rect 31760 37324 31812 37330
rect 31760 37266 31812 37272
rect 31772 36038 31800 37266
rect 31956 36582 31984 39034
rect 32036 37868 32088 37874
rect 32036 37810 32088 37816
rect 32048 37262 32076 37810
rect 32036 37256 32088 37262
rect 32036 37198 32088 37204
rect 31944 36576 31996 36582
rect 31944 36518 31996 36524
rect 32048 36258 32076 37198
rect 31864 36242 32076 36258
rect 31852 36236 32076 36242
rect 31904 36230 32076 36236
rect 31852 36178 31904 36184
rect 31944 36168 31996 36174
rect 31944 36110 31996 36116
rect 31760 36032 31812 36038
rect 31760 35974 31812 35980
rect 31956 35154 31984 36110
rect 32048 35290 32076 36230
rect 32036 35284 32088 35290
rect 32036 35226 32088 35232
rect 31944 35148 31996 35154
rect 31944 35090 31996 35096
rect 32048 35086 32076 35226
rect 32036 35080 32088 35086
rect 32036 35022 32088 35028
rect 32140 35018 32168 40054
rect 32312 40044 32364 40050
rect 32312 39986 32364 39992
rect 32324 38758 32352 39986
rect 32416 39098 32444 40310
rect 32494 40287 32550 40296
rect 32508 40227 32536 40287
rect 32692 39506 32720 40666
rect 32770 39944 32826 39953
rect 32770 39879 32826 39888
rect 32680 39500 32732 39506
rect 32680 39442 32732 39448
rect 32784 39137 32812 39879
rect 32864 39840 32916 39846
rect 32864 39782 32916 39788
rect 32770 39128 32826 39137
rect 32404 39092 32456 39098
rect 32770 39063 32826 39072
rect 32404 39034 32456 39040
rect 32784 39030 32812 39063
rect 32772 39024 32824 39030
rect 32772 38966 32824 38972
rect 32496 38956 32548 38962
rect 32496 38898 32548 38904
rect 32404 38820 32456 38826
rect 32404 38762 32456 38768
rect 32312 38752 32364 38758
rect 32312 38694 32364 38700
rect 32324 36718 32352 38694
rect 32312 36712 32364 36718
rect 32312 36654 32364 36660
rect 32220 36032 32272 36038
rect 32220 35974 32272 35980
rect 32232 35698 32260 35974
rect 32220 35692 32272 35698
rect 32220 35634 32272 35640
rect 31944 35012 31996 35018
rect 31944 34954 31996 34960
rect 32128 35012 32180 35018
rect 32128 34954 32180 34960
rect 31760 34944 31812 34950
rect 31760 34886 31812 34892
rect 31772 34610 31800 34886
rect 31760 34604 31812 34610
rect 31760 34546 31812 34552
rect 31956 33590 31984 34954
rect 32218 34912 32274 34921
rect 32218 34847 32274 34856
rect 32232 34746 32260 34847
rect 32220 34740 32272 34746
rect 32220 34682 32272 34688
rect 32324 34066 32352 36654
rect 32416 36650 32444 38762
rect 32508 37194 32536 38898
rect 32876 38826 32904 39782
rect 33048 39500 33100 39506
rect 33048 39442 33100 39448
rect 32864 38820 32916 38826
rect 32864 38762 32916 38768
rect 32876 38554 32904 38762
rect 32864 38548 32916 38554
rect 32864 38490 32916 38496
rect 33060 38434 33088 39442
rect 33152 39370 33180 41958
rect 33612 41614 33640 42094
rect 33704 41682 33732 43318
rect 33796 42702 33824 44814
rect 33876 44736 33928 44742
rect 33876 44678 33928 44684
rect 33888 42702 33916 44678
rect 33980 44538 34008 46514
rect 34072 46170 34100 46514
rect 34060 46164 34112 46170
rect 34060 46106 34112 46112
rect 34060 45280 34112 45286
rect 34060 45222 34112 45228
rect 34072 44878 34100 45222
rect 34060 44872 34112 44878
rect 34060 44814 34112 44820
rect 33968 44532 34020 44538
rect 33968 44474 34020 44480
rect 34072 43858 34100 44814
rect 34060 43852 34112 43858
rect 34060 43794 34112 43800
rect 34060 43648 34112 43654
rect 34060 43590 34112 43596
rect 34072 42906 34100 43590
rect 34060 42900 34112 42906
rect 34060 42842 34112 42848
rect 33784 42696 33836 42702
rect 33784 42638 33836 42644
rect 33876 42696 33928 42702
rect 33876 42638 33928 42644
rect 33888 42090 33916 42638
rect 34244 42628 34296 42634
rect 34244 42570 34296 42576
rect 34152 42288 34204 42294
rect 34152 42230 34204 42236
rect 33876 42084 33928 42090
rect 33876 42026 33928 42032
rect 33692 41676 33744 41682
rect 33692 41618 33744 41624
rect 33888 41614 33916 42026
rect 33416 41608 33468 41614
rect 33416 41550 33468 41556
rect 33600 41608 33652 41614
rect 33600 41550 33652 41556
rect 33876 41608 33928 41614
rect 33876 41550 33928 41556
rect 33324 41472 33376 41478
rect 33324 41414 33376 41420
rect 33232 40928 33284 40934
rect 33232 40870 33284 40876
rect 33244 40526 33272 40870
rect 33336 40594 33364 41414
rect 33324 40588 33376 40594
rect 33324 40530 33376 40536
rect 33232 40520 33284 40526
rect 33232 40462 33284 40468
rect 33244 40050 33272 40462
rect 33232 40044 33284 40050
rect 33232 39986 33284 39992
rect 33428 39914 33456 41550
rect 33612 41414 33640 41550
rect 33784 41472 33836 41478
rect 33784 41414 33836 41420
rect 33888 41414 33916 41550
rect 33612 41386 33732 41414
rect 33508 40928 33560 40934
rect 33508 40870 33560 40876
rect 33520 40089 33548 40870
rect 33600 40588 33652 40594
rect 33600 40530 33652 40536
rect 33506 40080 33562 40089
rect 33612 40050 33640 40530
rect 33506 40015 33562 40024
rect 33600 40044 33652 40050
rect 33600 39986 33652 39992
rect 33704 39930 33732 41386
rect 33796 41274 33824 41414
rect 33888 41386 34100 41414
rect 33784 41268 33836 41274
rect 33784 41210 33836 41216
rect 33876 40656 33928 40662
rect 33876 40598 33928 40604
rect 33784 40044 33836 40050
rect 33784 39986 33836 39992
rect 33416 39908 33468 39914
rect 33416 39850 33468 39856
rect 33612 39902 33732 39930
rect 33612 39370 33640 39902
rect 33692 39432 33744 39438
rect 33692 39374 33744 39380
rect 33140 39364 33192 39370
rect 33140 39306 33192 39312
rect 33416 39364 33468 39370
rect 33416 39306 33468 39312
rect 33600 39364 33652 39370
rect 33600 39306 33652 39312
rect 33428 39098 33456 39306
rect 33508 39296 33560 39302
rect 33508 39238 33560 39244
rect 33416 39092 33468 39098
rect 33416 39034 33468 39040
rect 33520 39030 33548 39238
rect 33508 39024 33560 39030
rect 33508 38966 33560 38972
rect 33600 39024 33652 39030
rect 33600 38966 33652 38972
rect 32876 38406 33180 38434
rect 32772 38344 32824 38350
rect 32692 38292 32772 38298
rect 32692 38286 32824 38292
rect 32692 38270 32812 38286
rect 32588 37868 32640 37874
rect 32588 37810 32640 37816
rect 32600 37466 32628 37810
rect 32692 37738 32720 38270
rect 32770 37904 32826 37913
rect 32770 37839 32772 37848
rect 32824 37839 32826 37848
rect 32772 37810 32824 37816
rect 32680 37732 32732 37738
rect 32680 37674 32732 37680
rect 32588 37460 32640 37466
rect 32588 37402 32640 37408
rect 32586 37224 32642 37233
rect 32496 37188 32548 37194
rect 32876 37194 32904 38406
rect 33152 38350 33180 38406
rect 33232 38412 33284 38418
rect 33232 38354 33284 38360
rect 33048 38344 33100 38350
rect 33048 38286 33100 38292
rect 33140 38344 33192 38350
rect 33140 38286 33192 38292
rect 32956 38208 33008 38214
rect 32956 38150 33008 38156
rect 32586 37159 32642 37168
rect 32864 37188 32916 37194
rect 32496 37130 32548 37136
rect 32496 36780 32548 36786
rect 32600 36768 32628 37159
rect 32864 37130 32916 37136
rect 32772 36848 32824 36854
rect 32772 36790 32824 36796
rect 32548 36740 32628 36768
rect 32496 36722 32548 36728
rect 32404 36644 32456 36650
rect 32404 36586 32456 36592
rect 32496 36576 32548 36582
rect 32496 36518 32548 36524
rect 32404 35692 32456 35698
rect 32404 35634 32456 35640
rect 32416 35057 32444 35634
rect 32402 35048 32458 35057
rect 32402 34983 32404 34992
rect 32456 34983 32458 34992
rect 32404 34954 32456 34960
rect 32402 34232 32458 34241
rect 32402 34167 32404 34176
rect 32456 34167 32458 34176
rect 32404 34138 32456 34144
rect 32312 34060 32364 34066
rect 32312 34002 32364 34008
rect 32508 33810 32536 36518
rect 32784 36378 32812 36790
rect 32968 36786 32996 38150
rect 33060 38010 33088 38286
rect 33048 38004 33100 38010
rect 33048 37946 33100 37952
rect 33140 38004 33192 38010
rect 33140 37946 33192 37952
rect 33048 36916 33100 36922
rect 33048 36858 33100 36864
rect 32956 36780 33008 36786
rect 32956 36722 33008 36728
rect 32772 36372 32824 36378
rect 32772 36314 32824 36320
rect 33060 36174 33088 36858
rect 33048 36168 33100 36174
rect 33048 36110 33100 36116
rect 33152 35834 33180 37946
rect 33140 35828 33192 35834
rect 33140 35770 33192 35776
rect 33244 35290 33272 38354
rect 33416 38276 33468 38282
rect 33416 38218 33468 38224
rect 33428 37466 33456 38218
rect 33520 38010 33548 38966
rect 33612 38758 33640 38966
rect 33704 38962 33732 39374
rect 33692 38956 33744 38962
rect 33692 38898 33744 38904
rect 33704 38826 33732 38898
rect 33692 38820 33744 38826
rect 33692 38762 33744 38768
rect 33600 38752 33652 38758
rect 33600 38694 33652 38700
rect 33600 38480 33652 38486
rect 33600 38422 33652 38428
rect 33508 38004 33560 38010
rect 33508 37946 33560 37952
rect 33508 37868 33560 37874
rect 33508 37810 33560 37816
rect 33416 37460 33468 37466
rect 33416 37402 33468 37408
rect 33520 37126 33548 37810
rect 33612 37670 33640 38422
rect 33704 38350 33732 38762
rect 33692 38344 33744 38350
rect 33692 38286 33744 38292
rect 33796 38298 33824 39986
rect 33888 38400 33916 40598
rect 33968 40112 34020 40118
rect 33968 40054 34020 40060
rect 33980 39574 34008 40054
rect 33968 39568 34020 39574
rect 33968 39510 34020 39516
rect 33968 39432 34020 39438
rect 33968 39374 34020 39380
rect 33980 38554 34008 39374
rect 33968 38548 34020 38554
rect 33968 38490 34020 38496
rect 33888 38372 34008 38400
rect 33980 38321 34008 38372
rect 33966 38312 34022 38321
rect 33796 38270 33916 38298
rect 33600 37664 33652 37670
rect 33600 37606 33652 37612
rect 33692 37664 33744 37670
rect 33692 37606 33744 37612
rect 33704 37262 33732 37606
rect 33888 37346 33916 38270
rect 33966 38247 34022 38256
rect 33796 37318 33916 37346
rect 33692 37256 33744 37262
rect 33692 37198 33744 37204
rect 33508 37120 33560 37126
rect 33508 37062 33560 37068
rect 33520 36854 33548 37062
rect 33508 36848 33560 36854
rect 33508 36790 33560 36796
rect 33324 36576 33376 36582
rect 33324 36518 33376 36524
rect 33232 35284 33284 35290
rect 33232 35226 33284 35232
rect 33336 34610 33364 36518
rect 33416 35828 33468 35834
rect 33416 35770 33468 35776
rect 33428 35086 33456 35770
rect 33520 35698 33548 36790
rect 33600 36780 33652 36786
rect 33600 36722 33652 36728
rect 33508 35692 33560 35698
rect 33508 35634 33560 35640
rect 33520 35290 33548 35634
rect 33612 35630 33640 36722
rect 33692 36168 33744 36174
rect 33692 36110 33744 36116
rect 33704 35834 33732 36110
rect 33796 35986 33824 37318
rect 33876 37256 33928 37262
rect 33876 37198 33928 37204
rect 33888 37097 33916 37198
rect 33874 37088 33930 37097
rect 33874 37023 33930 37032
rect 33876 36576 33928 36582
rect 33876 36518 33928 36524
rect 33888 36417 33916 36518
rect 33874 36408 33930 36417
rect 33874 36343 33930 36352
rect 33888 36174 33916 36343
rect 33876 36168 33928 36174
rect 33876 36110 33928 36116
rect 33796 35958 33916 35986
rect 33692 35828 33744 35834
rect 33692 35770 33744 35776
rect 33600 35624 33652 35630
rect 33600 35566 33652 35572
rect 33508 35284 33560 35290
rect 33508 35226 33560 35232
rect 33612 35222 33640 35566
rect 33600 35216 33652 35222
rect 33600 35158 33652 35164
rect 33416 35080 33468 35086
rect 33416 35022 33468 35028
rect 33784 35080 33836 35086
rect 33784 35022 33836 35028
rect 33414 34776 33470 34785
rect 33414 34711 33416 34720
rect 33468 34711 33470 34720
rect 33416 34682 33468 34688
rect 33324 34604 33376 34610
rect 33324 34546 33376 34552
rect 33600 34604 33652 34610
rect 33600 34546 33652 34552
rect 33046 34232 33102 34241
rect 33046 34167 33102 34176
rect 33060 33930 33088 34167
rect 33140 34060 33192 34066
rect 33140 34002 33192 34008
rect 33048 33924 33100 33930
rect 33048 33866 33100 33872
rect 32324 33782 32536 33810
rect 31944 33584 31996 33590
rect 31944 33526 31996 33532
rect 32128 33448 32180 33454
rect 32128 33390 32180 33396
rect 32140 32978 32168 33390
rect 32220 33312 32272 33318
rect 32220 33254 32272 33260
rect 32128 32972 32180 32978
rect 32128 32914 32180 32920
rect 32128 32496 32180 32502
rect 32128 32438 32180 32444
rect 32140 31822 32168 32438
rect 32232 31890 32260 33254
rect 32220 31884 32272 31890
rect 32220 31826 32272 31832
rect 32128 31816 32180 31822
rect 32128 31758 32180 31764
rect 32140 31346 32168 31758
rect 32220 31748 32272 31754
rect 32220 31690 32272 31696
rect 32128 31340 32180 31346
rect 32128 31282 32180 31288
rect 32232 30734 32260 31690
rect 32220 30728 32272 30734
rect 32220 30670 32272 30676
rect 32036 30660 32088 30666
rect 32036 30602 32088 30608
rect 32048 29510 32076 30602
rect 32232 30258 32260 30670
rect 32220 30252 32272 30258
rect 32220 30194 32272 30200
rect 32036 29504 32088 29510
rect 32036 29446 32088 29452
rect 31944 28960 31996 28966
rect 31944 28902 31996 28908
rect 31852 28552 31904 28558
rect 31852 28494 31904 28500
rect 31864 28218 31892 28494
rect 31852 28212 31904 28218
rect 31852 28154 31904 28160
rect 31956 28150 31984 28902
rect 32048 28694 32076 29446
rect 32036 28688 32088 28694
rect 32036 28630 32088 28636
rect 32232 28218 32260 30194
rect 32324 28642 32352 33782
rect 32404 33516 32456 33522
rect 32404 33458 32456 33464
rect 32588 33516 32640 33522
rect 32588 33458 32640 33464
rect 32416 32842 32444 33458
rect 32404 32836 32456 32842
rect 32404 32778 32456 32784
rect 32416 32366 32444 32778
rect 32404 32360 32456 32366
rect 32404 32302 32456 32308
rect 32600 32026 32628 33458
rect 32956 33448 33008 33454
rect 32956 33390 33008 33396
rect 32680 33040 32732 33046
rect 32680 32982 32732 32988
rect 32692 32366 32720 32982
rect 32772 32904 32824 32910
rect 32772 32846 32824 32852
rect 32864 32904 32916 32910
rect 32864 32846 32916 32852
rect 32784 32570 32812 32846
rect 32772 32564 32824 32570
rect 32772 32506 32824 32512
rect 32680 32360 32732 32366
rect 32680 32302 32732 32308
rect 32588 32020 32640 32026
rect 32588 31962 32640 31968
rect 32692 31346 32720 32302
rect 32876 31482 32904 32846
rect 32968 32570 32996 33390
rect 33152 33114 33180 34002
rect 33324 33992 33376 33998
rect 33324 33934 33376 33940
rect 33232 33312 33284 33318
rect 33232 33254 33284 33260
rect 33140 33108 33192 33114
rect 33140 33050 33192 33056
rect 32956 32564 33008 32570
rect 32956 32506 33008 32512
rect 32956 31680 33008 31686
rect 32956 31622 33008 31628
rect 32864 31476 32916 31482
rect 32864 31418 32916 31424
rect 32680 31340 32732 31346
rect 32680 31282 32732 31288
rect 32772 31340 32824 31346
rect 32772 31282 32824 31288
rect 32692 30802 32720 31282
rect 32680 30796 32732 30802
rect 32680 30738 32732 30744
rect 32496 30660 32548 30666
rect 32496 30602 32548 30608
rect 32508 30258 32536 30602
rect 32784 30394 32812 31282
rect 32968 30734 32996 31622
rect 33140 31340 33192 31346
rect 33140 31282 33192 31288
rect 33152 30938 33180 31282
rect 33140 30932 33192 30938
rect 33140 30874 33192 30880
rect 33244 30802 33272 33254
rect 33336 32366 33364 33934
rect 33612 33658 33640 34546
rect 33692 34468 33744 34474
rect 33692 34410 33744 34416
rect 33704 33998 33732 34410
rect 33796 34202 33824 35022
rect 33784 34196 33836 34202
rect 33784 34138 33836 34144
rect 33692 33992 33744 33998
rect 33692 33934 33744 33940
rect 33784 33856 33836 33862
rect 33784 33798 33836 33804
rect 33600 33652 33652 33658
rect 33600 33594 33652 33600
rect 33796 33046 33824 33798
rect 33784 33040 33836 33046
rect 33784 32982 33836 32988
rect 33416 32836 33468 32842
rect 33416 32778 33468 32784
rect 33428 32502 33456 32778
rect 33416 32496 33468 32502
rect 33416 32438 33468 32444
rect 33784 32428 33836 32434
rect 33784 32370 33836 32376
rect 33324 32360 33376 32366
rect 33324 32302 33376 32308
rect 33324 31680 33376 31686
rect 33324 31622 33376 31628
rect 33336 31210 33364 31622
rect 33796 31414 33824 32370
rect 33888 31754 33916 35958
rect 33980 34542 34008 38247
rect 34072 37738 34100 41386
rect 34164 41206 34192 42230
rect 34256 41818 34284 42570
rect 34244 41812 34296 41818
rect 34244 41754 34296 41760
rect 34348 41698 34376 47194
rect 34808 46646 34836 49200
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 37200 47274 37228 49286
rect 38658 49200 38714 50000
rect 40590 49200 40646 50000
rect 42522 49314 42578 50000
rect 42522 49286 42748 49314
rect 42522 49200 42578 49286
rect 37372 47660 37424 47666
rect 37372 47602 37424 47608
rect 37200 47258 37320 47274
rect 37200 47252 37332 47258
rect 37200 47246 37280 47252
rect 37280 47194 37332 47200
rect 35900 46980 35952 46986
rect 35900 46922 35952 46928
rect 34796 46640 34848 46646
rect 34796 46582 34848 46588
rect 34704 46436 34756 46442
rect 34704 46378 34756 46384
rect 34428 46368 34480 46374
rect 34428 46310 34480 46316
rect 34440 44538 34468 46310
rect 34716 45937 34744 46378
rect 34808 46170 34836 46582
rect 35912 46374 35940 46922
rect 35900 46368 35952 46374
rect 35900 46310 35952 46316
rect 36820 46368 36872 46374
rect 36820 46310 36872 46316
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 34796 46164 34848 46170
rect 34796 46106 34848 46112
rect 34702 45928 34758 45937
rect 34702 45863 34758 45872
rect 34612 45484 34664 45490
rect 34612 45426 34664 45432
rect 34624 44810 34652 45426
rect 35532 45416 35584 45422
rect 35532 45358 35584 45364
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34704 44940 34756 44946
rect 34704 44882 34756 44888
rect 34612 44804 34664 44810
rect 34612 44746 34664 44752
rect 34716 44690 34744 44882
rect 34624 44662 34744 44690
rect 35440 44736 35492 44742
rect 35440 44678 35492 44684
rect 34428 44532 34480 44538
rect 34428 44474 34480 44480
rect 34624 43790 34652 44662
rect 35452 44402 35480 44678
rect 35544 44402 35572 45358
rect 36084 44736 36136 44742
rect 36084 44678 36136 44684
rect 34704 44396 34756 44402
rect 34704 44338 34756 44344
rect 35440 44396 35492 44402
rect 35440 44338 35492 44344
rect 35532 44396 35584 44402
rect 35532 44338 35584 44344
rect 34612 43784 34664 43790
rect 34612 43726 34664 43732
rect 34520 43444 34572 43450
rect 34520 43386 34572 43392
rect 34428 42764 34480 42770
rect 34428 42706 34480 42712
rect 34256 41670 34376 41698
rect 34152 41200 34204 41206
rect 34152 41142 34204 41148
rect 34152 40928 34204 40934
rect 34152 40870 34204 40876
rect 34164 40730 34192 40870
rect 34152 40724 34204 40730
rect 34152 40666 34204 40672
rect 34152 40452 34204 40458
rect 34152 40394 34204 40400
rect 34164 40361 34192 40394
rect 34150 40352 34206 40361
rect 34150 40287 34206 40296
rect 34152 38956 34204 38962
rect 34152 38898 34204 38904
rect 34060 37732 34112 37738
rect 34060 37674 34112 37680
rect 34060 37324 34112 37330
rect 34060 37266 34112 37272
rect 34072 35766 34100 37266
rect 34164 37194 34192 38898
rect 34256 38894 34284 41670
rect 34336 41540 34388 41546
rect 34336 41482 34388 41488
rect 34348 40594 34376 41482
rect 34440 40662 34468 42706
rect 34532 41750 34560 43386
rect 34624 42838 34652 43726
rect 34612 42832 34664 42838
rect 34612 42774 34664 42780
rect 34716 42770 34744 44338
rect 34796 44328 34848 44334
rect 34796 44270 34848 44276
rect 34808 43994 34836 44270
rect 35348 44192 35400 44198
rect 35348 44134 35400 44140
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 34796 43988 34848 43994
rect 34796 43930 34848 43936
rect 35360 43858 35388 44134
rect 35348 43852 35400 43858
rect 35348 43794 35400 43800
rect 35164 43784 35216 43790
rect 35164 43726 35216 43732
rect 35176 43110 35204 43726
rect 35544 43722 35572 44338
rect 35900 44260 35952 44266
rect 35900 44202 35952 44208
rect 35624 43784 35676 43790
rect 35624 43726 35676 43732
rect 35532 43716 35584 43722
rect 35532 43658 35584 43664
rect 35544 43382 35572 43658
rect 35532 43376 35584 43382
rect 35532 43318 35584 43324
rect 35164 43104 35216 43110
rect 35164 43046 35216 43052
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 35438 42800 35494 42809
rect 34704 42764 34756 42770
rect 35438 42735 35494 42744
rect 34704 42706 34756 42712
rect 35452 42702 35480 42735
rect 35164 42696 35216 42702
rect 35164 42638 35216 42644
rect 35440 42696 35492 42702
rect 35440 42638 35492 42644
rect 35176 42022 35204 42638
rect 35348 42628 35400 42634
rect 35348 42570 35400 42576
rect 35360 42362 35388 42570
rect 35348 42356 35400 42362
rect 35348 42298 35400 42304
rect 35348 42220 35400 42226
rect 35348 42162 35400 42168
rect 35164 42016 35216 42022
rect 35164 41958 35216 41964
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 35360 41818 35388 42162
rect 35452 42158 35480 42638
rect 35544 42362 35572 43318
rect 35636 43314 35664 43726
rect 35912 43450 35940 44202
rect 35992 43716 36044 43722
rect 35992 43658 36044 43664
rect 35900 43444 35952 43450
rect 35900 43386 35952 43392
rect 35624 43308 35676 43314
rect 35624 43250 35676 43256
rect 35636 42566 35664 43250
rect 36004 43246 36032 43658
rect 35992 43240 36044 43246
rect 35992 43182 36044 43188
rect 35900 43172 35952 43178
rect 35900 43114 35952 43120
rect 35912 42566 35940 43114
rect 36004 42702 36032 43182
rect 36096 42809 36124 44678
rect 36728 44192 36780 44198
rect 36728 44134 36780 44140
rect 36188 43858 36492 43874
rect 36176 43852 36492 43858
rect 36228 43846 36492 43852
rect 36176 43794 36228 43800
rect 36268 43784 36320 43790
rect 36268 43726 36320 43732
rect 36082 42800 36138 42809
rect 36082 42735 36138 42744
rect 36280 42702 36308 43726
rect 36464 43722 36492 43846
rect 36452 43716 36504 43722
rect 36452 43658 36504 43664
rect 36636 43716 36688 43722
rect 36636 43658 36688 43664
rect 35992 42696 36044 42702
rect 35992 42638 36044 42644
rect 36268 42696 36320 42702
rect 36268 42638 36320 42644
rect 35624 42560 35676 42566
rect 35624 42502 35676 42508
rect 35900 42560 35952 42566
rect 35900 42502 35952 42508
rect 36004 42362 36032 42638
rect 36464 42566 36492 43658
rect 36648 43178 36676 43658
rect 36740 43246 36768 44134
rect 36728 43240 36780 43246
rect 36728 43182 36780 43188
rect 36636 43172 36688 43178
rect 36636 43114 36688 43120
rect 36452 42560 36504 42566
rect 36452 42502 36504 42508
rect 36544 42560 36596 42566
rect 36544 42502 36596 42508
rect 35532 42356 35584 42362
rect 35532 42298 35584 42304
rect 35992 42356 36044 42362
rect 35992 42298 36044 42304
rect 35440 42152 35492 42158
rect 35440 42094 35492 42100
rect 36360 42152 36412 42158
rect 36360 42094 36412 42100
rect 35808 42016 35860 42022
rect 35808 41958 35860 41964
rect 35348 41812 35400 41818
rect 35348 41754 35400 41760
rect 34520 41744 34572 41750
rect 34520 41686 34572 41692
rect 34888 41744 34940 41750
rect 34888 41686 34940 41692
rect 34612 41472 34664 41478
rect 34612 41414 34664 41420
rect 34520 41064 34572 41070
rect 34520 41006 34572 41012
rect 34428 40656 34480 40662
rect 34428 40598 34480 40604
rect 34336 40588 34388 40594
rect 34336 40530 34388 40536
rect 34532 40066 34560 41006
rect 34336 40044 34388 40050
rect 34336 39986 34388 39992
rect 34440 40038 34560 40066
rect 34348 39642 34376 39986
rect 34336 39636 34388 39642
rect 34336 39578 34388 39584
rect 34336 39432 34388 39438
rect 34336 39374 34388 39380
rect 34348 39273 34376 39374
rect 34334 39264 34390 39273
rect 34334 39199 34390 39208
rect 34440 39030 34468 40038
rect 34520 39976 34572 39982
rect 34520 39918 34572 39924
rect 34532 39846 34560 39918
rect 34520 39840 34572 39846
rect 34520 39782 34572 39788
rect 34428 39024 34480 39030
rect 34428 38966 34480 38972
rect 34244 38888 34296 38894
rect 34244 38830 34296 38836
rect 34336 38752 34388 38758
rect 34336 38694 34388 38700
rect 34242 38584 34298 38593
rect 34242 38519 34298 38528
rect 34256 37262 34284 38519
rect 34348 37942 34376 38694
rect 34532 38049 34560 39782
rect 34518 38040 34574 38049
rect 34518 37975 34574 37984
rect 34336 37936 34388 37942
rect 34336 37878 34388 37884
rect 34520 37868 34572 37874
rect 34520 37810 34572 37816
rect 34336 37324 34388 37330
rect 34336 37266 34388 37272
rect 34244 37256 34296 37262
rect 34244 37198 34296 37204
rect 34152 37188 34204 37194
rect 34152 37130 34204 37136
rect 34256 37074 34284 37198
rect 34164 37046 34284 37074
rect 34164 36553 34192 37046
rect 34242 36952 34298 36961
rect 34242 36887 34298 36896
rect 34256 36582 34284 36887
rect 34244 36576 34296 36582
rect 34150 36544 34206 36553
rect 34244 36518 34296 36524
rect 34150 36479 34206 36488
rect 34164 35873 34192 36479
rect 34150 35864 34206 35873
rect 34150 35799 34206 35808
rect 34060 35760 34112 35766
rect 34060 35702 34112 35708
rect 34244 35692 34296 35698
rect 34244 35634 34296 35640
rect 34152 35148 34204 35154
rect 34152 35090 34204 35096
rect 34164 34746 34192 35090
rect 34152 34740 34204 34746
rect 34152 34682 34204 34688
rect 34256 34542 34284 35634
rect 33968 34536 34020 34542
rect 33968 34478 34020 34484
rect 34244 34536 34296 34542
rect 34244 34478 34296 34484
rect 33968 34400 34020 34406
rect 33968 34342 34020 34348
rect 33980 33998 34008 34342
rect 33968 33992 34020 33998
rect 33968 33934 34020 33940
rect 33980 33862 34008 33934
rect 33968 33856 34020 33862
rect 33968 33798 34020 33804
rect 33980 32570 34008 33798
rect 34060 33108 34112 33114
rect 34060 33050 34112 33056
rect 33968 32564 34020 32570
rect 33968 32506 34020 32512
rect 34072 32434 34100 33050
rect 34060 32428 34112 32434
rect 34060 32370 34112 32376
rect 33968 32224 34020 32230
rect 33968 32166 34020 32172
rect 33980 31890 34008 32166
rect 34072 32026 34100 32370
rect 34060 32020 34112 32026
rect 34060 31962 34112 31968
rect 33968 31884 34020 31890
rect 33968 31826 34020 31832
rect 33888 31726 34192 31754
rect 33784 31408 33836 31414
rect 33784 31350 33836 31356
rect 33416 31340 33468 31346
rect 33416 31282 33468 31288
rect 33324 31204 33376 31210
rect 33324 31146 33376 31152
rect 33232 30796 33284 30802
rect 33232 30738 33284 30744
rect 32956 30728 33008 30734
rect 32956 30670 33008 30676
rect 32772 30388 32824 30394
rect 32772 30330 32824 30336
rect 32968 30326 32996 30670
rect 33244 30598 33272 30738
rect 33428 30716 33456 31282
rect 34164 31278 34192 31726
rect 34152 31272 34204 31278
rect 34152 31214 34204 31220
rect 33508 30728 33560 30734
rect 33428 30688 33508 30716
rect 33508 30670 33560 30676
rect 33232 30592 33284 30598
rect 33232 30534 33284 30540
rect 32956 30320 33008 30326
rect 32956 30262 33008 30268
rect 32496 30252 32548 30258
rect 32496 30194 32548 30200
rect 33140 30252 33192 30258
rect 33140 30194 33192 30200
rect 33152 29714 33180 30194
rect 33140 29708 33192 29714
rect 33140 29650 33192 29656
rect 32496 29640 32548 29646
rect 32496 29582 32548 29588
rect 32680 29640 32732 29646
rect 32680 29582 32732 29588
rect 32508 29238 32536 29582
rect 32496 29232 32548 29238
rect 32496 29174 32548 29180
rect 32692 29170 32720 29582
rect 33152 29306 33180 29650
rect 33140 29300 33192 29306
rect 33140 29242 33192 29248
rect 32680 29164 32732 29170
rect 32680 29106 32732 29112
rect 32324 28614 32444 28642
rect 32312 28484 32364 28490
rect 32312 28426 32364 28432
rect 32220 28212 32272 28218
rect 32220 28154 32272 28160
rect 31944 28144 31996 28150
rect 31944 28086 31996 28092
rect 32128 28144 32180 28150
rect 32128 28086 32180 28092
rect 32140 27470 32168 28086
rect 32128 27464 32180 27470
rect 32128 27406 32180 27412
rect 32036 27396 32088 27402
rect 32036 27338 32088 27344
rect 32048 27130 32076 27338
rect 32324 27334 32352 28426
rect 32312 27328 32364 27334
rect 32312 27270 32364 27276
rect 32324 27130 32352 27270
rect 32036 27124 32088 27130
rect 32036 27066 32088 27072
rect 32312 27124 32364 27130
rect 32312 27066 32364 27072
rect 32036 26920 32088 26926
rect 32036 26862 32088 26868
rect 32048 25702 32076 26862
rect 32036 25696 32088 25702
rect 32036 25638 32088 25644
rect 31668 10056 31720 10062
rect 31668 9998 31720 10004
rect 31116 9920 31168 9926
rect 31116 9862 31168 9868
rect 28448 2508 28500 2514
rect 28448 2450 28500 2456
rect 30656 2508 30708 2514
rect 30656 2450 30708 2456
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 28356 2372 28408 2378
rect 28356 2314 28408 2320
rect 27160 2032 27212 2038
rect 27160 1974 27212 1980
rect 28368 800 28396 2314
rect 30300 800 30328 2382
rect 32048 2106 32076 25638
rect 32416 22094 32444 28614
rect 32496 28552 32548 28558
rect 32496 28494 32548 28500
rect 32508 28218 32536 28494
rect 32496 28212 32548 28218
rect 32496 28154 32548 28160
rect 32508 27470 32536 28154
rect 32864 28076 32916 28082
rect 32864 28018 32916 28024
rect 32876 27674 32904 28018
rect 32864 27668 32916 27674
rect 32864 27610 32916 27616
rect 32496 27464 32548 27470
rect 32496 27406 32548 27412
rect 32772 27056 32824 27062
rect 32772 26998 32824 27004
rect 32784 26926 32812 26998
rect 33048 26988 33100 26994
rect 33048 26930 33100 26936
rect 32772 26920 32824 26926
rect 32772 26862 32824 26868
rect 32784 26042 32812 26862
rect 33060 26586 33088 26930
rect 33048 26580 33100 26586
rect 33048 26522 33100 26528
rect 33244 26382 33272 30534
rect 33324 30048 33376 30054
rect 33324 29990 33376 29996
rect 33336 29782 33364 29990
rect 33520 29850 33548 30670
rect 34060 30592 34112 30598
rect 34060 30534 34112 30540
rect 34072 30258 34100 30534
rect 33600 30252 33652 30258
rect 33600 30194 33652 30200
rect 34060 30252 34112 30258
rect 34060 30194 34112 30200
rect 33508 29844 33560 29850
rect 33508 29786 33560 29792
rect 33324 29776 33376 29782
rect 33324 29718 33376 29724
rect 33612 29646 33640 30194
rect 34164 30190 34192 31214
rect 34152 30184 34204 30190
rect 34152 30126 34204 30132
rect 33692 30048 33744 30054
rect 33692 29990 33744 29996
rect 33704 29646 33732 29990
rect 34256 29850 34284 34478
rect 34348 33386 34376 37266
rect 34532 36825 34560 37810
rect 34518 36816 34574 36825
rect 34518 36751 34520 36760
rect 34572 36751 34574 36760
rect 34520 36722 34572 36728
rect 34428 36576 34480 36582
rect 34428 36518 34480 36524
rect 34440 35698 34468 36518
rect 34624 36378 34652 41414
rect 34704 41132 34756 41138
rect 34704 41074 34756 41080
rect 34716 40526 34744 41074
rect 34900 41070 34928 41686
rect 35716 41608 35768 41614
rect 35636 41556 35716 41562
rect 35636 41550 35768 41556
rect 35636 41534 35756 41550
rect 34888 41064 34940 41070
rect 34888 41006 34940 41012
rect 35348 40996 35400 41002
rect 35348 40938 35400 40944
rect 34796 40928 34848 40934
rect 34796 40870 34848 40876
rect 34704 40520 34756 40526
rect 34704 40462 34756 40468
rect 34704 40384 34756 40390
rect 34704 40326 34756 40332
rect 34716 37233 34744 40326
rect 34808 39488 34836 40870
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 35360 40526 35388 40938
rect 35348 40520 35400 40526
rect 35348 40462 35400 40468
rect 35532 40520 35584 40526
rect 35532 40462 35584 40468
rect 35348 40384 35400 40390
rect 35348 40326 35400 40332
rect 35440 40384 35492 40390
rect 35440 40326 35492 40332
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34980 39500 35032 39506
rect 34808 39460 34980 39488
rect 34980 39442 35032 39448
rect 35360 39438 35388 40326
rect 35452 40118 35480 40326
rect 35544 40186 35572 40462
rect 35532 40180 35584 40186
rect 35532 40122 35584 40128
rect 35440 40112 35492 40118
rect 35440 40054 35492 40060
rect 35530 40080 35586 40089
rect 35530 40015 35586 40024
rect 35440 39976 35492 39982
rect 35440 39918 35492 39924
rect 35452 39574 35480 39918
rect 35440 39568 35492 39574
rect 35440 39510 35492 39516
rect 35544 39438 35572 40015
rect 35348 39432 35400 39438
rect 35348 39374 35400 39380
rect 35532 39432 35584 39438
rect 35532 39374 35584 39380
rect 35348 39296 35400 39302
rect 34794 39264 34850 39273
rect 35348 39238 35400 39244
rect 34794 39199 34850 39208
rect 34808 38593 34836 39199
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34794 38584 34850 38593
rect 34934 38587 35242 38596
rect 34794 38519 34850 38528
rect 34808 38406 35020 38434
rect 35360 38418 35388 39238
rect 35440 38752 35492 38758
rect 35438 38720 35440 38729
rect 35492 38720 35494 38729
rect 35438 38655 35494 38664
rect 35438 38584 35494 38593
rect 35438 38519 35494 38528
rect 34808 38214 34836 38406
rect 34888 38276 34940 38282
rect 34888 38218 34940 38224
rect 34796 38208 34848 38214
rect 34796 38150 34848 38156
rect 34900 38010 34928 38218
rect 34992 38214 35020 38406
rect 35072 38412 35124 38418
rect 35072 38354 35124 38360
rect 35348 38412 35400 38418
rect 35348 38354 35400 38360
rect 35084 38321 35112 38354
rect 35070 38312 35126 38321
rect 35070 38247 35126 38256
rect 35348 38276 35400 38282
rect 35348 38218 35400 38224
rect 34980 38208 35032 38214
rect 34980 38150 35032 38156
rect 34888 38004 34940 38010
rect 34888 37946 34940 37952
rect 34794 37904 34850 37913
rect 34794 37839 34850 37848
rect 34702 37224 34758 37233
rect 34702 37159 34758 37168
rect 34716 37126 34744 37159
rect 34704 37120 34756 37126
rect 34704 37062 34756 37068
rect 34704 36644 34756 36650
rect 34704 36586 34756 36592
rect 34612 36372 34664 36378
rect 34612 36314 34664 36320
rect 34716 36242 34744 36586
rect 34808 36242 34836 37839
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35360 37466 35388 38218
rect 35348 37460 35400 37466
rect 35348 37402 35400 37408
rect 35452 36786 35480 38519
rect 35532 37936 35584 37942
rect 35532 37878 35584 37884
rect 35544 36854 35572 37878
rect 35636 37210 35664 41534
rect 35820 41426 35848 41958
rect 36372 41818 36400 42094
rect 36556 41834 36584 42502
rect 36360 41812 36412 41818
rect 36360 41754 36412 41760
rect 36464 41806 36584 41834
rect 36176 41744 36228 41750
rect 36176 41686 36228 41692
rect 35728 41398 35848 41426
rect 35728 39846 35756 41398
rect 35808 41132 35860 41138
rect 35808 41074 35860 41080
rect 35820 40934 35848 41074
rect 36188 41070 36216 41686
rect 36268 41200 36320 41206
rect 36268 41142 36320 41148
rect 35900 41064 35952 41070
rect 36084 41064 36136 41070
rect 35952 41024 36032 41052
rect 35900 41006 35952 41012
rect 35808 40928 35860 40934
rect 35808 40870 35860 40876
rect 35900 40928 35952 40934
rect 35900 40870 35952 40876
rect 35820 40594 35848 40870
rect 35808 40588 35860 40594
rect 35808 40530 35860 40536
rect 35820 39982 35848 40530
rect 35912 40526 35940 40870
rect 36004 40730 36032 41024
rect 36084 41006 36136 41012
rect 36176 41064 36228 41070
rect 36176 41006 36228 41012
rect 35992 40724 36044 40730
rect 35992 40666 36044 40672
rect 35900 40520 35952 40526
rect 35900 40462 35952 40468
rect 36004 40186 36032 40666
rect 35992 40180 36044 40186
rect 35992 40122 36044 40128
rect 35900 40044 35952 40050
rect 35900 39986 35952 39992
rect 35808 39976 35860 39982
rect 35808 39918 35860 39924
rect 35716 39840 35768 39846
rect 35716 39782 35768 39788
rect 35912 39642 35940 39986
rect 36004 39642 36032 40122
rect 36096 39914 36124 41006
rect 36176 40656 36228 40662
rect 36176 40598 36228 40604
rect 36188 40458 36216 40598
rect 36176 40452 36228 40458
rect 36176 40394 36228 40400
rect 36084 39908 36136 39914
rect 36084 39850 36136 39856
rect 35900 39636 35952 39642
rect 35900 39578 35952 39584
rect 35992 39636 36044 39642
rect 35992 39578 36044 39584
rect 36280 39506 36308 41142
rect 36360 40044 36412 40050
rect 36360 39986 36412 39992
rect 36372 39642 36400 39986
rect 36360 39636 36412 39642
rect 36360 39578 36412 39584
rect 36268 39500 36320 39506
rect 36268 39442 36320 39448
rect 36372 39438 36400 39578
rect 36360 39432 36412 39438
rect 36360 39374 36412 39380
rect 36464 39114 36492 41806
rect 36544 41676 36596 41682
rect 36544 41618 36596 41624
rect 36556 41274 36584 41618
rect 36544 41268 36596 41274
rect 36544 41210 36596 41216
rect 36636 40588 36688 40594
rect 36636 40530 36688 40536
rect 36544 40044 36596 40050
rect 36544 39986 36596 39992
rect 36556 39438 36584 39986
rect 36648 39982 36676 40530
rect 36636 39976 36688 39982
rect 36636 39918 36688 39924
rect 36740 39574 36768 43182
rect 36728 39568 36780 39574
rect 36728 39510 36780 39516
rect 36544 39432 36596 39438
rect 36542 39400 36544 39409
rect 36596 39400 36598 39409
rect 36542 39335 36598 39344
rect 36464 39086 36584 39114
rect 36176 38956 36228 38962
rect 36176 38898 36228 38904
rect 36452 38956 36504 38962
rect 36452 38898 36504 38904
rect 35716 38888 35768 38894
rect 35716 38830 35768 38836
rect 35728 38758 35756 38830
rect 35716 38752 35768 38758
rect 35716 38694 35768 38700
rect 35728 38593 35756 38694
rect 35714 38584 35770 38593
rect 35714 38519 35770 38528
rect 35716 38412 35768 38418
rect 35716 38354 35768 38360
rect 35728 38010 35756 38354
rect 36084 38344 36136 38350
rect 36082 38312 36084 38321
rect 36136 38312 36138 38321
rect 36082 38247 36138 38256
rect 35808 38208 35860 38214
rect 35808 38150 35860 38156
rect 35716 38004 35768 38010
rect 35716 37946 35768 37952
rect 35820 37262 35848 38150
rect 36188 37874 36216 38898
rect 36268 38752 36320 38758
rect 36268 38694 36320 38700
rect 36280 38350 36308 38694
rect 36360 38480 36412 38486
rect 36358 38448 36360 38457
rect 36412 38448 36414 38457
rect 36358 38383 36414 38392
rect 36268 38344 36320 38350
rect 36268 38286 36320 38292
rect 36280 37874 36308 38286
rect 36176 37868 36228 37874
rect 36176 37810 36228 37816
rect 36268 37868 36320 37874
rect 36268 37810 36320 37816
rect 35992 37800 36044 37806
rect 35992 37742 36044 37748
rect 35808 37256 35860 37262
rect 35636 37182 35756 37210
rect 35808 37198 35860 37204
rect 35624 37120 35676 37126
rect 35624 37062 35676 37068
rect 35532 36848 35584 36854
rect 35532 36790 35584 36796
rect 35440 36780 35492 36786
rect 35440 36722 35492 36728
rect 35348 36576 35400 36582
rect 35348 36518 35400 36524
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34704 36236 34756 36242
rect 34704 36178 34756 36184
rect 34796 36236 34848 36242
rect 34796 36178 34848 36184
rect 34428 35692 34480 35698
rect 34428 35634 34480 35640
rect 34716 35154 34744 36178
rect 34796 35488 34848 35494
rect 34796 35430 34848 35436
rect 34704 35148 34756 35154
rect 34704 35090 34756 35096
rect 34520 34944 34572 34950
rect 34808 34921 34836 35430
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34888 35080 34940 35086
rect 34888 35022 34940 35028
rect 34520 34886 34572 34892
rect 34794 34912 34850 34921
rect 34428 34196 34480 34202
rect 34428 34138 34480 34144
rect 34336 33380 34388 33386
rect 34336 33322 34388 33328
rect 34440 33318 34468 34138
rect 34532 33590 34560 34886
rect 34794 34847 34850 34856
rect 34900 34388 34928 35022
rect 34808 34360 34928 34388
rect 34520 33584 34572 33590
rect 34520 33526 34572 33532
rect 34520 33448 34572 33454
rect 34520 33390 34572 33396
rect 34428 33312 34480 33318
rect 34428 33254 34480 33260
rect 34532 32230 34560 33390
rect 34808 32910 34836 34360
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35360 34066 35388 36518
rect 35544 35834 35572 36790
rect 35636 36378 35664 37062
rect 35624 36372 35676 36378
rect 35624 36314 35676 36320
rect 35532 35828 35584 35834
rect 35532 35770 35584 35776
rect 35530 35184 35586 35193
rect 35530 35119 35586 35128
rect 35544 34610 35572 35119
rect 35532 34604 35584 34610
rect 35532 34546 35584 34552
rect 35440 34536 35492 34542
rect 35440 34478 35492 34484
rect 35452 34202 35480 34478
rect 35728 34474 35756 37182
rect 35808 37120 35860 37126
rect 35808 37062 35860 37068
rect 35820 36786 35848 37062
rect 36004 36786 36032 37742
rect 36464 37262 36492 38898
rect 36556 37806 36584 39086
rect 36832 38654 36860 46310
rect 37384 45554 37412 47602
rect 38672 47258 38700 49200
rect 40604 47258 40632 49200
rect 42720 48090 42748 49286
rect 44454 49200 44510 50000
rect 46386 49314 46442 50000
rect 46386 49286 46704 49314
rect 46386 49200 46442 49286
rect 42720 48062 42840 48090
rect 40776 47456 40828 47462
rect 40776 47398 40828 47404
rect 40788 47258 40816 47398
rect 42812 47258 42840 48062
rect 38660 47252 38712 47258
rect 38660 47194 38712 47200
rect 40592 47252 40644 47258
rect 40592 47194 40644 47200
rect 40776 47252 40828 47258
rect 40776 47194 40828 47200
rect 42800 47252 42852 47258
rect 42800 47194 42852 47200
rect 38672 47054 38700 47194
rect 40604 47054 40632 47194
rect 42432 47116 42484 47122
rect 42432 47058 42484 47064
rect 38660 47048 38712 47054
rect 38660 46990 38712 46996
rect 40592 47048 40644 47054
rect 40592 46990 40644 46996
rect 38752 46912 38804 46918
rect 38752 46854 38804 46860
rect 38764 45626 38792 46854
rect 42444 46714 42472 47058
rect 44468 46918 44496 49200
rect 46676 47258 46704 49286
rect 48318 49200 48374 50000
rect 49606 49200 49662 50000
rect 48042 48376 48098 48385
rect 48042 48311 48098 48320
rect 46664 47252 46716 47258
rect 46664 47194 46716 47200
rect 46204 47048 46256 47054
rect 46204 46990 46256 46996
rect 45468 46980 45520 46986
rect 45468 46922 45520 46928
rect 44456 46912 44508 46918
rect 44456 46854 44508 46860
rect 45192 46912 45244 46918
rect 45192 46854 45244 46860
rect 45204 46714 45232 46854
rect 42432 46708 42484 46714
rect 42432 46650 42484 46656
rect 45192 46708 45244 46714
rect 45192 46650 45244 46656
rect 43260 46504 43312 46510
rect 43260 46446 43312 46452
rect 38752 45620 38804 45626
rect 38752 45562 38804 45568
rect 37292 45526 37412 45554
rect 37292 44198 37320 45526
rect 43272 45354 43300 46446
rect 43260 45348 43312 45354
rect 43260 45290 43312 45296
rect 37280 44192 37332 44198
rect 37280 44134 37332 44140
rect 37740 44192 37792 44198
rect 37740 44134 37792 44140
rect 37924 44192 37976 44198
rect 37924 44134 37976 44140
rect 37752 43722 37780 44134
rect 37936 43790 37964 44134
rect 37924 43784 37976 43790
rect 37924 43726 37976 43732
rect 37740 43716 37792 43722
rect 37740 43658 37792 43664
rect 37832 43648 37884 43654
rect 37832 43590 37884 43596
rect 38384 43648 38436 43654
rect 38384 43590 38436 43596
rect 38568 43648 38620 43654
rect 38568 43590 38620 43596
rect 37844 43314 37872 43590
rect 38396 43314 38424 43590
rect 38580 43314 38608 43590
rect 37832 43308 37884 43314
rect 37832 43250 37884 43256
rect 38292 43308 38344 43314
rect 38292 43250 38344 43256
rect 38384 43308 38436 43314
rect 38384 43250 38436 43256
rect 38568 43308 38620 43314
rect 38568 43250 38620 43256
rect 38304 43110 38332 43250
rect 38016 43104 38068 43110
rect 38016 43046 38068 43052
rect 38292 43104 38344 43110
rect 38292 43046 38344 43052
rect 37280 42764 37332 42770
rect 37280 42706 37332 42712
rect 37292 42673 37320 42706
rect 38028 42702 38056 43046
rect 38304 42770 38332 43046
rect 38292 42764 38344 42770
rect 38292 42706 38344 42712
rect 37464 42696 37516 42702
rect 37278 42664 37334 42673
rect 37188 42628 37240 42634
rect 37464 42638 37516 42644
rect 38016 42696 38068 42702
rect 38016 42638 38068 42644
rect 37278 42599 37334 42608
rect 37188 42570 37240 42576
rect 37200 42090 37228 42570
rect 37292 42158 37320 42599
rect 37476 42226 37504 42638
rect 37740 42560 37792 42566
rect 37740 42502 37792 42508
rect 37464 42220 37516 42226
rect 37464 42162 37516 42168
rect 37280 42152 37332 42158
rect 37280 42094 37332 42100
rect 37188 42084 37240 42090
rect 37188 42026 37240 42032
rect 37648 42084 37700 42090
rect 37648 42026 37700 42032
rect 37660 41614 37688 42026
rect 37752 41682 37780 42502
rect 38292 42220 38344 42226
rect 38292 42162 38344 42168
rect 37924 42016 37976 42022
rect 37924 41958 37976 41964
rect 37740 41676 37792 41682
rect 37740 41618 37792 41624
rect 37648 41608 37700 41614
rect 37648 41550 37700 41556
rect 37004 41472 37056 41478
rect 37004 41414 37056 41420
rect 36912 40452 36964 40458
rect 36912 40394 36964 40400
rect 36924 40186 36952 40394
rect 36912 40180 36964 40186
rect 36912 40122 36964 40128
rect 37016 39370 37044 41414
rect 37740 41132 37792 41138
rect 37740 41074 37792 41080
rect 37832 41132 37884 41138
rect 37832 41074 37884 41080
rect 37280 40928 37332 40934
rect 37280 40870 37332 40876
rect 37096 40724 37148 40730
rect 37096 40666 37148 40672
rect 37108 40458 37136 40666
rect 37096 40452 37148 40458
rect 37096 40394 37148 40400
rect 37292 39953 37320 40870
rect 37752 40730 37780 41074
rect 37844 41002 37872 41074
rect 37832 40996 37884 41002
rect 37832 40938 37884 40944
rect 37740 40724 37792 40730
rect 37740 40666 37792 40672
rect 37844 40610 37872 40938
rect 37752 40582 37872 40610
rect 37464 40384 37516 40390
rect 37464 40326 37516 40332
rect 37476 40050 37504 40326
rect 37464 40044 37516 40050
rect 37464 39986 37516 39992
rect 37372 39976 37424 39982
rect 37278 39944 37334 39953
rect 37372 39918 37424 39924
rect 37278 39879 37334 39888
rect 37004 39364 37056 39370
rect 37004 39306 37056 39312
rect 36740 38626 36860 38654
rect 36544 37800 36596 37806
rect 36544 37742 36596 37748
rect 36636 37460 36688 37466
rect 36636 37402 36688 37408
rect 36452 37256 36504 37262
rect 36452 37198 36504 37204
rect 36268 37188 36320 37194
rect 36268 37130 36320 37136
rect 35808 36780 35860 36786
rect 35808 36722 35860 36728
rect 35992 36780 36044 36786
rect 35992 36722 36044 36728
rect 35820 36106 35848 36722
rect 36280 36174 36308 37130
rect 36648 36718 36676 37402
rect 36740 37330 36768 38626
rect 37384 38418 37412 39918
rect 37464 39840 37516 39846
rect 37464 39782 37516 39788
rect 37372 38412 37424 38418
rect 37372 38354 37424 38360
rect 37384 37738 37412 38354
rect 37476 38010 37504 39782
rect 37648 39364 37700 39370
rect 37648 39306 37700 39312
rect 37660 39098 37688 39306
rect 37648 39092 37700 39098
rect 37648 39034 37700 39040
rect 37554 38992 37610 39001
rect 37554 38927 37610 38936
rect 37464 38004 37516 38010
rect 37464 37946 37516 37952
rect 37464 37868 37516 37874
rect 37464 37810 37516 37816
rect 37372 37732 37424 37738
rect 37372 37674 37424 37680
rect 37372 37392 37424 37398
rect 37370 37360 37372 37369
rect 37424 37360 37426 37369
rect 36728 37324 36780 37330
rect 36728 37266 36780 37272
rect 37280 37324 37332 37330
rect 37370 37295 37426 37304
rect 37280 37266 37332 37272
rect 37096 37188 37148 37194
rect 37096 37130 37148 37136
rect 36636 36712 36688 36718
rect 36636 36654 36688 36660
rect 36648 36174 36676 36654
rect 36268 36168 36320 36174
rect 36268 36110 36320 36116
rect 36636 36168 36688 36174
rect 36636 36110 36688 36116
rect 37004 36168 37056 36174
rect 37004 36110 37056 36116
rect 35808 36100 35860 36106
rect 35808 36042 35860 36048
rect 36280 35834 36308 36110
rect 36452 36100 36504 36106
rect 36452 36042 36504 36048
rect 36268 35828 36320 35834
rect 36268 35770 36320 35776
rect 36464 35698 36492 36042
rect 37016 35698 37044 36110
rect 36452 35692 36504 35698
rect 36452 35634 36504 35640
rect 36544 35692 36596 35698
rect 36544 35634 36596 35640
rect 37004 35692 37056 35698
rect 37004 35634 37056 35640
rect 36556 35222 36584 35634
rect 36544 35216 36596 35222
rect 36544 35158 36596 35164
rect 36268 35148 36320 35154
rect 36268 35090 36320 35096
rect 36280 34746 36308 35090
rect 37004 34944 37056 34950
rect 37004 34886 37056 34892
rect 36268 34740 36320 34746
rect 36268 34682 36320 34688
rect 35900 34672 35952 34678
rect 35900 34614 35952 34620
rect 36728 34672 36780 34678
rect 37016 34649 37044 34886
rect 36728 34614 36780 34620
rect 37002 34640 37058 34649
rect 35716 34468 35768 34474
rect 35716 34410 35768 34416
rect 35440 34196 35492 34202
rect 35440 34138 35492 34144
rect 35348 34060 35400 34066
rect 35348 34002 35400 34008
rect 35532 34060 35584 34066
rect 35532 34002 35584 34008
rect 35544 33590 35572 34002
rect 35808 33992 35860 33998
rect 35808 33934 35860 33940
rect 35532 33584 35584 33590
rect 35532 33526 35584 33532
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34796 32904 34848 32910
rect 34796 32846 34848 32852
rect 34980 32904 35032 32910
rect 34980 32846 35032 32852
rect 34704 32768 34756 32774
rect 34704 32710 34756 32716
rect 34716 32502 34744 32710
rect 34704 32496 34756 32502
rect 34704 32438 34756 32444
rect 34520 32224 34572 32230
rect 34520 32166 34572 32172
rect 34716 31890 34744 32438
rect 34796 32428 34848 32434
rect 34796 32370 34848 32376
rect 34808 32026 34836 32370
rect 34992 32366 35020 32846
rect 35348 32564 35400 32570
rect 35348 32506 35400 32512
rect 34980 32360 35032 32366
rect 34980 32302 35032 32308
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34796 32020 34848 32026
rect 34796 31962 34848 31968
rect 34704 31884 34756 31890
rect 34704 31826 34756 31832
rect 34520 31816 34572 31822
rect 34520 31758 34572 31764
rect 34532 31482 34560 31758
rect 35360 31754 35388 32506
rect 35440 32428 35492 32434
rect 35440 32370 35492 32376
rect 35452 31958 35480 32370
rect 35440 31952 35492 31958
rect 35440 31894 35492 31900
rect 35348 31748 35400 31754
rect 35348 31690 35400 31696
rect 34520 31476 34572 31482
rect 34520 31418 34572 31424
rect 35360 31414 35388 31690
rect 35348 31408 35400 31414
rect 35348 31350 35400 31356
rect 35452 31278 35480 31894
rect 35544 31482 35572 33526
rect 35624 33448 35676 33454
rect 35624 33390 35676 33396
rect 35532 31476 35584 31482
rect 35532 31418 35584 31424
rect 35440 31272 35492 31278
rect 35440 31214 35492 31220
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34704 30660 34756 30666
rect 34704 30602 34756 30608
rect 34716 30258 34744 30602
rect 34704 30252 34756 30258
rect 34704 30194 34756 30200
rect 35256 30252 35308 30258
rect 35256 30194 35308 30200
rect 34796 30184 34848 30190
rect 34796 30126 34848 30132
rect 34244 29844 34296 29850
rect 34244 29786 34296 29792
rect 34256 29714 34284 29786
rect 34244 29708 34296 29714
rect 34244 29650 34296 29656
rect 33600 29640 33652 29646
rect 33600 29582 33652 29588
rect 33692 29640 33744 29646
rect 33692 29582 33744 29588
rect 33704 29510 33732 29582
rect 34612 29572 34664 29578
rect 34612 29514 34664 29520
rect 33416 29504 33468 29510
rect 33416 29446 33468 29452
rect 33692 29504 33744 29510
rect 33692 29446 33744 29452
rect 33428 29102 33456 29446
rect 33968 29232 34020 29238
rect 33968 29174 34020 29180
rect 33416 29096 33468 29102
rect 33416 29038 33468 29044
rect 33428 28558 33456 29038
rect 33416 28552 33468 28558
rect 33416 28494 33468 28500
rect 33508 28076 33560 28082
rect 33508 28018 33560 28024
rect 33520 27606 33548 28018
rect 33508 27600 33560 27606
rect 33508 27542 33560 27548
rect 33600 27600 33652 27606
rect 33600 27542 33652 27548
rect 33612 26450 33640 27542
rect 33980 27334 34008 29174
rect 34520 29096 34572 29102
rect 34520 29038 34572 29044
rect 34336 29028 34388 29034
rect 34336 28970 34388 28976
rect 34348 28642 34376 28970
rect 34532 28762 34560 29038
rect 34520 28756 34572 28762
rect 34520 28698 34572 28704
rect 34624 28694 34652 29514
rect 34808 29306 34836 30126
rect 35268 30002 35296 30194
rect 35268 29974 35388 30002
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35360 29782 35388 29974
rect 35348 29776 35400 29782
rect 35348 29718 35400 29724
rect 34796 29300 34848 29306
rect 34796 29242 34848 29248
rect 34796 28960 34848 28966
rect 34796 28902 34848 28908
rect 34612 28688 34664 28694
rect 34348 28614 34560 28642
rect 34612 28630 34664 28636
rect 34060 28552 34112 28558
rect 34060 28494 34112 28500
rect 34072 28082 34100 28494
rect 34532 28150 34560 28614
rect 34624 28218 34652 28630
rect 34808 28626 34836 28902
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34796 28620 34848 28626
rect 34796 28562 34848 28568
rect 34612 28212 34664 28218
rect 34612 28154 34664 28160
rect 34520 28144 34572 28150
rect 34520 28086 34572 28092
rect 34060 28076 34112 28082
rect 34060 28018 34112 28024
rect 34072 27470 34100 28018
rect 34808 27538 34836 28562
rect 35360 28558 35388 29718
rect 35452 28694 35480 31214
rect 35440 28688 35492 28694
rect 35440 28630 35492 28636
rect 35348 28552 35400 28558
rect 35348 28494 35400 28500
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34796 27532 34848 27538
rect 34796 27474 34848 27480
rect 34060 27464 34112 27470
rect 34060 27406 34112 27412
rect 33968 27328 34020 27334
rect 33968 27270 34020 27276
rect 33600 26444 33652 26450
rect 33600 26386 33652 26392
rect 33232 26376 33284 26382
rect 33232 26318 33284 26324
rect 32772 26036 32824 26042
rect 32772 25978 32824 25984
rect 32416 22066 32628 22094
rect 32600 3194 32628 22066
rect 32588 3188 32640 3194
rect 32588 3130 32640 3136
rect 32600 2446 32628 3130
rect 32588 2440 32640 2446
rect 32588 2382 32640 2388
rect 32220 2304 32272 2310
rect 32220 2246 32272 2252
rect 32036 2100 32088 2106
rect 32036 2042 32088 2048
rect 32232 800 32260 2246
rect 33980 1970 34008 27270
rect 34072 27062 34100 27406
rect 34060 27056 34112 27062
rect 34060 26998 34112 27004
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35636 13870 35664 33390
rect 35716 32904 35768 32910
rect 35716 32846 35768 32852
rect 35728 32434 35756 32846
rect 35716 32428 35768 32434
rect 35716 32370 35768 32376
rect 35728 31890 35756 32370
rect 35820 32298 35848 33934
rect 35912 33930 35940 34614
rect 36452 34604 36504 34610
rect 36452 34546 36504 34552
rect 36268 34536 36320 34542
rect 36268 34478 36320 34484
rect 36280 34202 36308 34478
rect 36268 34196 36320 34202
rect 36268 34138 36320 34144
rect 36464 33998 36492 34546
rect 36176 33992 36228 33998
rect 36176 33934 36228 33940
rect 36452 33992 36504 33998
rect 36452 33934 36504 33940
rect 35900 33924 35952 33930
rect 35900 33866 35952 33872
rect 35912 32570 35940 33866
rect 36084 33856 36136 33862
rect 36084 33798 36136 33804
rect 36096 33114 36124 33798
rect 36188 33658 36216 33934
rect 36176 33652 36228 33658
rect 36176 33594 36228 33600
rect 36268 33652 36320 33658
rect 36268 33594 36320 33600
rect 36176 33516 36228 33522
rect 36280 33504 36308 33594
rect 36464 33590 36492 33934
rect 36452 33584 36504 33590
rect 36452 33526 36504 33532
rect 36228 33476 36308 33504
rect 36176 33458 36228 33464
rect 36188 33386 36216 33458
rect 36176 33380 36228 33386
rect 36176 33322 36228 33328
rect 36084 33108 36136 33114
rect 36084 33050 36136 33056
rect 35900 32564 35952 32570
rect 35900 32506 35952 32512
rect 35900 32360 35952 32366
rect 35900 32302 35952 32308
rect 35808 32292 35860 32298
rect 35808 32234 35860 32240
rect 35912 31958 35940 32302
rect 36544 32224 36596 32230
rect 36544 32166 36596 32172
rect 35900 31952 35952 31958
rect 35900 31894 35952 31900
rect 35716 31884 35768 31890
rect 35716 31826 35768 31832
rect 35728 30394 35756 31826
rect 35912 31822 35940 31894
rect 36556 31890 36584 32166
rect 36544 31884 36596 31890
rect 36544 31826 36596 31832
rect 36740 31822 36768 34614
rect 37002 34575 37058 34584
rect 35900 31816 35952 31822
rect 35900 31758 35952 31764
rect 36728 31816 36780 31822
rect 36728 31758 36780 31764
rect 36082 31648 36138 31657
rect 36082 31583 36138 31592
rect 36096 31142 36124 31583
rect 36084 31136 36136 31142
rect 36084 31078 36136 31084
rect 36452 31136 36504 31142
rect 36452 31078 36504 31084
rect 35900 30592 35952 30598
rect 35900 30534 35952 30540
rect 35992 30592 36044 30598
rect 35992 30534 36044 30540
rect 35716 30388 35768 30394
rect 35716 30330 35768 30336
rect 35912 29714 35940 30534
rect 36004 29850 36032 30534
rect 35992 29844 36044 29850
rect 35992 29786 36044 29792
rect 35900 29708 35952 29714
rect 35900 29650 35952 29656
rect 35808 29640 35860 29646
rect 35808 29582 35860 29588
rect 35820 29306 35848 29582
rect 35808 29300 35860 29306
rect 35808 29242 35860 29248
rect 35624 13864 35676 13870
rect 35624 13806 35676 13812
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 36096 2922 36124 31078
rect 36464 30734 36492 31078
rect 36452 30728 36504 30734
rect 36452 30670 36504 30676
rect 36544 30252 36596 30258
rect 36544 30194 36596 30200
rect 36556 29510 36584 30194
rect 36544 29504 36596 29510
rect 36544 29446 36596 29452
rect 36556 29170 36584 29446
rect 36544 29164 36596 29170
rect 36544 29106 36596 29112
rect 36544 27464 36596 27470
rect 36544 27406 36596 27412
rect 36360 26784 36412 26790
rect 36360 26726 36412 26732
rect 36084 2916 36136 2922
rect 36084 2858 36136 2864
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 36372 2650 36400 26726
rect 36556 26518 36584 27406
rect 36544 26512 36596 26518
rect 36544 26454 36596 26460
rect 37016 22030 37044 34575
rect 37108 30938 37136 37130
rect 37292 36922 37320 37266
rect 37476 37262 37504 37810
rect 37568 37806 37596 38927
rect 37556 37800 37608 37806
rect 37556 37742 37608 37748
rect 37464 37256 37516 37262
rect 37464 37198 37516 37204
rect 37568 37194 37596 37742
rect 37556 37188 37608 37194
rect 37556 37130 37608 37136
rect 37280 36916 37332 36922
rect 37280 36858 37332 36864
rect 37278 36680 37334 36689
rect 37278 36615 37280 36624
rect 37332 36615 37334 36624
rect 37280 36586 37332 36592
rect 37464 36168 37516 36174
rect 37464 36110 37516 36116
rect 37476 35698 37504 36110
rect 37464 35692 37516 35698
rect 37464 35634 37516 35640
rect 37372 35080 37424 35086
rect 37372 35022 37424 35028
rect 37384 33998 37412 35022
rect 37556 34604 37608 34610
rect 37556 34546 37608 34552
rect 37568 34134 37596 34546
rect 37556 34128 37608 34134
rect 37556 34070 37608 34076
rect 37372 33992 37424 33998
rect 37372 33934 37424 33940
rect 37384 33114 37412 33934
rect 37568 33658 37596 34070
rect 37556 33652 37608 33658
rect 37556 33594 37608 33600
rect 37660 33538 37688 39034
rect 37752 36174 37780 40582
rect 37936 40526 37964 41958
rect 38304 41818 38332 42162
rect 38292 41812 38344 41818
rect 38292 41754 38344 41760
rect 38396 41698 38424 43250
rect 38580 42566 38608 43250
rect 39948 43172 40000 43178
rect 39948 43114 40000 43120
rect 39120 43104 39172 43110
rect 39120 43046 39172 43052
rect 38568 42560 38620 42566
rect 38568 42502 38620 42508
rect 38476 42220 38528 42226
rect 38476 42162 38528 42168
rect 38568 42220 38620 42226
rect 38568 42162 38620 42168
rect 38304 41670 38424 41698
rect 38304 41478 38332 41670
rect 38016 41472 38068 41478
rect 38016 41414 38068 41420
rect 38292 41472 38344 41478
rect 38292 41414 38344 41420
rect 38028 41386 38332 41414
rect 37924 40520 37976 40526
rect 37924 40462 37976 40468
rect 37936 39982 37964 40462
rect 37924 39976 37976 39982
rect 37924 39918 37976 39924
rect 38016 39976 38068 39982
rect 38016 39918 38068 39924
rect 38028 38826 38056 39918
rect 38108 39432 38160 39438
rect 38108 39374 38160 39380
rect 38120 38894 38148 39374
rect 38108 38888 38160 38894
rect 38108 38830 38160 38836
rect 38016 38820 38068 38826
rect 38016 38762 38068 38768
rect 38200 38752 38252 38758
rect 38200 38694 38252 38700
rect 37922 38584 37978 38593
rect 37922 38519 37978 38528
rect 37832 38276 37884 38282
rect 37832 38218 37884 38224
rect 37844 37670 37872 38218
rect 37832 37664 37884 37670
rect 37832 37606 37884 37612
rect 37936 37466 37964 38519
rect 38212 38350 38240 38694
rect 38108 38344 38160 38350
rect 38106 38312 38108 38321
rect 38200 38344 38252 38350
rect 38160 38312 38162 38321
rect 38200 38286 38252 38292
rect 38106 38247 38162 38256
rect 38304 38026 38332 41386
rect 38488 41206 38516 42162
rect 38580 41750 38608 42162
rect 39132 42158 39160 43046
rect 39960 42906 39988 43114
rect 40224 43104 40276 43110
rect 40224 43046 40276 43052
rect 39948 42900 40000 42906
rect 39948 42842 40000 42848
rect 40040 42560 40092 42566
rect 40040 42502 40092 42508
rect 39120 42152 39172 42158
rect 39120 42094 39172 42100
rect 40052 42022 40080 42502
rect 40236 42022 40264 43046
rect 39304 42016 39356 42022
rect 39304 41958 39356 41964
rect 40040 42016 40092 42022
rect 40040 41958 40092 41964
rect 40224 42016 40276 42022
rect 40224 41958 40276 41964
rect 38568 41744 38620 41750
rect 38568 41686 38620 41692
rect 38476 41200 38528 41206
rect 38476 41142 38528 41148
rect 38384 39500 38436 39506
rect 38384 39442 38436 39448
rect 38028 37998 38332 38026
rect 38396 38010 38424 39442
rect 38384 38004 38436 38010
rect 37924 37460 37976 37466
rect 37924 37402 37976 37408
rect 37740 36168 37792 36174
rect 37740 36110 37792 36116
rect 37924 35080 37976 35086
rect 37924 35022 37976 35028
rect 37832 33856 37884 33862
rect 37832 33798 37884 33804
rect 37568 33510 37688 33538
rect 37738 33552 37794 33561
rect 37372 33108 37424 33114
rect 37372 33050 37424 33056
rect 37464 32428 37516 32434
rect 37464 32370 37516 32376
rect 37476 31822 37504 32370
rect 37464 31816 37516 31822
rect 37464 31758 37516 31764
rect 37280 31136 37332 31142
rect 37280 31078 37332 31084
rect 37096 30932 37148 30938
rect 37096 30874 37148 30880
rect 37108 30666 37136 30874
rect 37096 30660 37148 30666
rect 37096 30602 37148 30608
rect 37108 30394 37136 30602
rect 37096 30388 37148 30394
rect 37096 30330 37148 30336
rect 37292 30258 37320 31078
rect 37280 30252 37332 30258
rect 37280 30194 37332 30200
rect 37292 29102 37320 30194
rect 37476 29850 37504 31758
rect 37464 29844 37516 29850
rect 37464 29786 37516 29792
rect 37280 29096 37332 29102
rect 37280 29038 37332 29044
rect 37568 28218 37596 33510
rect 37738 33487 37740 33496
rect 37792 33487 37794 33496
rect 37740 33458 37792 33464
rect 37648 32904 37700 32910
rect 37648 32846 37700 32852
rect 37660 32570 37688 32846
rect 37740 32836 37792 32842
rect 37740 32778 37792 32784
rect 37648 32564 37700 32570
rect 37648 32506 37700 32512
rect 37752 32434 37780 32778
rect 37740 32428 37792 32434
rect 37740 32370 37792 32376
rect 37648 31748 37700 31754
rect 37648 31690 37700 31696
rect 37660 31482 37688 31690
rect 37648 31476 37700 31482
rect 37648 31418 37700 31424
rect 37648 31340 37700 31346
rect 37752 31328 37780 32370
rect 37844 31890 37872 33798
rect 37936 33114 37964 35022
rect 38028 33454 38056 37998
rect 38384 37946 38436 37952
rect 38108 37936 38160 37942
rect 38488 37890 38516 41142
rect 38580 41138 38608 41686
rect 39316 41614 39344 41958
rect 40052 41818 40080 41958
rect 40040 41812 40092 41818
rect 40040 41754 40092 41760
rect 38752 41608 38804 41614
rect 38752 41550 38804 41556
rect 39304 41608 39356 41614
rect 39304 41550 39356 41556
rect 38764 41274 38792 41550
rect 38752 41268 38804 41274
rect 38752 41210 38804 41216
rect 38568 41132 38620 41138
rect 38568 41074 38620 41080
rect 40052 41002 40080 41754
rect 40236 41750 40264 41958
rect 40224 41744 40276 41750
rect 40224 41686 40276 41692
rect 40236 41274 40264 41686
rect 40500 41472 40552 41478
rect 40500 41414 40552 41420
rect 40224 41268 40276 41274
rect 40224 41210 40276 41216
rect 40040 40996 40092 41002
rect 40040 40938 40092 40944
rect 39672 40928 39724 40934
rect 39672 40870 39724 40876
rect 39684 40390 39712 40870
rect 38660 40384 38712 40390
rect 38660 40326 38712 40332
rect 39672 40384 39724 40390
rect 39672 40326 39724 40332
rect 38672 39642 38700 40326
rect 38844 40044 38896 40050
rect 38844 39986 38896 39992
rect 39488 40044 39540 40050
rect 39488 39986 39540 39992
rect 38856 39642 38884 39986
rect 39120 39908 39172 39914
rect 39120 39850 39172 39856
rect 39132 39642 39160 39850
rect 38660 39636 38712 39642
rect 38660 39578 38712 39584
rect 38844 39636 38896 39642
rect 38844 39578 38896 39584
rect 39028 39636 39080 39642
rect 39028 39578 39080 39584
rect 39120 39636 39172 39642
rect 39120 39578 39172 39584
rect 38672 39522 38700 39578
rect 39040 39522 39068 39578
rect 38672 39494 39068 39522
rect 38660 39364 38712 39370
rect 38660 39306 38712 39312
rect 38672 39030 38700 39306
rect 38752 39296 38804 39302
rect 38752 39238 38804 39244
rect 38568 39024 38620 39030
rect 38566 38992 38568 39001
rect 38660 39024 38712 39030
rect 38620 38992 38622 39001
rect 38660 38966 38712 38972
rect 38566 38927 38622 38936
rect 38580 38418 38608 38927
rect 38568 38412 38620 38418
rect 38568 38354 38620 38360
rect 38764 38350 38792 39238
rect 38752 38344 38804 38350
rect 38752 38286 38804 38292
rect 38108 37878 38160 37884
rect 38120 37398 38148 37878
rect 38304 37862 38516 37890
rect 38108 37392 38160 37398
rect 38108 37334 38160 37340
rect 38120 36922 38148 37334
rect 38108 36916 38160 36922
rect 38108 36858 38160 36864
rect 38120 35222 38148 36858
rect 38200 36576 38252 36582
rect 38200 36518 38252 36524
rect 38212 36174 38240 36518
rect 38200 36168 38252 36174
rect 38200 36110 38252 36116
rect 38212 35834 38240 36110
rect 38304 35850 38332 37862
rect 38476 37800 38528 37806
rect 38476 37742 38528 37748
rect 38488 36854 38516 37742
rect 38568 37256 38620 37262
rect 38568 37198 38620 37204
rect 38476 36848 38528 36854
rect 38476 36790 38528 36796
rect 38580 36786 38608 37198
rect 38384 36780 38436 36786
rect 38384 36722 38436 36728
rect 38568 36780 38620 36786
rect 38568 36722 38620 36728
rect 38396 36378 38424 36722
rect 38660 36644 38712 36650
rect 38660 36586 38712 36592
rect 38384 36372 38436 36378
rect 38384 36314 38436 36320
rect 38672 36310 38700 36586
rect 38660 36304 38712 36310
rect 38660 36246 38712 36252
rect 38200 35828 38252 35834
rect 38304 35822 38424 35850
rect 38856 35834 38884 39494
rect 39118 39400 39174 39409
rect 39118 39335 39120 39344
rect 39172 39335 39174 39344
rect 39120 39306 39172 39312
rect 38936 39092 38988 39098
rect 38936 39034 38988 39040
rect 38948 38350 38976 39034
rect 39500 39030 39528 39986
rect 40052 39914 40080 40938
rect 40236 40730 40264 41210
rect 40224 40724 40276 40730
rect 40224 40666 40276 40672
rect 40512 40050 40540 41414
rect 43168 40928 43220 40934
rect 43168 40870 43220 40876
rect 41052 40656 41104 40662
rect 41052 40598 41104 40604
rect 41064 40390 41092 40598
rect 41604 40452 41656 40458
rect 41604 40394 41656 40400
rect 41052 40384 41104 40390
rect 41052 40326 41104 40332
rect 41512 40384 41564 40390
rect 41512 40326 41564 40332
rect 40500 40044 40552 40050
rect 40500 39986 40552 39992
rect 40224 39976 40276 39982
rect 40224 39918 40276 39924
rect 40040 39908 40092 39914
rect 40040 39850 40092 39856
rect 39856 39840 39908 39846
rect 39856 39782 39908 39788
rect 39868 39438 39896 39782
rect 39856 39432 39908 39438
rect 39762 39400 39818 39409
rect 39856 39374 39908 39380
rect 39762 39335 39818 39344
rect 39488 39024 39540 39030
rect 39488 38966 39540 38972
rect 39028 38956 39080 38962
rect 39028 38898 39080 38904
rect 38936 38344 38988 38350
rect 38936 38286 38988 38292
rect 39040 37670 39068 38898
rect 39672 38752 39724 38758
rect 39672 38694 39724 38700
rect 39684 38214 39712 38694
rect 39672 38208 39724 38214
rect 39672 38150 39724 38156
rect 39120 37868 39172 37874
rect 39120 37810 39172 37816
rect 39028 37664 39080 37670
rect 39028 37606 39080 37612
rect 39132 37262 39160 37810
rect 39210 37768 39266 37777
rect 39210 37703 39212 37712
rect 39264 37703 39266 37712
rect 39212 37674 39264 37680
rect 39120 37256 39172 37262
rect 39120 37198 39172 37204
rect 39488 37256 39540 37262
rect 39488 37198 39540 37204
rect 39132 36582 39160 37198
rect 39500 36786 39528 37198
rect 39488 36780 39540 36786
rect 39488 36722 39540 36728
rect 39120 36576 39172 36582
rect 39120 36518 39172 36524
rect 39212 36168 39264 36174
rect 39212 36110 39264 36116
rect 38200 35770 38252 35776
rect 38292 35760 38344 35766
rect 38292 35702 38344 35708
rect 38108 35216 38160 35222
rect 38108 35158 38160 35164
rect 38200 35080 38252 35086
rect 38200 35022 38252 35028
rect 38108 34944 38160 34950
rect 38108 34886 38160 34892
rect 38120 34610 38148 34886
rect 38108 34604 38160 34610
rect 38108 34546 38160 34552
rect 38120 33998 38148 34546
rect 38212 34066 38240 35022
rect 38304 34746 38332 35702
rect 38292 34740 38344 34746
rect 38292 34682 38344 34688
rect 38200 34060 38252 34066
rect 38200 34002 38252 34008
rect 38108 33992 38160 33998
rect 38108 33934 38160 33940
rect 38396 33590 38424 35822
rect 38844 35828 38896 35834
rect 38844 35770 38896 35776
rect 38856 35698 38884 35770
rect 38844 35692 38896 35698
rect 38844 35634 38896 35640
rect 39028 35692 39080 35698
rect 39028 35634 39080 35640
rect 38856 35222 38884 35634
rect 39040 35494 39068 35634
rect 39224 35562 39252 36110
rect 39302 35864 39358 35873
rect 39302 35799 39358 35808
rect 39212 35556 39264 35562
rect 39212 35498 39264 35504
rect 39028 35488 39080 35494
rect 39028 35430 39080 35436
rect 38568 35216 38620 35222
rect 38568 35158 38620 35164
rect 38844 35216 38896 35222
rect 38844 35158 38896 35164
rect 38384 33584 38436 33590
rect 38384 33526 38436 33532
rect 38108 33516 38160 33522
rect 38108 33458 38160 33464
rect 38016 33448 38068 33454
rect 38016 33390 38068 33396
rect 37924 33108 37976 33114
rect 37924 33050 37976 33056
rect 37832 31884 37884 31890
rect 37832 31826 37884 31832
rect 37844 31346 37872 31826
rect 37700 31300 37780 31328
rect 37832 31340 37884 31346
rect 37648 31282 37700 31288
rect 37832 31282 37884 31288
rect 38028 30938 38056 33390
rect 38120 32910 38148 33458
rect 38396 32910 38424 33526
rect 38108 32904 38160 32910
rect 38108 32846 38160 32852
rect 38384 32904 38436 32910
rect 38384 32846 38436 32852
rect 38120 32434 38148 32846
rect 38108 32428 38160 32434
rect 38108 32370 38160 32376
rect 38396 32366 38424 32846
rect 38384 32360 38436 32366
rect 38384 32302 38436 32308
rect 38396 32026 38424 32302
rect 38580 32298 38608 35158
rect 39040 34746 39068 35430
rect 39120 35012 39172 35018
rect 39120 34954 39172 34960
rect 38660 34740 38712 34746
rect 38660 34682 38712 34688
rect 39028 34740 39080 34746
rect 39028 34682 39080 34688
rect 38672 34066 38700 34682
rect 39132 34610 39160 34954
rect 39316 34950 39344 35799
rect 39304 34944 39356 34950
rect 39304 34886 39356 34892
rect 39120 34604 39172 34610
rect 39120 34546 39172 34552
rect 39304 34604 39356 34610
rect 39304 34546 39356 34552
rect 38660 34060 38712 34066
rect 38660 34002 38712 34008
rect 38672 33658 38700 34002
rect 38660 33652 38712 33658
rect 38660 33594 38712 33600
rect 39132 33522 39160 34546
rect 39316 33522 39344 34546
rect 39120 33516 39172 33522
rect 39120 33458 39172 33464
rect 39304 33516 39356 33522
rect 39304 33458 39356 33464
rect 38660 32768 38712 32774
rect 38660 32710 38712 32716
rect 38672 32502 38700 32710
rect 38660 32496 38712 32502
rect 38660 32438 38712 32444
rect 38568 32292 38620 32298
rect 38568 32234 38620 32240
rect 38384 32020 38436 32026
rect 38384 31962 38436 31968
rect 38476 31884 38528 31890
rect 38580 31872 38608 32234
rect 38672 31890 38700 32438
rect 38752 32428 38804 32434
rect 38752 32370 38804 32376
rect 38528 31844 38608 31872
rect 38476 31826 38528 31832
rect 38580 31754 38608 31844
rect 38660 31884 38712 31890
rect 38660 31826 38712 31832
rect 38580 31726 38700 31754
rect 38580 31414 38608 31726
rect 38568 31408 38620 31414
rect 38568 31350 38620 31356
rect 38672 31142 38700 31726
rect 38764 31142 38792 32370
rect 38844 31816 38896 31822
rect 38844 31758 38896 31764
rect 38856 31482 38884 31758
rect 38844 31476 38896 31482
rect 38844 31418 38896 31424
rect 38660 31136 38712 31142
rect 38660 31078 38712 31084
rect 38752 31136 38804 31142
rect 38752 31078 38804 31084
rect 38016 30932 38068 30938
rect 38016 30874 38068 30880
rect 38672 30394 38700 31078
rect 38764 30938 38792 31078
rect 38752 30932 38804 30938
rect 38752 30874 38804 30880
rect 38660 30388 38712 30394
rect 38660 30330 38712 30336
rect 39396 30388 39448 30394
rect 39396 30330 39448 30336
rect 37556 28212 37608 28218
rect 37556 28154 37608 28160
rect 37004 22024 37056 22030
rect 37004 21966 37056 21972
rect 39408 20058 39436 30330
rect 39500 30190 39528 36722
rect 39684 34202 39712 38150
rect 39776 35086 39804 39335
rect 39856 39296 39908 39302
rect 39856 39238 39908 39244
rect 39868 39098 39896 39238
rect 39856 39092 39908 39098
rect 39856 39034 39908 39040
rect 40236 38962 40264 39918
rect 40960 39840 41012 39846
rect 40960 39782 41012 39788
rect 40972 39574 41000 39782
rect 40960 39568 41012 39574
rect 40960 39510 41012 39516
rect 40592 39296 40644 39302
rect 40592 39238 40644 39244
rect 40224 38956 40276 38962
rect 40224 38898 40276 38904
rect 40604 38350 40632 39238
rect 40868 38956 40920 38962
rect 40868 38898 40920 38904
rect 40592 38344 40644 38350
rect 40592 38286 40644 38292
rect 39856 38208 39908 38214
rect 39856 38150 39908 38156
rect 39868 37913 39896 38150
rect 39854 37904 39910 37913
rect 39854 37839 39910 37848
rect 40132 37868 40184 37874
rect 40132 37810 40184 37816
rect 39948 37256 40000 37262
rect 39948 37198 40000 37204
rect 39960 36718 39988 37198
rect 40144 37194 40172 37810
rect 40604 37466 40632 38286
rect 40592 37460 40644 37466
rect 40592 37402 40644 37408
rect 40776 37256 40828 37262
rect 40880 37244 40908 38898
rect 41064 38010 41092 40326
rect 41328 39908 41380 39914
rect 41328 39850 41380 39856
rect 41052 38004 41104 38010
rect 41052 37946 41104 37952
rect 41144 37800 41196 37806
rect 41144 37742 41196 37748
rect 41156 37466 41184 37742
rect 41144 37460 41196 37466
rect 41144 37402 41196 37408
rect 41236 37392 41288 37398
rect 41236 37334 41288 37340
rect 40828 37216 40908 37244
rect 40776 37198 40828 37204
rect 40132 37188 40184 37194
rect 40132 37130 40184 37136
rect 40040 37120 40092 37126
rect 40040 37062 40092 37068
rect 39948 36712 40000 36718
rect 39948 36654 40000 36660
rect 39856 36576 39908 36582
rect 39856 36518 39908 36524
rect 39868 36174 39896 36518
rect 40052 36310 40080 37062
rect 40040 36304 40092 36310
rect 40040 36246 40092 36252
rect 39856 36168 39908 36174
rect 39856 36110 39908 36116
rect 39856 36032 39908 36038
rect 39856 35974 39908 35980
rect 39764 35080 39816 35086
rect 39764 35022 39816 35028
rect 39764 34944 39816 34950
rect 39764 34886 39816 34892
rect 39672 34196 39724 34202
rect 39672 34138 39724 34144
rect 39580 33516 39632 33522
rect 39580 33458 39632 33464
rect 39592 32366 39620 33458
rect 39672 32768 39724 32774
rect 39672 32710 39724 32716
rect 39684 32502 39712 32710
rect 39672 32496 39724 32502
rect 39672 32438 39724 32444
rect 39580 32360 39632 32366
rect 39580 32302 39632 32308
rect 39488 30184 39540 30190
rect 39488 30126 39540 30132
rect 39592 26994 39620 32302
rect 39580 26988 39632 26994
rect 39580 26930 39632 26936
rect 39684 26874 39712 32438
rect 39500 26846 39712 26874
rect 39396 20052 39448 20058
rect 39396 19994 39448 20000
rect 39500 4146 39528 26846
rect 39580 26784 39632 26790
rect 39580 26726 39632 26732
rect 39592 15910 39620 26726
rect 39776 24410 39804 34886
rect 39868 34406 39896 35974
rect 40052 35698 40080 36246
rect 40144 36174 40172 37130
rect 40224 37120 40276 37126
rect 40224 37062 40276 37068
rect 40236 36922 40264 37062
rect 40224 36916 40276 36922
rect 40224 36858 40276 36864
rect 40880 36854 40908 37216
rect 40408 36848 40460 36854
rect 40408 36790 40460 36796
rect 40868 36848 40920 36854
rect 40868 36790 40920 36796
rect 40316 36644 40368 36650
rect 40316 36586 40368 36592
rect 40132 36168 40184 36174
rect 40132 36110 40184 36116
rect 40040 35692 40092 35698
rect 40040 35634 40092 35640
rect 40144 35494 40172 36110
rect 40328 36038 40356 36586
rect 40420 36378 40448 36790
rect 40408 36372 40460 36378
rect 40408 36314 40460 36320
rect 40880 36174 40908 36790
rect 41248 36786 41276 37334
rect 41236 36780 41288 36786
rect 41236 36722 41288 36728
rect 40868 36168 40920 36174
rect 41248 36152 41276 36722
rect 40868 36110 40920 36116
rect 41236 36146 41288 36152
rect 41236 36088 41288 36094
rect 40316 36032 40368 36038
rect 40316 35974 40368 35980
rect 40328 35698 40356 35974
rect 40316 35692 40368 35698
rect 40316 35634 40368 35640
rect 40132 35488 40184 35494
rect 40132 35430 40184 35436
rect 40132 35148 40184 35154
rect 40132 35090 40184 35096
rect 39946 35048 40002 35057
rect 39946 34983 39948 34992
rect 40000 34983 40002 34992
rect 39948 34954 40000 34960
rect 39960 34746 39988 34954
rect 39948 34740 40000 34746
rect 39948 34682 40000 34688
rect 39856 34400 39908 34406
rect 39856 34342 39908 34348
rect 39946 34096 40002 34105
rect 39946 34031 40002 34040
rect 39856 33380 39908 33386
rect 39856 33322 39908 33328
rect 39868 33046 39896 33322
rect 39856 33040 39908 33046
rect 39856 32982 39908 32988
rect 39868 32570 39896 32982
rect 39960 32910 39988 34031
rect 40144 33522 40172 35090
rect 40868 35080 40920 35086
rect 40868 35022 40920 35028
rect 40408 34604 40460 34610
rect 40408 34546 40460 34552
rect 40592 34604 40644 34610
rect 40592 34546 40644 34552
rect 40316 34128 40368 34134
rect 40316 34070 40368 34076
rect 40132 33516 40184 33522
rect 40132 33458 40184 33464
rect 40040 33448 40092 33454
rect 40040 33390 40092 33396
rect 40052 33114 40080 33390
rect 40040 33108 40092 33114
rect 40040 33050 40092 33056
rect 40328 32910 40356 34070
rect 40420 33590 40448 34546
rect 40604 34066 40632 34546
rect 40788 34134 40816 34165
rect 40776 34128 40828 34134
rect 40774 34096 40776 34105
rect 40828 34096 40830 34105
rect 40592 34060 40644 34066
rect 40774 34031 40830 34040
rect 40592 34002 40644 34008
rect 40788 33998 40816 34031
rect 40776 33992 40828 33998
rect 40776 33934 40828 33940
rect 40684 33856 40736 33862
rect 40684 33798 40736 33804
rect 40408 33584 40460 33590
rect 40408 33526 40460 33532
rect 40696 33522 40724 33798
rect 40684 33516 40736 33522
rect 40684 33458 40736 33464
rect 40408 33312 40460 33318
rect 40408 33254 40460 33260
rect 40420 32910 40448 33254
rect 40696 32978 40724 33458
rect 40788 33318 40816 33934
rect 40880 33522 40908 35022
rect 41248 34746 41276 36088
rect 41236 34740 41288 34746
rect 41236 34682 41288 34688
rect 41052 33652 41104 33658
rect 41052 33594 41104 33600
rect 41064 33522 41092 33594
rect 40868 33516 40920 33522
rect 41052 33516 41104 33522
rect 40920 33476 41000 33504
rect 40868 33458 40920 33464
rect 40776 33312 40828 33318
rect 40776 33254 40828 33260
rect 40868 33312 40920 33318
rect 40868 33254 40920 33260
rect 40880 33114 40908 33254
rect 40868 33108 40920 33114
rect 40868 33050 40920 33056
rect 40684 32972 40736 32978
rect 40684 32914 40736 32920
rect 39948 32904 40000 32910
rect 39948 32846 40000 32852
rect 40316 32904 40368 32910
rect 40316 32846 40368 32852
rect 40408 32904 40460 32910
rect 40408 32846 40460 32852
rect 39856 32564 39908 32570
rect 39856 32506 39908 32512
rect 39960 31482 39988 32846
rect 40408 32224 40460 32230
rect 40408 32166 40460 32172
rect 40420 32026 40448 32166
rect 40696 32026 40724 32914
rect 40972 32366 41000 33476
rect 41052 33458 41104 33464
rect 40960 32360 41012 32366
rect 40960 32302 41012 32308
rect 40408 32020 40460 32026
rect 40408 31962 40460 31968
rect 40684 32020 40736 32026
rect 40684 31962 40736 31968
rect 39948 31476 40000 31482
rect 39948 31418 40000 31424
rect 39764 24404 39816 24410
rect 39764 24346 39816 24352
rect 41340 22094 41368 39850
rect 41524 39438 41552 40326
rect 41616 40186 41644 40394
rect 42064 40384 42116 40390
rect 42064 40326 42116 40332
rect 41604 40180 41656 40186
rect 41604 40122 41656 40128
rect 41696 40044 41748 40050
rect 41696 39986 41748 39992
rect 41512 39432 41564 39438
rect 41512 39374 41564 39380
rect 41602 39400 41658 39409
rect 41602 39335 41604 39344
rect 41656 39335 41658 39344
rect 41604 39306 41656 39312
rect 41708 38010 41736 39986
rect 42076 39846 42104 40326
rect 43180 39846 43208 40870
rect 42064 39840 42116 39846
rect 42064 39782 42116 39788
rect 43168 39840 43220 39846
rect 43168 39782 43220 39788
rect 42076 39370 42104 39782
rect 42064 39364 42116 39370
rect 42064 39306 42116 39312
rect 42708 39296 42760 39302
rect 42708 39238 42760 39244
rect 42720 38894 42748 39238
rect 43180 39030 43208 39782
rect 43536 39500 43588 39506
rect 43536 39442 43588 39448
rect 43548 39098 43576 39442
rect 43536 39092 43588 39098
rect 43536 39034 43588 39040
rect 43168 39024 43220 39030
rect 43168 38966 43220 38972
rect 42708 38888 42760 38894
rect 42628 38836 42708 38842
rect 42628 38830 42760 38836
rect 42628 38814 42748 38830
rect 42628 38554 42656 38814
rect 42708 38752 42760 38758
rect 42708 38694 42760 38700
rect 42984 38752 43036 38758
rect 42984 38694 43036 38700
rect 42616 38548 42668 38554
rect 42616 38490 42668 38496
rect 42156 38276 42208 38282
rect 42156 38218 42208 38224
rect 41696 38004 41748 38010
rect 41696 37946 41748 37952
rect 41420 35488 41472 35494
rect 41420 35430 41472 35436
rect 41512 35488 41564 35494
rect 41512 35430 41564 35436
rect 41432 35086 41460 35430
rect 41524 35290 41552 35430
rect 41512 35284 41564 35290
rect 41512 35226 41564 35232
rect 41420 35080 41472 35086
rect 41420 35022 41472 35028
rect 41512 35012 41564 35018
rect 41512 34954 41564 34960
rect 41420 33380 41472 33386
rect 41420 33322 41472 33328
rect 41432 33046 41460 33322
rect 41420 33040 41472 33046
rect 41420 32982 41472 32988
rect 41524 32774 41552 34954
rect 41708 34950 41736 37946
rect 42168 37398 42196 38218
rect 42156 37392 42208 37398
rect 42156 37334 42208 37340
rect 41880 36372 41932 36378
rect 41880 36314 41932 36320
rect 41892 35018 41920 36314
rect 42168 35494 42196 37334
rect 42628 36922 42656 38490
rect 42720 38350 42748 38694
rect 42996 38486 43024 38694
rect 42984 38480 43036 38486
rect 42984 38422 43036 38428
rect 42708 38344 42760 38350
rect 42708 38286 42760 38292
rect 42996 38010 43024 38422
rect 43180 38214 43208 38966
rect 43352 38344 43404 38350
rect 43352 38286 43404 38292
rect 43168 38208 43220 38214
rect 43168 38150 43220 38156
rect 42984 38004 43036 38010
rect 42984 37946 43036 37952
rect 42616 36916 42668 36922
rect 42616 36858 42668 36864
rect 42628 36378 42656 36858
rect 42616 36372 42668 36378
rect 42616 36314 42668 36320
rect 42984 36032 43036 36038
rect 42984 35974 43036 35980
rect 42996 35494 43024 35974
rect 42156 35488 42208 35494
rect 42156 35430 42208 35436
rect 42984 35488 43036 35494
rect 42984 35430 43036 35436
rect 41972 35080 42024 35086
rect 41972 35022 42024 35028
rect 41880 35012 41932 35018
rect 41880 34954 41932 34960
rect 41696 34944 41748 34950
rect 41696 34886 41748 34892
rect 41984 34082 42012 35022
rect 43076 34944 43128 34950
rect 43076 34886 43128 34892
rect 42064 34536 42116 34542
rect 42064 34478 42116 34484
rect 42076 34202 42104 34478
rect 42064 34196 42116 34202
rect 42064 34138 42116 34144
rect 42524 34128 42576 34134
rect 41984 34054 42104 34082
rect 42524 34070 42576 34076
rect 41512 32768 41564 32774
rect 41512 32710 41564 32716
rect 41972 32768 42024 32774
rect 41972 32710 42024 32716
rect 41984 32230 42012 32710
rect 41972 32224 42024 32230
rect 41972 32166 42024 32172
rect 41248 22066 41368 22094
rect 41248 18290 41276 22066
rect 41236 18284 41288 18290
rect 41236 18226 41288 18232
rect 42076 16250 42104 34054
rect 42536 33046 42564 34070
rect 43088 33590 43116 34886
rect 43180 33862 43208 38150
rect 43364 37466 43392 38286
rect 43352 37460 43404 37466
rect 43352 37402 43404 37408
rect 43364 36922 43392 37402
rect 43352 36916 43404 36922
rect 43352 36858 43404 36864
rect 44180 36848 44232 36854
rect 44178 36816 44180 36825
rect 44232 36816 44234 36825
rect 44178 36751 44234 36760
rect 45480 35737 45508 46922
rect 46216 46374 46244 46990
rect 47124 46980 47176 46986
rect 47124 46922 47176 46928
rect 46756 46436 46808 46442
rect 46756 46378 46808 46384
rect 46204 46368 46256 46374
rect 46204 46310 46256 46316
rect 46216 45830 46244 46310
rect 46204 45824 46256 45830
rect 46204 45766 46256 45772
rect 45466 35728 45522 35737
rect 45466 35663 45522 35672
rect 43260 35488 43312 35494
rect 43260 35430 43312 35436
rect 43536 35488 43588 35494
rect 43536 35430 43588 35436
rect 43168 33856 43220 33862
rect 43168 33798 43220 33804
rect 43076 33584 43128 33590
rect 43076 33526 43128 33532
rect 43180 33318 43208 33798
rect 43168 33312 43220 33318
rect 43168 33254 43220 33260
rect 42524 33040 42576 33046
rect 42524 32982 42576 32988
rect 43272 32434 43300 35430
rect 43548 35290 43576 35430
rect 43536 35284 43588 35290
rect 43536 35226 43588 35232
rect 44180 33312 44232 33318
rect 44180 33254 44232 33260
rect 43260 32428 43312 32434
rect 43260 32370 43312 32376
rect 42064 16244 42116 16250
rect 42064 16186 42116 16192
rect 39580 15904 39632 15910
rect 39580 15846 39632 15852
rect 39488 4140 39540 4146
rect 39488 4082 39540 4088
rect 40040 2848 40092 2854
rect 40040 2790 40092 2796
rect 36360 2644 36412 2650
rect 36360 2586 36412 2592
rect 40052 2446 40080 2790
rect 44192 2582 44220 33254
rect 46768 31249 46796 46378
rect 47032 45892 47084 45898
rect 47032 45834 47084 45840
rect 47044 44441 47072 45834
rect 47030 44432 47086 44441
rect 47030 44367 47086 44376
rect 47136 39506 47164 46922
rect 47216 46640 47268 46646
rect 47216 46582 47268 46588
rect 47228 46102 47256 46582
rect 47216 46096 47268 46102
rect 47216 46038 47268 46044
rect 48056 45966 48084 48311
rect 48332 47054 48360 49200
rect 48320 47048 48372 47054
rect 48320 46990 48372 46996
rect 48136 46572 48188 46578
rect 48136 46514 48188 46520
rect 48148 46345 48176 46514
rect 48134 46336 48190 46345
rect 48134 46271 48190 46280
rect 48148 46170 48176 46271
rect 48136 46164 48188 46170
rect 48136 46106 48188 46112
rect 48044 45960 48096 45966
rect 48044 45902 48096 45908
rect 48056 45626 48084 45902
rect 48044 45620 48096 45626
rect 48044 45562 48096 45568
rect 48332 45554 48360 46990
rect 49620 46646 49648 49200
rect 49608 46640 49660 46646
rect 49608 46582 49660 46588
rect 48148 45526 48360 45554
rect 48148 45082 48176 45526
rect 47952 45076 48004 45082
rect 47952 45018 48004 45024
rect 48136 45076 48188 45082
rect 48136 45018 48188 45024
rect 47964 44538 47992 45018
rect 47952 44532 48004 44538
rect 47952 44474 48004 44480
rect 48044 44396 48096 44402
rect 48044 44338 48096 44344
rect 48056 44305 48084 44338
rect 48042 44296 48098 44305
rect 48042 44231 48098 44240
rect 48056 43994 48084 44231
rect 48044 43988 48096 43994
rect 48044 43930 48096 43936
rect 48136 42696 48188 42702
rect 48136 42638 48188 42644
rect 47952 42560 48004 42566
rect 47952 42502 48004 42508
rect 47306 40488 47362 40497
rect 47306 40423 47308 40432
rect 47360 40423 47362 40432
rect 47308 40394 47360 40400
rect 47124 39500 47176 39506
rect 47124 39442 47176 39448
rect 47768 37120 47820 37126
rect 47582 37088 47638 37097
rect 47768 37062 47820 37068
rect 47582 37023 47638 37032
rect 47596 36854 47624 37023
rect 47584 36848 47636 36854
rect 47584 36790 47636 36796
rect 47780 36786 47808 37062
rect 47964 36786 47992 42502
rect 48148 42265 48176 42638
rect 48134 42256 48190 42265
rect 48134 42191 48190 42200
rect 48044 40384 48096 40390
rect 48044 40326 48096 40332
rect 48056 40225 48084 40326
rect 48042 40216 48098 40225
rect 48042 40151 48098 40160
rect 48044 38208 48096 38214
rect 48042 38176 48044 38185
rect 48096 38176 48098 38185
rect 48042 38111 48098 38120
rect 47768 36780 47820 36786
rect 47768 36722 47820 36728
rect 47952 36780 48004 36786
rect 47952 36722 48004 36728
rect 47780 36650 47808 36722
rect 47216 36644 47268 36650
rect 47216 36586 47268 36592
rect 47768 36644 47820 36650
rect 47768 36586 47820 36592
rect 47228 36378 47256 36586
rect 47216 36372 47268 36378
rect 47216 36314 47268 36320
rect 47780 35894 47808 36586
rect 47858 36136 47914 36145
rect 47858 36071 47860 36080
rect 47912 36071 47914 36080
rect 48042 36136 48098 36145
rect 48042 36071 48044 36080
rect 47860 36042 47912 36048
rect 48096 36071 48098 36080
rect 48044 36042 48096 36048
rect 47780 35866 47992 35894
rect 47860 33992 47912 33998
rect 47860 33934 47912 33940
rect 47872 33522 47900 33934
rect 47860 33516 47912 33522
rect 47860 33458 47912 33464
rect 47860 32768 47912 32774
rect 47860 32710 47912 32716
rect 47676 32428 47728 32434
rect 47676 32370 47728 32376
rect 47688 32026 47716 32370
rect 47676 32020 47728 32026
rect 47676 31962 47728 31968
rect 46754 31240 46810 31249
rect 46754 31175 46810 31184
rect 46388 29640 46440 29646
rect 46388 29582 46440 29588
rect 45284 28416 45336 28422
rect 45284 28358 45336 28364
rect 45296 2650 45324 28358
rect 46400 27606 46428 29582
rect 46388 27600 46440 27606
rect 46388 27542 46440 27548
rect 47676 18284 47728 18290
rect 47676 18226 47728 18232
rect 47688 17882 47716 18226
rect 47676 17876 47728 17882
rect 47676 17818 47728 17824
rect 47872 16574 47900 32710
rect 47780 16546 47900 16574
rect 47780 11898 47808 16546
rect 47858 13968 47914 13977
rect 47858 13903 47860 13912
rect 47912 13903 47914 13912
rect 47860 13874 47912 13880
rect 47872 13530 47900 13874
rect 47860 13524 47912 13530
rect 47860 13466 47912 13472
rect 47768 11892 47820 11898
rect 47768 11834 47820 11840
rect 47964 8090 47992 35866
rect 48056 35834 48084 36042
rect 48044 35828 48096 35834
rect 48044 35770 48096 35776
rect 48134 34096 48190 34105
rect 48134 34031 48136 34040
rect 48188 34031 48190 34040
rect 48136 34002 48188 34008
rect 48148 33658 48176 34002
rect 48136 33652 48188 33658
rect 48136 33594 48188 33600
rect 48044 32224 48096 32230
rect 48044 32166 48096 32172
rect 48056 32065 48084 32166
rect 48042 32056 48098 32065
rect 48042 31991 48098 32000
rect 48134 30016 48190 30025
rect 48134 29951 48190 29960
rect 48148 29714 48176 29951
rect 48136 29708 48188 29714
rect 48136 29650 48188 29656
rect 48148 29306 48176 29650
rect 48136 29300 48188 29306
rect 48136 29242 48188 29248
rect 48134 27976 48190 27985
rect 48134 27911 48190 27920
rect 48148 27538 48176 27911
rect 48136 27532 48188 27538
rect 48136 27474 48188 27480
rect 48148 27130 48176 27474
rect 48136 27124 48188 27130
rect 48136 27066 48188 27072
rect 48136 26376 48188 26382
rect 48136 26318 48188 26324
rect 48148 25974 48176 26318
rect 48136 25968 48188 25974
rect 48134 25936 48136 25945
rect 48188 25936 48190 25945
rect 48134 25871 48190 25880
rect 48148 25845 48176 25871
rect 48136 24132 48188 24138
rect 48136 24074 48188 24080
rect 48148 23905 48176 24074
rect 48134 23896 48190 23905
rect 48134 23831 48136 23840
rect 48188 23831 48190 23840
rect 48136 23802 48188 23808
rect 48044 21888 48096 21894
rect 48042 21856 48044 21865
rect 48096 21856 48098 21865
rect 48042 21791 48098 21800
rect 48042 19816 48098 19825
rect 48042 19751 48098 19760
rect 48056 19718 48084 19751
rect 48044 19712 48096 19718
rect 48044 19654 48096 19660
rect 48044 18080 48096 18086
rect 48044 18022 48096 18028
rect 48056 17785 48084 18022
rect 48042 17776 48098 17785
rect 48042 17711 48098 17720
rect 48136 16108 48188 16114
rect 48136 16050 48188 16056
rect 48148 15745 48176 16050
rect 48134 15736 48190 15745
rect 48134 15671 48136 15680
rect 48188 15671 48190 15680
rect 48136 15642 48188 15648
rect 48044 13728 48096 13734
rect 48042 13696 48044 13705
rect 48096 13696 48098 13705
rect 48042 13631 48098 13640
rect 48136 11756 48188 11762
rect 48136 11698 48188 11704
rect 48148 11665 48176 11698
rect 48134 11656 48190 11665
rect 48134 11591 48190 11600
rect 48148 11354 48176 11591
rect 48136 11348 48188 11354
rect 48136 11290 48188 11296
rect 48044 9920 48096 9926
rect 48044 9862 48096 9868
rect 48056 9625 48084 9862
rect 48042 9616 48098 9625
rect 48042 9551 48098 9560
rect 47952 8084 48004 8090
rect 47952 8026 48004 8032
rect 48044 7812 48096 7818
rect 48044 7754 48096 7760
rect 48056 7585 48084 7754
rect 48042 7576 48098 7585
rect 48042 7511 48098 7520
rect 48044 5636 48096 5642
rect 48044 5578 48096 5584
rect 48056 5545 48084 5578
rect 48042 5536 48098 5545
rect 48042 5471 48098 5480
rect 47768 4140 47820 4146
rect 47768 4082 47820 4088
rect 47306 3632 47362 3641
rect 47306 3567 47308 3576
rect 47360 3567 47362 3576
rect 47308 3538 47360 3544
rect 46572 2984 46624 2990
rect 46570 2952 46572 2961
rect 46624 2952 46626 2961
rect 46570 2887 46626 2896
rect 45284 2644 45336 2650
rect 45284 2586 45336 2592
rect 44180 2576 44232 2582
rect 44180 2518 44232 2524
rect 45296 2446 45324 2586
rect 46584 2446 46612 2887
rect 47780 2446 47808 4082
rect 48042 3496 48098 3505
rect 48042 3431 48098 3440
rect 48320 3460 48372 3466
rect 48056 3398 48084 3431
rect 48320 3402 48372 3408
rect 48044 3392 48096 3398
rect 48044 3334 48096 3340
rect 48332 3058 48360 3402
rect 48320 3052 48372 3058
rect 48320 2994 48372 3000
rect 49608 3052 49660 3058
rect 49608 2994 49660 3000
rect 40040 2440 40092 2446
rect 40040 2382 40092 2388
rect 45284 2440 45336 2446
rect 45284 2382 45336 2388
rect 46572 2440 46624 2446
rect 46572 2382 46624 2388
rect 47768 2440 47820 2446
rect 47768 2382 47820 2388
rect 36084 2372 36136 2378
rect 36084 2314 36136 2320
rect 34152 2304 34204 2310
rect 34152 2246 34204 2252
rect 33968 1964 34020 1970
rect 33968 1906 34020 1912
rect 34164 800 34192 2246
rect 36096 800 36124 2314
rect 38016 2304 38068 2310
rect 38016 2246 38068 2252
rect 38028 800 38056 2246
rect 40052 1714 40080 2382
rect 43812 2372 43864 2378
rect 43812 2314 43864 2320
rect 40224 2304 40276 2310
rect 40224 2246 40276 2252
rect 41880 2304 41932 2310
rect 41880 2246 41932 2252
rect 42616 2304 42668 2310
rect 42616 2246 42668 2252
rect 40236 1902 40264 2246
rect 40224 1896 40276 1902
rect 40224 1838 40276 1844
rect 39960 1686 40080 1714
rect 39960 800 39988 1686
rect 41892 800 41920 2246
rect 42628 2038 42656 2246
rect 42616 2032 42668 2038
rect 42616 1974 42668 1980
rect 43824 800 43852 2314
rect 45744 2304 45796 2310
rect 45744 2246 45796 2252
rect 46848 2304 46900 2310
rect 46848 2246 46900 2252
rect 47676 2304 47728 2310
rect 47676 2246 47728 2252
rect 45756 800 45784 2246
rect 46860 1465 46888 2246
rect 46846 1456 46902 1465
rect 46846 1391 46902 1400
rect 47688 800 47716 2246
rect 49620 800 49648 2994
rect 18 0 74 800
rect 1306 0 1362 800
rect 3238 0 3294 800
rect 5170 0 5226 800
rect 7102 0 7158 800
rect 9034 0 9090 800
rect 10966 0 11022 800
rect 12898 0 12954 800
rect 14830 0 14886 800
rect 16762 0 16818 800
rect 18694 0 18750 800
rect 20626 0 20682 800
rect 22558 0 22614 800
rect 24490 0 24546 800
rect 26422 0 26478 800
rect 28354 0 28410 800
rect 30286 0 30342 800
rect 32218 0 32274 800
rect 34150 0 34206 800
rect 36082 0 36138 800
rect 38014 0 38070 800
rect 39946 0 40002 800
rect 41878 0 41934 800
rect 43810 0 43866 800
rect 45742 0 45798 800
rect 47674 0 47730 800
rect 49606 0 49662 800
<< via2 >>
rect 2778 48320 2834 48376
rect 1398 46280 1454 46336
rect 1398 44240 1454 44296
rect 1490 42200 1546 42256
rect 1582 40180 1638 40216
rect 1582 40160 1584 40180
rect 1584 40160 1636 40180
rect 1636 40160 1638 40180
rect 1582 38120 1638 38176
rect 1490 36080 1546 36136
rect 1582 34076 1584 34096
rect 1584 34076 1636 34096
rect 1636 34076 1638 34096
rect 1582 34040 1638 34076
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 2686 38936 2742 38992
rect 1674 33496 1730 33552
rect 1582 32020 1638 32056
rect 1582 32000 1584 32020
rect 1584 32000 1636 32020
rect 1636 32000 1638 32020
rect 1582 29960 1638 30016
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 8022 34040 8078 34096
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 2870 28056 2926 28112
rect 1490 27940 1546 27976
rect 1490 27920 1492 27940
rect 1492 27920 1544 27940
rect 1544 27920 1546 27940
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 1582 25916 1584 25936
rect 1584 25916 1636 25936
rect 1636 25916 1638 25936
rect 1582 25880 1638 25916
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 1490 23840 1546 23896
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 1582 21800 1638 21856
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 1858 19780 1914 19816
rect 1858 19760 1860 19780
rect 1860 19760 1912 19780
rect 1912 19760 1914 19780
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 1582 17756 1584 17776
rect 1584 17756 1636 17776
rect 1636 17756 1638 17776
rect 1582 17720 1638 17756
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 1582 15700 1638 15736
rect 1582 15680 1584 15700
rect 1584 15680 1636 15700
rect 1636 15680 1638 15700
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 1398 13640 1454 13696
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 1490 11620 1546 11656
rect 1490 11600 1492 11620
rect 1492 11600 1544 11620
rect 1544 11600 1546 11620
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 1582 9596 1584 9616
rect 1584 9596 1636 9616
rect 1636 9596 1638 9616
rect 1582 9560 1638 9596
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 1490 7520 1546 7576
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 1582 5480 1638 5536
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 1490 3440 1546 3496
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 1398 1400 1454 1456
rect 11886 45500 11888 45520
rect 11888 45500 11940 45520
rect 11940 45500 11942 45520
rect 11886 45464 11942 45500
rect 12714 46588 12716 46608
rect 12716 46588 12768 46608
rect 12768 46588 12770 46608
rect 12714 46552 12770 46588
rect 13818 44804 13874 44840
rect 13818 44784 13820 44804
rect 13820 44784 13872 44804
rect 13872 44784 13874 44804
rect 12990 43832 13046 43888
rect 12438 36760 12494 36816
rect 14646 44804 14702 44840
rect 14646 44784 14648 44804
rect 14648 44784 14700 44804
rect 14700 44784 14702 44804
rect 14462 44376 14518 44432
rect 11794 31728 11850 31784
rect 11978 2916 12034 2952
rect 11978 2896 11980 2916
rect 11980 2896 12032 2916
rect 12032 2896 12034 2916
rect 16486 43832 16542 43888
rect 18326 45484 18382 45520
rect 18326 45464 18328 45484
rect 18328 45464 18380 45484
rect 18380 45464 18382 45484
rect 17498 45328 17554 45384
rect 17498 44396 17554 44432
rect 17498 44376 17500 44396
rect 17500 44376 17552 44396
rect 17552 44376 17554 44396
rect 14002 41248 14058 41304
rect 15014 40468 15016 40488
rect 15016 40468 15068 40488
rect 15068 40468 15070 40488
rect 15014 40432 15070 40468
rect 14554 37712 14610 37768
rect 15474 40024 15530 40080
rect 18142 44396 18198 44432
rect 18142 44376 18144 44396
rect 18144 44376 18196 44396
rect 18196 44376 18198 44396
rect 18142 43832 18198 43888
rect 17866 43188 17868 43208
rect 17868 43188 17920 43208
rect 17920 43188 17922 43208
rect 17866 43152 17922 43188
rect 17866 40468 17868 40488
rect 17868 40468 17920 40488
rect 17920 40468 17922 40488
rect 17866 40432 17922 40468
rect 15106 37440 15162 37496
rect 15014 37204 15016 37224
rect 15016 37204 15068 37224
rect 15068 37204 15070 37224
rect 15014 37168 15070 37204
rect 15934 37304 15990 37360
rect 15842 36624 15898 36680
rect 17406 40024 17462 40080
rect 17038 37848 17094 37904
rect 16578 37576 16634 37632
rect 16118 36524 16120 36544
rect 16120 36524 16172 36544
rect 16172 36524 16174 36544
rect 16118 36488 16174 36524
rect 15382 31748 15438 31784
rect 15382 31728 15384 31748
rect 15384 31728 15436 31748
rect 15436 31728 15438 31748
rect 17590 38292 17592 38312
rect 17592 38292 17644 38312
rect 17644 38292 17646 38312
rect 17590 38256 17646 38292
rect 18694 43716 18750 43752
rect 18694 43696 18696 43716
rect 18696 43696 18748 43716
rect 18748 43696 18750 43716
rect 18326 43308 18382 43344
rect 18326 43288 18328 43308
rect 18328 43288 18380 43308
rect 18380 43288 18382 43308
rect 18602 41112 18658 41168
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19982 46436 20038 46472
rect 19982 46416 19984 46436
rect 19984 46416 20036 46436
rect 20036 46416 20038 46436
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19338 45464 19394 45520
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19430 41384 19486 41440
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19338 40160 19394 40216
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 20718 46572 20774 46608
rect 20718 46552 20720 46572
rect 20720 46552 20772 46572
rect 20772 46552 20774 46572
rect 21086 45328 21142 45384
rect 20718 44512 20774 44568
rect 20442 41132 20498 41168
rect 20442 41112 20444 41132
rect 20444 41112 20496 41132
rect 20496 41112 20498 41132
rect 21730 45872 21786 45928
rect 19430 39888 19486 39944
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 18510 38292 18512 38312
rect 18512 38292 18564 38312
rect 18564 38292 18566 38312
rect 18510 38256 18566 38292
rect 18694 37748 18696 37768
rect 18696 37748 18748 37768
rect 18748 37748 18750 37768
rect 18694 37712 18750 37748
rect 19614 38256 19670 38312
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19890 37612 19892 37632
rect 19892 37612 19944 37632
rect 19944 37612 19946 37632
rect 19890 37576 19946 37612
rect 18602 36624 18658 36680
rect 18786 35672 18842 35728
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19706 36780 19762 36816
rect 19706 36760 19708 36780
rect 19708 36760 19760 36780
rect 19760 36760 19762 36780
rect 19890 36624 19946 36680
rect 20718 40024 20774 40080
rect 20166 37068 20168 37088
rect 20168 37068 20220 37088
rect 20220 37068 20222 37088
rect 20166 37032 20222 37068
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 18418 33224 18474 33280
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19338 31592 19394 31648
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 20166 31728 20222 31784
rect 20534 36488 20590 36544
rect 20442 35944 20498 36000
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 20626 29588 20628 29608
rect 20628 29588 20680 29608
rect 20680 29588 20682 29608
rect 20626 29552 20682 29588
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 20350 27104 20406 27160
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 15198 2488 15254 2544
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 22006 42628 22062 42664
rect 22006 42608 22008 42628
rect 22008 42608 22060 42628
rect 22060 42608 22062 42628
rect 21086 41248 21142 41304
rect 21822 41248 21878 41304
rect 21822 40160 21878 40216
rect 22098 40432 22154 40488
rect 22374 41928 22430 41984
rect 22282 41112 22338 41168
rect 22006 39888 22062 39944
rect 21546 37032 21602 37088
rect 21454 36080 21510 36136
rect 21914 33224 21970 33280
rect 24490 45908 24492 45928
rect 24492 45908 24544 45928
rect 24544 45908 24546 45928
rect 24490 45872 24546 45908
rect 23294 37884 23296 37904
rect 23296 37884 23348 37904
rect 23348 37884 23350 37904
rect 23294 37848 23350 37884
rect 23018 35808 23074 35864
rect 23938 40160 23994 40216
rect 23846 38548 23902 38584
rect 23846 38528 23848 38548
rect 23848 38528 23900 38548
rect 23900 38528 23902 38548
rect 23846 37576 23902 37632
rect 24030 37712 24086 37768
rect 24674 40996 24730 41032
rect 24674 40976 24676 40996
rect 24676 40976 24728 40996
rect 24728 40976 24730 40996
rect 24030 36896 24086 36952
rect 24674 37984 24730 38040
rect 24306 37712 24362 37768
rect 24490 37324 24546 37360
rect 24490 37304 24492 37324
rect 24492 37304 24544 37324
rect 24544 37304 24546 37324
rect 24490 35536 24546 35592
rect 22006 31184 22062 31240
rect 20994 28056 21050 28112
rect 22282 28076 22338 28112
rect 22282 28056 22284 28076
rect 22284 28056 22336 28076
rect 22336 28056 22338 28076
rect 23018 31184 23074 31240
rect 25226 45600 25282 45656
rect 26238 45872 26294 45928
rect 25502 45328 25558 45384
rect 25410 35828 25466 35864
rect 26238 40060 26240 40080
rect 26240 40060 26292 40080
rect 26292 40060 26294 40080
rect 26238 40024 26294 40060
rect 25410 35808 25412 35828
rect 25412 35808 25464 35828
rect 25464 35808 25466 35828
rect 25042 34584 25098 34640
rect 25870 35536 25926 35592
rect 26698 37304 26754 37360
rect 27158 41792 27214 41848
rect 27342 41248 27398 41304
rect 27618 41656 27674 41712
rect 27526 41384 27582 41440
rect 27802 41520 27858 41576
rect 27434 38292 27436 38312
rect 27436 38292 27488 38312
rect 27488 38292 27490 38312
rect 27434 38256 27490 38292
rect 26974 37204 26976 37224
rect 26976 37204 27028 37224
rect 27028 37204 27030 37224
rect 26974 37168 27030 37204
rect 26882 36760 26938 36816
rect 27802 37440 27858 37496
rect 27066 34856 27122 34912
rect 28354 44512 28410 44568
rect 27894 35808 27950 35864
rect 27894 34856 27950 34912
rect 28446 37748 28448 37768
rect 28448 37748 28500 37768
rect 28500 37748 28502 37768
rect 28446 37712 28502 37748
rect 28630 41656 28686 41712
rect 30838 46960 30894 47016
rect 28906 41928 28962 41984
rect 29642 46416 29698 46472
rect 28906 41248 28962 41304
rect 28906 40432 28962 40488
rect 28630 37440 28686 37496
rect 28170 34856 28226 34912
rect 29182 38528 29238 38584
rect 29550 36624 29606 36680
rect 30286 45600 30342 45656
rect 30470 43288 30526 43344
rect 30378 41656 30434 41712
rect 30286 37712 30342 37768
rect 30102 37168 30158 37224
rect 30102 36488 30158 36544
rect 30010 35128 30066 35184
rect 29918 34720 29974 34776
rect 30378 36780 30434 36816
rect 30378 36760 30380 36780
rect 30380 36760 30432 36780
rect 30432 36760 30434 36780
rect 30562 37032 30618 37088
rect 30746 36352 30802 36408
rect 30930 37712 30986 37768
rect 31206 41676 31262 41712
rect 31206 41656 31208 41676
rect 31208 41656 31260 41676
rect 31260 41656 31262 41676
rect 31114 37304 31170 37360
rect 30930 34856 30986 34912
rect 30746 34604 30802 34640
rect 30746 34584 30748 34604
rect 30748 34584 30800 34604
rect 30800 34584 30802 34604
rect 31114 36896 31170 36952
rect 31758 40976 31814 41032
rect 32034 45348 32090 45384
rect 32034 45328 32036 45348
rect 32036 45328 32088 45348
rect 32088 45328 32090 45348
rect 32218 40568 32274 40624
rect 33230 43696 33286 43752
rect 33322 43152 33378 43208
rect 32494 41420 32496 41440
rect 32496 41420 32548 41440
rect 32548 41420 32550 41440
rect 32494 41384 32550 41420
rect 31390 38412 31446 38448
rect 31390 38392 31392 38412
rect 31392 38392 31444 38412
rect 31444 38392 31446 38412
rect 31482 37984 31538 38040
rect 31390 37032 31446 37088
rect 31298 36780 31354 36816
rect 31298 36760 31300 36780
rect 31300 36760 31352 36780
rect 31352 36760 31354 36780
rect 31206 34584 31262 34640
rect 30838 28076 30894 28112
rect 30838 28056 30840 28076
rect 30840 28056 30892 28076
rect 30892 28056 30894 28076
rect 31298 31628 31300 31648
rect 31300 31628 31352 31648
rect 31352 31628 31354 31648
rect 31298 31592 31354 31628
rect 31758 37848 31814 37904
rect 32494 40296 32550 40352
rect 32770 39888 32826 39944
rect 32770 39072 32826 39128
rect 32218 34856 32274 34912
rect 33506 40024 33562 40080
rect 32770 37868 32826 37904
rect 32770 37848 32772 37868
rect 32772 37848 32824 37868
rect 32824 37848 32826 37868
rect 32586 37168 32642 37224
rect 32402 35012 32458 35048
rect 32402 34992 32404 35012
rect 32404 34992 32456 35012
rect 32456 34992 32458 35012
rect 32402 34196 32458 34232
rect 32402 34176 32404 34196
rect 32404 34176 32456 34196
rect 32456 34176 32458 34196
rect 33966 38256 34022 38312
rect 33874 37032 33930 37088
rect 33874 36352 33930 36408
rect 33414 34740 33470 34776
rect 33414 34720 33416 34740
rect 33416 34720 33468 34740
rect 33468 34720 33470 34740
rect 33046 34176 33102 34232
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34702 45872 34758 45928
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34150 40296 34206 40352
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 35438 42744 35494 42800
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 36082 42744 36138 42800
rect 34334 39208 34390 39264
rect 34242 38528 34298 38584
rect 34518 37984 34574 38040
rect 34242 36896 34298 36952
rect 34150 36488 34206 36544
rect 34150 35808 34206 35864
rect 34518 36780 34574 36816
rect 34518 36760 34520 36780
rect 34520 36760 34572 36780
rect 34572 36760 34574 36780
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 35530 40024 35586 40080
rect 34794 39208 34850 39264
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34794 38528 34850 38584
rect 35438 38700 35440 38720
rect 35440 38700 35492 38720
rect 35492 38700 35494 38720
rect 35438 38664 35494 38700
rect 35438 38528 35494 38584
rect 35070 38256 35126 38312
rect 34794 37848 34850 37904
rect 34702 37168 34758 37224
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 36542 39380 36544 39400
rect 36544 39380 36596 39400
rect 36596 39380 36598 39400
rect 36542 39344 36598 39380
rect 35714 38528 35770 38584
rect 36082 38292 36084 38312
rect 36084 38292 36136 38312
rect 36136 38292 36138 38312
rect 36082 38256 36138 38292
rect 36358 38428 36360 38448
rect 36360 38428 36412 38448
rect 36412 38428 36414 38448
rect 36358 38392 36414 38428
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34794 34856 34850 34912
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 35530 35128 35586 35184
rect 48042 48320 48098 48376
rect 37278 42608 37334 42664
rect 37278 39888 37334 39944
rect 37554 38936 37610 38992
rect 37370 37340 37372 37360
rect 37372 37340 37424 37360
rect 37424 37340 37426 37360
rect 37370 37304 37426 37340
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 37002 34584 37058 34640
rect 36082 31592 36138 31648
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 37278 36644 37334 36680
rect 37278 36624 37280 36644
rect 37280 36624 37332 36644
rect 37332 36624 37334 36644
rect 37922 38528 37978 38584
rect 38106 38292 38108 38312
rect 38108 38292 38160 38312
rect 38160 38292 38162 38312
rect 38106 38256 38162 38292
rect 37738 33516 37794 33552
rect 37738 33496 37740 33516
rect 37740 33496 37792 33516
rect 37792 33496 37794 33516
rect 38566 38972 38568 38992
rect 38568 38972 38620 38992
rect 38620 38972 38622 38992
rect 38566 38936 38622 38972
rect 39118 39364 39174 39400
rect 39118 39344 39120 39364
rect 39120 39344 39172 39364
rect 39172 39344 39174 39364
rect 39762 39344 39818 39400
rect 39210 37732 39266 37768
rect 39210 37712 39212 37732
rect 39212 37712 39264 37732
rect 39264 37712 39266 37732
rect 39302 35808 39358 35864
rect 39854 37848 39910 37904
rect 39946 35012 40002 35048
rect 39946 34992 39948 35012
rect 39948 34992 40000 35012
rect 40000 34992 40002 35012
rect 39946 34040 40002 34096
rect 40774 34076 40776 34096
rect 40776 34076 40828 34096
rect 40828 34076 40830 34096
rect 40774 34040 40830 34076
rect 41602 39364 41658 39400
rect 41602 39344 41604 39364
rect 41604 39344 41656 39364
rect 41656 39344 41658 39364
rect 44178 36796 44180 36816
rect 44180 36796 44232 36816
rect 44232 36796 44234 36816
rect 44178 36760 44234 36796
rect 45466 35672 45522 35728
rect 47030 44376 47086 44432
rect 48134 46280 48190 46336
rect 48042 44240 48098 44296
rect 47306 40452 47362 40488
rect 47306 40432 47308 40452
rect 47308 40432 47360 40452
rect 47360 40432 47362 40452
rect 47582 37032 47638 37088
rect 48134 42200 48190 42256
rect 48042 40160 48098 40216
rect 48042 38156 48044 38176
rect 48044 38156 48096 38176
rect 48096 38156 48098 38176
rect 48042 38120 48098 38156
rect 47858 36100 47914 36136
rect 47858 36080 47860 36100
rect 47860 36080 47912 36100
rect 47912 36080 47914 36100
rect 48042 36100 48098 36136
rect 48042 36080 48044 36100
rect 48044 36080 48096 36100
rect 48096 36080 48098 36100
rect 46754 31184 46810 31240
rect 47858 13932 47914 13968
rect 47858 13912 47860 13932
rect 47860 13912 47912 13932
rect 47912 13912 47914 13932
rect 48134 34060 48190 34096
rect 48134 34040 48136 34060
rect 48136 34040 48188 34060
rect 48188 34040 48190 34060
rect 48042 32000 48098 32056
rect 48134 29960 48190 30016
rect 48134 27920 48190 27976
rect 48134 25916 48136 25936
rect 48136 25916 48188 25936
rect 48188 25916 48190 25936
rect 48134 25880 48190 25916
rect 48134 23860 48190 23896
rect 48134 23840 48136 23860
rect 48136 23840 48188 23860
rect 48188 23840 48190 23860
rect 48042 21836 48044 21856
rect 48044 21836 48096 21856
rect 48096 21836 48098 21856
rect 48042 21800 48098 21836
rect 48042 19760 48098 19816
rect 48042 17720 48098 17776
rect 48134 15700 48190 15736
rect 48134 15680 48136 15700
rect 48136 15680 48188 15700
rect 48188 15680 48190 15700
rect 48042 13676 48044 13696
rect 48044 13676 48096 13696
rect 48096 13676 48098 13696
rect 48042 13640 48098 13676
rect 48134 11600 48190 11656
rect 48042 9560 48098 9616
rect 48042 7520 48098 7576
rect 48042 5480 48098 5536
rect 47306 3596 47362 3632
rect 47306 3576 47308 3596
rect 47308 3576 47360 3596
rect 47360 3576 47362 3596
rect 46570 2932 46572 2952
rect 46572 2932 46624 2952
rect 46624 2932 46626 2952
rect 46570 2896 46626 2932
rect 48042 3440 48098 3496
rect 46846 1400 46902 1456
<< metal3 >>
rect 0 48378 800 48408
rect 2773 48378 2839 48381
rect 0 48376 2839 48378
rect 0 48320 2778 48376
rect 2834 48320 2839 48376
rect 0 48318 2839 48320
rect 0 48288 800 48318
rect 2773 48315 2839 48318
rect 48037 48378 48103 48381
rect 49200 48378 50000 48408
rect 48037 48376 50000 48378
rect 48037 48320 48042 48376
rect 48098 48320 50000 48376
rect 48037 48318 50000 48320
rect 48037 48315 48103 48318
rect 49200 48288 50000 48318
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 30833 47018 30899 47021
rect 30966 47018 30972 47020
rect 30833 47016 30972 47018
rect 30833 46960 30838 47016
rect 30894 46960 30972 47016
rect 30833 46958 30972 46960
rect 30833 46955 30899 46958
rect 30966 46956 30972 46958
rect 31036 46956 31042 47020
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 12709 46610 12775 46613
rect 20713 46610 20779 46613
rect 12709 46608 20779 46610
rect 12709 46552 12714 46608
rect 12770 46552 20718 46608
rect 20774 46552 20779 46608
rect 12709 46550 20779 46552
rect 12709 46547 12775 46550
rect 20713 46547 20779 46550
rect 19977 46474 20043 46477
rect 29637 46474 29703 46477
rect 19977 46472 29703 46474
rect 19977 46416 19982 46472
rect 20038 46416 29642 46472
rect 29698 46416 29703 46472
rect 19977 46414 29703 46416
rect 19977 46411 20043 46414
rect 29637 46411 29703 46414
rect 0 46338 800 46368
rect 1393 46338 1459 46341
rect 0 46336 1459 46338
rect 0 46280 1398 46336
rect 1454 46280 1459 46336
rect 0 46278 1459 46280
rect 0 46248 800 46278
rect 1393 46275 1459 46278
rect 48129 46338 48195 46341
rect 49200 46338 50000 46368
rect 48129 46336 50000 46338
rect 48129 46280 48134 46336
rect 48190 46280 50000 46336
rect 48129 46278 50000 46280
rect 48129 46275 48195 46278
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 49200 46248 50000 46278
rect 34930 46207 35246 46208
rect 21725 45930 21791 45933
rect 24485 45930 24551 45933
rect 26233 45930 26299 45933
rect 34697 45932 34763 45933
rect 34646 45930 34652 45932
rect 21725 45928 26299 45930
rect 21725 45872 21730 45928
rect 21786 45872 24490 45928
rect 24546 45872 26238 45928
rect 26294 45872 26299 45928
rect 21725 45870 26299 45872
rect 34606 45870 34652 45930
rect 34716 45928 34763 45932
rect 34758 45872 34763 45928
rect 21725 45867 21791 45870
rect 24485 45867 24551 45870
rect 26233 45867 26299 45870
rect 34646 45868 34652 45870
rect 34716 45868 34763 45872
rect 34697 45867 34763 45868
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 25221 45660 25287 45661
rect 25221 45656 25268 45660
rect 25332 45658 25338 45660
rect 25221 45600 25226 45656
rect 25221 45596 25268 45600
rect 25332 45598 25378 45658
rect 25332 45596 25338 45598
rect 30046 45596 30052 45660
rect 30116 45658 30122 45660
rect 30281 45658 30347 45661
rect 30116 45656 30347 45658
rect 30116 45600 30286 45656
rect 30342 45600 30347 45656
rect 30116 45598 30347 45600
rect 30116 45596 30122 45598
rect 25221 45595 25287 45596
rect 30281 45595 30347 45598
rect 11881 45522 11947 45525
rect 18321 45522 18387 45525
rect 19333 45522 19399 45525
rect 11881 45520 19399 45522
rect 11881 45464 11886 45520
rect 11942 45464 18326 45520
rect 18382 45464 19338 45520
rect 19394 45464 19399 45520
rect 11881 45462 19399 45464
rect 11881 45459 11947 45462
rect 18321 45459 18387 45462
rect 19333 45459 19399 45462
rect 17493 45386 17559 45389
rect 21081 45386 21147 45389
rect 17493 45384 21147 45386
rect 17493 45328 17498 45384
rect 17554 45328 21086 45384
rect 21142 45328 21147 45384
rect 17493 45326 21147 45328
rect 17493 45323 17559 45326
rect 21081 45323 21147 45326
rect 25497 45386 25563 45389
rect 32029 45386 32095 45389
rect 25497 45384 32095 45386
rect 25497 45328 25502 45384
rect 25558 45328 32034 45384
rect 32090 45328 32095 45384
rect 25497 45326 32095 45328
rect 25497 45323 25563 45326
rect 32029 45323 32095 45326
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 13813 44842 13879 44845
rect 14641 44842 14707 44845
rect 13813 44840 14707 44842
rect 13813 44784 13818 44840
rect 13874 44784 14646 44840
rect 14702 44784 14707 44840
rect 13813 44782 14707 44784
rect 13813 44779 13879 44782
rect 14641 44779 14707 44782
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 20713 44570 20779 44573
rect 28349 44570 28415 44573
rect 20713 44568 28415 44570
rect 20713 44512 20718 44568
rect 20774 44512 28354 44568
rect 28410 44512 28415 44568
rect 20713 44510 28415 44512
rect 20713 44507 20779 44510
rect 28349 44507 28415 44510
rect 14457 44434 14523 44437
rect 17493 44434 17559 44437
rect 14457 44432 17559 44434
rect 14457 44376 14462 44432
rect 14518 44376 17498 44432
rect 17554 44376 17559 44432
rect 14457 44374 17559 44376
rect 14457 44371 14523 44374
rect 17493 44371 17559 44374
rect 18137 44434 18203 44437
rect 47025 44434 47091 44437
rect 18137 44432 47091 44434
rect 18137 44376 18142 44432
rect 18198 44376 47030 44432
rect 47086 44376 47091 44432
rect 18137 44374 47091 44376
rect 18137 44371 18203 44374
rect 47025 44371 47091 44374
rect 0 44298 800 44328
rect 1393 44298 1459 44301
rect 0 44296 1459 44298
rect 0 44240 1398 44296
rect 1454 44240 1459 44296
rect 0 44238 1459 44240
rect 0 44208 800 44238
rect 1393 44235 1459 44238
rect 48037 44298 48103 44301
rect 49200 44298 50000 44328
rect 48037 44296 50000 44298
rect 48037 44240 48042 44296
rect 48098 44240 50000 44296
rect 48037 44238 50000 44240
rect 48037 44235 48103 44238
rect 49200 44208 50000 44238
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 12985 43890 13051 43893
rect 16481 43890 16547 43893
rect 18137 43890 18203 43893
rect 12985 43888 18203 43890
rect 12985 43832 12990 43888
rect 13046 43832 16486 43888
rect 16542 43832 18142 43888
rect 18198 43832 18203 43888
rect 12985 43830 18203 43832
rect 12985 43827 13051 43830
rect 16481 43827 16547 43830
rect 18137 43827 18203 43830
rect 18689 43754 18755 43757
rect 33225 43754 33291 43757
rect 18689 43752 33291 43754
rect 18689 43696 18694 43752
rect 18750 43696 33230 43752
rect 33286 43696 33291 43752
rect 18689 43694 33291 43696
rect 18689 43691 18755 43694
rect 33225 43691 33291 43694
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 18321 43346 18387 43349
rect 30465 43346 30531 43349
rect 18321 43344 30531 43346
rect 18321 43288 18326 43344
rect 18382 43288 30470 43344
rect 30526 43288 30531 43344
rect 18321 43286 30531 43288
rect 18321 43283 18387 43286
rect 30465 43283 30531 43286
rect 17861 43210 17927 43213
rect 33317 43210 33383 43213
rect 17861 43208 33383 43210
rect 17861 43152 17866 43208
rect 17922 43152 33322 43208
rect 33378 43152 33383 43208
rect 17861 43150 33383 43152
rect 17861 43147 17927 43150
rect 33317 43147 33383 43150
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 35433 42802 35499 42805
rect 36077 42802 36143 42805
rect 35433 42800 36143 42802
rect 35433 42744 35438 42800
rect 35494 42744 36082 42800
rect 36138 42744 36143 42800
rect 35433 42742 36143 42744
rect 35433 42739 35499 42742
rect 36077 42739 36143 42742
rect 22001 42666 22067 42669
rect 37273 42666 37339 42669
rect 22001 42664 37339 42666
rect 22001 42608 22006 42664
rect 22062 42608 37278 42664
rect 37334 42608 37339 42664
rect 22001 42606 37339 42608
rect 22001 42603 22067 42606
rect 37273 42603 37339 42606
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 0 42258 800 42288
rect 1485 42258 1551 42261
rect 0 42256 1551 42258
rect 0 42200 1490 42256
rect 1546 42200 1551 42256
rect 0 42198 1551 42200
rect 0 42168 800 42198
rect 1485 42195 1551 42198
rect 48129 42258 48195 42261
rect 49200 42258 50000 42288
rect 48129 42256 50000 42258
rect 48129 42200 48134 42256
rect 48190 42200 50000 42256
rect 48129 42198 50000 42200
rect 48129 42195 48195 42198
rect 49200 42168 50000 42198
rect 22369 41986 22435 41989
rect 28901 41986 28967 41989
rect 22369 41984 28967 41986
rect 22369 41928 22374 41984
rect 22430 41928 28906 41984
rect 28962 41928 28967 41984
rect 22369 41926 28967 41928
rect 22369 41923 22435 41926
rect 28901 41923 28967 41926
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 26734 41788 26740 41852
rect 26804 41850 26810 41852
rect 27153 41850 27219 41853
rect 26804 41848 27219 41850
rect 26804 41792 27158 41848
rect 27214 41792 27219 41848
rect 26804 41790 27219 41792
rect 26804 41788 26810 41790
rect 27153 41787 27219 41790
rect 27613 41714 27679 41717
rect 28625 41714 28691 41717
rect 30373 41716 30439 41717
rect 28758 41714 28764 41716
rect 27613 41712 28764 41714
rect 27613 41656 27618 41712
rect 27674 41656 28630 41712
rect 28686 41656 28764 41712
rect 27613 41654 28764 41656
rect 27613 41651 27679 41654
rect 28625 41651 28691 41654
rect 28758 41652 28764 41654
rect 28828 41652 28834 41716
rect 30373 41712 30420 41716
rect 30484 41714 30490 41716
rect 31201 41714 31267 41717
rect 35382 41714 35388 41716
rect 30373 41656 30378 41712
rect 30373 41652 30420 41656
rect 30484 41654 30530 41714
rect 30606 41712 35388 41714
rect 30606 41656 31206 41712
rect 31262 41656 35388 41712
rect 30606 41654 35388 41656
rect 30484 41652 30490 41654
rect 30373 41651 30439 41652
rect 27797 41578 27863 41581
rect 28390 41578 28396 41580
rect 27797 41576 28396 41578
rect 27797 41520 27802 41576
rect 27858 41520 28396 41576
rect 27797 41518 28396 41520
rect 27797 41515 27863 41518
rect 28390 41516 28396 41518
rect 28460 41578 28466 41580
rect 30606 41578 30666 41654
rect 31201 41651 31267 41654
rect 35382 41652 35388 41654
rect 35452 41652 35458 41716
rect 33358 41578 33364 41580
rect 28460 41518 30666 41578
rect 31710 41518 33364 41578
rect 28460 41516 28466 41518
rect 19425 41444 19491 41445
rect 19374 41442 19380 41444
rect 19334 41382 19380 41442
rect 19444 41440 19491 41444
rect 19486 41384 19491 41440
rect 19374 41380 19380 41382
rect 19444 41380 19491 41384
rect 19425 41379 19491 41380
rect 27521 41442 27587 41445
rect 31710 41442 31770 41518
rect 33358 41516 33364 41518
rect 33428 41516 33434 41580
rect 32489 41444 32555 41445
rect 27521 41440 31770 41442
rect 27521 41384 27526 41440
rect 27582 41384 31770 41440
rect 27521 41382 31770 41384
rect 27521 41379 27587 41382
rect 32438 41380 32444 41444
rect 32508 41442 32555 41444
rect 32508 41440 32600 41442
rect 32550 41384 32600 41440
rect 32508 41382 32600 41384
rect 32508 41380 32555 41382
rect 32489 41379 32555 41380
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 13997 41306 14063 41309
rect 21081 41306 21147 41309
rect 21817 41306 21883 41309
rect 13997 41304 16590 41306
rect 13997 41248 14002 41304
rect 14058 41248 16590 41304
rect 13997 41246 16590 41248
rect 13997 41243 14063 41246
rect 16530 41170 16590 41246
rect 21081 41304 21883 41306
rect 21081 41248 21086 41304
rect 21142 41248 21822 41304
rect 21878 41248 21883 41304
rect 21081 41246 21883 41248
rect 21081 41243 21147 41246
rect 21817 41243 21883 41246
rect 27337 41306 27403 41309
rect 28901 41306 28967 41309
rect 27337 41304 28967 41306
rect 27337 41248 27342 41304
rect 27398 41248 28906 41304
rect 28962 41248 28967 41304
rect 27337 41246 28967 41248
rect 27337 41243 27403 41246
rect 28901 41243 28967 41246
rect 18597 41170 18663 41173
rect 20437 41170 20503 41173
rect 22277 41170 22343 41173
rect 16530 41168 22343 41170
rect 16530 41112 18602 41168
rect 18658 41112 20442 41168
rect 20498 41112 22282 41168
rect 22338 41112 22343 41168
rect 16530 41110 22343 41112
rect 18597 41107 18663 41110
rect 20437 41107 20503 41110
rect 22277 41107 22343 41110
rect 24669 41034 24735 41037
rect 31753 41034 31819 41037
rect 24669 41032 31819 41034
rect 24669 40976 24674 41032
rect 24730 40976 31758 41032
rect 31814 40976 31819 41032
rect 24669 40974 31819 40976
rect 24669 40971 24735 40974
rect 31753 40971 31819 40974
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 32213 40626 32279 40629
rect 16070 40624 32279 40626
rect 16070 40568 32218 40624
rect 32274 40568 32279 40624
rect 16070 40566 32279 40568
rect 15009 40492 15075 40493
rect 14958 40428 14964 40492
rect 15028 40490 15075 40492
rect 16070 40490 16130 40566
rect 32213 40563 32279 40566
rect 15028 40488 16130 40490
rect 15070 40432 16130 40488
rect 15028 40430 16130 40432
rect 17861 40490 17927 40493
rect 22093 40490 22159 40493
rect 17861 40488 22159 40490
rect 17861 40432 17866 40488
rect 17922 40432 22098 40488
rect 22154 40432 22159 40488
rect 17861 40430 22159 40432
rect 15028 40428 15075 40430
rect 15009 40427 15075 40428
rect 17861 40427 17927 40430
rect 22093 40427 22159 40430
rect 28901 40490 28967 40493
rect 47301 40490 47367 40493
rect 28901 40488 47367 40490
rect 28901 40432 28906 40488
rect 28962 40432 47306 40488
rect 47362 40432 47367 40488
rect 28901 40430 47367 40432
rect 28901 40427 28967 40430
rect 47301 40427 47367 40430
rect 32489 40354 32555 40357
rect 34145 40354 34211 40357
rect 32489 40352 34346 40354
rect 32489 40296 32494 40352
rect 32550 40296 34150 40352
rect 34206 40296 34346 40352
rect 32489 40294 34346 40296
rect 32489 40291 32555 40294
rect 34145 40291 34211 40294
rect 19570 40288 19886 40289
rect 0 40218 800 40248
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 1577 40218 1643 40221
rect 0 40216 1643 40218
rect 0 40160 1582 40216
rect 1638 40160 1643 40216
rect 0 40158 1643 40160
rect 0 40128 800 40158
rect 1577 40155 1643 40158
rect 19333 40220 19399 40221
rect 19333 40216 19380 40220
rect 19444 40218 19450 40220
rect 21817 40218 21883 40221
rect 23933 40218 23999 40221
rect 19333 40160 19338 40216
rect 19333 40156 19380 40160
rect 19444 40158 19490 40218
rect 21817 40216 23999 40218
rect 21817 40160 21822 40216
rect 21878 40160 23938 40216
rect 23994 40160 23999 40216
rect 21817 40158 23999 40160
rect 19444 40156 19450 40158
rect 19333 40155 19399 40156
rect 21817 40155 21883 40158
rect 23933 40155 23999 40158
rect 15469 40082 15535 40085
rect 17401 40082 17467 40085
rect 15469 40080 17467 40082
rect 15469 40024 15474 40080
rect 15530 40024 17406 40080
rect 17462 40024 17467 40080
rect 15469 40022 17467 40024
rect 15469 40019 15535 40022
rect 17401 40019 17467 40022
rect 20713 40082 20779 40085
rect 26233 40082 26299 40085
rect 20713 40080 26299 40082
rect 20713 40024 20718 40080
rect 20774 40024 26238 40080
rect 26294 40024 26299 40080
rect 20713 40022 26299 40024
rect 20713 40019 20779 40022
rect 26233 40019 26299 40022
rect 33174 40020 33180 40084
rect 33244 40082 33250 40084
rect 33501 40082 33567 40085
rect 33244 40080 33567 40082
rect 33244 40024 33506 40080
rect 33562 40024 33567 40080
rect 33244 40022 33567 40024
rect 34286 40082 34346 40294
rect 48037 40218 48103 40221
rect 49200 40218 50000 40248
rect 48037 40216 50000 40218
rect 48037 40160 48042 40216
rect 48098 40160 50000 40216
rect 48037 40158 50000 40160
rect 48037 40155 48103 40158
rect 49200 40128 50000 40158
rect 35525 40082 35591 40085
rect 34286 40080 35591 40082
rect 34286 40024 35530 40080
rect 35586 40024 35591 40080
rect 34286 40022 35591 40024
rect 33244 40020 33250 40022
rect 33501 40019 33567 40022
rect 35525 40019 35591 40022
rect 19425 39946 19491 39949
rect 22001 39946 22067 39949
rect 19425 39944 22067 39946
rect 19425 39888 19430 39944
rect 19486 39888 22006 39944
rect 22062 39888 22067 39944
rect 19425 39886 22067 39888
rect 19425 39883 19491 39886
rect 22001 39883 22067 39886
rect 32765 39946 32831 39949
rect 37273 39946 37339 39949
rect 32765 39944 37339 39946
rect 32765 39888 32770 39944
rect 32826 39888 37278 39944
rect 37334 39888 37339 39944
rect 32765 39886 37339 39888
rect 32765 39883 32831 39886
rect 37273 39883 37339 39886
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 36537 39402 36603 39405
rect 39113 39402 39179 39405
rect 39757 39402 39823 39405
rect 41597 39402 41663 39405
rect 36537 39400 41663 39402
rect 36537 39344 36542 39400
rect 36598 39344 39118 39400
rect 39174 39344 39762 39400
rect 39818 39344 41602 39400
rect 41658 39344 41663 39400
rect 36537 39342 41663 39344
rect 36537 39339 36603 39342
rect 39113 39339 39179 39342
rect 39757 39339 39823 39342
rect 41597 39339 41663 39342
rect 34329 39266 34395 39269
rect 34789 39266 34855 39269
rect 34329 39264 34855 39266
rect 34329 39208 34334 39264
rect 34390 39208 34794 39264
rect 34850 39208 34855 39264
rect 34329 39206 34855 39208
rect 34329 39203 34395 39206
rect 34789 39203 34855 39206
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 26734 39068 26740 39132
rect 26804 39130 26810 39132
rect 32765 39130 32831 39133
rect 26804 39128 32831 39130
rect 26804 39072 32770 39128
rect 32826 39072 32831 39128
rect 26804 39070 32831 39072
rect 26804 39068 26810 39070
rect 32765 39067 32831 39070
rect 2681 38994 2747 38997
rect 37549 38994 37615 38997
rect 38561 38994 38627 38997
rect 2681 38992 38627 38994
rect 2681 38936 2686 38992
rect 2742 38936 37554 38992
rect 37610 38936 38566 38992
rect 38622 38936 38627 38992
rect 2681 38934 38627 38936
rect 2681 38931 2747 38934
rect 37549 38931 37615 38934
rect 38561 38931 38627 38934
rect 35433 38724 35499 38725
rect 35382 38660 35388 38724
rect 35452 38722 35499 38724
rect 35452 38720 35544 38722
rect 35494 38664 35544 38720
rect 35452 38662 35544 38664
rect 35452 38660 35499 38662
rect 35433 38659 35499 38660
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 23841 38586 23907 38589
rect 29177 38586 29243 38589
rect 23841 38584 29243 38586
rect 23841 38528 23846 38584
rect 23902 38528 29182 38584
rect 29238 38528 29243 38584
rect 23841 38526 29243 38528
rect 23841 38523 23907 38526
rect 29177 38523 29243 38526
rect 34237 38586 34303 38589
rect 34789 38586 34855 38589
rect 34237 38584 34855 38586
rect 34237 38528 34242 38584
rect 34298 38528 34794 38584
rect 34850 38528 34855 38584
rect 34237 38526 34855 38528
rect 34237 38523 34303 38526
rect 34789 38523 34855 38526
rect 35433 38586 35499 38589
rect 35709 38586 35775 38589
rect 37917 38586 37983 38589
rect 35433 38584 37983 38586
rect 35433 38528 35438 38584
rect 35494 38528 35714 38584
rect 35770 38528 37922 38584
rect 37978 38528 37983 38584
rect 35433 38526 37983 38528
rect 35433 38523 35499 38526
rect 35709 38523 35775 38526
rect 37917 38523 37983 38526
rect 31385 38450 31451 38453
rect 36353 38450 36419 38453
rect 31385 38448 36419 38450
rect 31385 38392 31390 38448
rect 31446 38392 36358 38448
rect 36414 38392 36419 38448
rect 31385 38390 36419 38392
rect 31385 38387 31451 38390
rect 36353 38387 36419 38390
rect 17585 38314 17651 38317
rect 18505 38314 18571 38317
rect 17585 38312 18571 38314
rect 17585 38256 17590 38312
rect 17646 38256 18510 38312
rect 18566 38256 18571 38312
rect 17585 38254 18571 38256
rect 17585 38251 17651 38254
rect 18505 38251 18571 38254
rect 19609 38314 19675 38317
rect 27429 38314 27495 38317
rect 19609 38312 27495 38314
rect 19609 38256 19614 38312
rect 19670 38256 27434 38312
rect 27490 38256 27495 38312
rect 19609 38254 27495 38256
rect 19609 38251 19675 38254
rect 27429 38251 27495 38254
rect 33961 38314 34027 38317
rect 35065 38314 35131 38317
rect 33961 38312 35131 38314
rect 33961 38256 33966 38312
rect 34022 38256 35070 38312
rect 35126 38256 35131 38312
rect 33961 38254 35131 38256
rect 33961 38251 34027 38254
rect 35065 38251 35131 38254
rect 36077 38314 36143 38317
rect 38101 38314 38167 38317
rect 36077 38312 38167 38314
rect 36077 38256 36082 38312
rect 36138 38256 38106 38312
rect 38162 38256 38167 38312
rect 36077 38254 38167 38256
rect 36077 38251 36143 38254
rect 38101 38251 38167 38254
rect 0 38178 800 38208
rect 1577 38178 1643 38181
rect 0 38176 1643 38178
rect 0 38120 1582 38176
rect 1638 38120 1643 38176
rect 0 38118 1643 38120
rect 0 38088 800 38118
rect 1577 38115 1643 38118
rect 48037 38178 48103 38181
rect 49200 38178 50000 38208
rect 48037 38176 50000 38178
rect 48037 38120 48042 38176
rect 48098 38120 50000 38176
rect 48037 38118 50000 38120
rect 48037 38115 48103 38118
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 49200 38088 50000 38118
rect 19570 38047 19886 38048
rect 24669 38042 24735 38045
rect 31477 38042 31543 38045
rect 34513 38042 34579 38045
rect 24669 38040 34579 38042
rect 24669 37984 24674 38040
rect 24730 37984 31482 38040
rect 31538 37984 34518 38040
rect 34574 37984 34579 38040
rect 24669 37982 34579 37984
rect 24669 37979 24735 37982
rect 31477 37979 31543 37982
rect 34513 37979 34579 37982
rect 17033 37906 17099 37909
rect 23289 37906 23355 37909
rect 17033 37904 23355 37906
rect 17033 37848 17038 37904
rect 17094 37848 23294 37904
rect 23350 37848 23355 37904
rect 17033 37846 23355 37848
rect 17033 37843 17099 37846
rect 23289 37843 23355 37846
rect 31753 37906 31819 37909
rect 32765 37906 32831 37909
rect 34789 37906 34855 37909
rect 39849 37906 39915 37909
rect 31753 37904 39915 37906
rect 31753 37848 31758 37904
rect 31814 37848 32770 37904
rect 32826 37848 34794 37904
rect 34850 37848 39854 37904
rect 39910 37848 39915 37904
rect 31753 37846 39915 37848
rect 31753 37843 31819 37846
rect 32765 37843 32831 37846
rect 34789 37843 34855 37846
rect 39849 37843 39915 37846
rect 14549 37770 14615 37773
rect 18689 37770 18755 37773
rect 14549 37768 18755 37770
rect 14549 37712 14554 37768
rect 14610 37712 18694 37768
rect 18750 37712 18755 37768
rect 14549 37710 18755 37712
rect 14549 37707 14615 37710
rect 18689 37707 18755 37710
rect 24025 37770 24091 37773
rect 24301 37770 24367 37773
rect 28441 37772 28507 37773
rect 24025 37768 24367 37770
rect 24025 37712 24030 37768
rect 24086 37712 24306 37768
rect 24362 37712 24367 37768
rect 24025 37710 24367 37712
rect 24025 37707 24091 37710
rect 24301 37707 24367 37710
rect 28390 37708 28396 37772
rect 28460 37770 28507 37772
rect 30281 37770 30347 37773
rect 30925 37770 30991 37773
rect 39205 37770 39271 37773
rect 28460 37768 28552 37770
rect 28502 37712 28552 37768
rect 28460 37710 28552 37712
rect 30281 37768 39271 37770
rect 30281 37712 30286 37768
rect 30342 37712 30930 37768
rect 30986 37712 39210 37768
rect 39266 37712 39271 37768
rect 30281 37710 39271 37712
rect 28460 37708 28507 37710
rect 28441 37707 28507 37708
rect 30281 37707 30347 37710
rect 30925 37707 30991 37710
rect 39205 37707 39271 37710
rect 16573 37634 16639 37637
rect 19885 37634 19951 37637
rect 23841 37634 23907 37637
rect 16573 37632 23907 37634
rect 16573 37576 16578 37632
rect 16634 37576 19890 37632
rect 19946 37576 23846 37632
rect 23902 37576 23907 37632
rect 16573 37574 23907 37576
rect 16573 37571 16639 37574
rect 19885 37571 19951 37574
rect 23841 37571 23907 37574
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 15101 37498 15167 37501
rect 27797 37498 27863 37501
rect 28625 37498 28691 37501
rect 15101 37496 28691 37498
rect 15101 37440 15106 37496
rect 15162 37440 27802 37496
rect 27858 37440 28630 37496
rect 28686 37440 28691 37496
rect 15101 37438 28691 37440
rect 15101 37435 15167 37438
rect 27797 37435 27863 37438
rect 28625 37435 28691 37438
rect 15929 37362 15995 37365
rect 24485 37362 24551 37365
rect 15929 37360 24551 37362
rect 15929 37304 15934 37360
rect 15990 37304 24490 37360
rect 24546 37304 24551 37360
rect 15929 37302 24551 37304
rect 15929 37299 15995 37302
rect 24485 37299 24551 37302
rect 26693 37362 26759 37365
rect 31109 37362 31175 37365
rect 37365 37362 37431 37365
rect 26693 37360 37431 37362
rect 26693 37304 26698 37360
rect 26754 37304 31114 37360
rect 31170 37304 37370 37360
rect 37426 37304 37431 37360
rect 26693 37302 37431 37304
rect 26693 37299 26759 37302
rect 15009 37226 15075 37229
rect 26969 37226 27035 37229
rect 28390 37226 28396 37228
rect 15009 37224 28396 37226
rect 15009 37168 15014 37224
rect 15070 37168 26974 37224
rect 27030 37168 28396 37224
rect 15009 37166 28396 37168
rect 15009 37163 15075 37166
rect 26969 37163 27035 37166
rect 28390 37164 28396 37166
rect 28460 37164 28466 37228
rect 30097 37226 30163 37229
rect 30238 37228 30298 37302
rect 31109 37299 31175 37302
rect 37365 37299 37431 37302
rect 30230 37226 30236 37228
rect 30097 37224 30236 37226
rect 30097 37168 30102 37224
rect 30158 37168 30236 37224
rect 30097 37166 30236 37168
rect 30097 37163 30163 37166
rect 30230 37164 30236 37166
rect 30300 37164 30306 37228
rect 32581 37226 32647 37229
rect 34697 37226 34763 37229
rect 32581 37224 34763 37226
rect 32581 37168 32586 37224
rect 32642 37168 34702 37224
rect 34758 37168 34763 37224
rect 32581 37166 34763 37168
rect 32581 37163 32647 37166
rect 34697 37163 34763 37166
rect 20161 37090 20227 37093
rect 21541 37090 21607 37093
rect 20161 37088 21607 37090
rect 20161 37032 20166 37088
rect 20222 37032 21546 37088
rect 21602 37032 21607 37088
rect 20161 37030 21607 37032
rect 20161 37027 20227 37030
rect 21541 37027 21607 37030
rect 30557 37090 30623 37093
rect 31385 37090 31451 37093
rect 33869 37090 33935 37093
rect 47577 37090 47643 37093
rect 30557 37088 47643 37090
rect 30557 37032 30562 37088
rect 30618 37032 31390 37088
rect 31446 37032 33874 37088
rect 33930 37032 47582 37088
rect 47638 37032 47643 37088
rect 30557 37030 47643 37032
rect 30557 37027 30623 37030
rect 31385 37027 31451 37030
rect 33869 37027 33935 37030
rect 47577 37027 47643 37030
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 24025 36954 24091 36957
rect 31109 36954 31175 36957
rect 34237 36954 34303 36957
rect 24025 36952 31175 36954
rect 24025 36896 24030 36952
rect 24086 36896 31114 36952
rect 31170 36896 31175 36952
rect 24025 36894 31175 36896
rect 24025 36891 24091 36894
rect 31109 36891 31175 36894
rect 31296 36952 34303 36954
rect 31296 36896 34242 36952
rect 34298 36896 34303 36952
rect 31296 36894 34303 36896
rect 31296 36821 31356 36894
rect 34237 36891 34303 36894
rect 12433 36818 12499 36821
rect 19701 36818 19767 36821
rect 12433 36816 19767 36818
rect 12433 36760 12438 36816
rect 12494 36760 19706 36816
rect 19762 36760 19767 36816
rect 12433 36758 19767 36760
rect 12433 36755 12499 36758
rect 19701 36755 19767 36758
rect 26877 36818 26943 36821
rect 30373 36818 30439 36821
rect 31293 36818 31359 36821
rect 26877 36816 31359 36818
rect 26877 36760 26882 36816
rect 26938 36760 30378 36816
rect 30434 36760 31298 36816
rect 31354 36760 31359 36816
rect 26877 36758 31359 36760
rect 26877 36755 26943 36758
rect 30373 36755 30439 36758
rect 31293 36755 31359 36758
rect 34513 36818 34579 36821
rect 44173 36818 44239 36821
rect 34513 36816 44239 36818
rect 34513 36760 34518 36816
rect 34574 36760 44178 36816
rect 44234 36760 44239 36816
rect 34513 36758 44239 36760
rect 34513 36755 34579 36758
rect 44173 36755 44239 36758
rect 15837 36682 15903 36685
rect 18597 36682 18663 36685
rect 19885 36682 19951 36685
rect 15837 36680 19951 36682
rect 15837 36624 15842 36680
rect 15898 36624 18602 36680
rect 18658 36624 19890 36680
rect 19946 36624 19951 36680
rect 15837 36622 19951 36624
rect 15837 36619 15903 36622
rect 18597 36619 18663 36622
rect 19885 36619 19951 36622
rect 29545 36682 29611 36685
rect 32438 36682 32444 36684
rect 29545 36680 32444 36682
rect 29545 36624 29550 36680
rect 29606 36624 32444 36680
rect 29545 36622 32444 36624
rect 29545 36619 29611 36622
rect 32438 36620 32444 36622
rect 32508 36682 32514 36684
rect 37273 36682 37339 36685
rect 32508 36680 37339 36682
rect 32508 36624 37278 36680
rect 37334 36624 37339 36680
rect 32508 36622 37339 36624
rect 32508 36620 32514 36622
rect 37273 36619 37339 36622
rect 16113 36546 16179 36549
rect 20529 36546 20595 36549
rect 16113 36544 20595 36546
rect 16113 36488 16118 36544
rect 16174 36488 20534 36544
rect 20590 36488 20595 36544
rect 16113 36486 20595 36488
rect 16113 36483 16179 36486
rect 20529 36483 20595 36486
rect 30097 36546 30163 36549
rect 34145 36546 34211 36549
rect 30097 36544 34211 36546
rect 30097 36488 30102 36544
rect 30158 36488 34150 36544
rect 34206 36488 34211 36544
rect 30097 36486 34211 36488
rect 30097 36483 30163 36486
rect 34145 36483 34211 36486
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 30741 36410 30807 36413
rect 33869 36410 33935 36413
rect 30741 36408 33935 36410
rect 30741 36352 30746 36408
rect 30802 36352 33874 36408
rect 33930 36352 33935 36408
rect 30741 36350 33935 36352
rect 30741 36347 30807 36350
rect 33869 36347 33935 36350
rect 0 36138 800 36168
rect 1485 36138 1551 36141
rect 0 36136 1551 36138
rect 0 36080 1490 36136
rect 1546 36080 1551 36136
rect 0 36078 1551 36080
rect 0 36048 800 36078
rect 1485 36075 1551 36078
rect 21449 36138 21515 36141
rect 47853 36138 47919 36141
rect 21449 36136 47919 36138
rect 21449 36080 21454 36136
rect 21510 36080 47858 36136
rect 47914 36080 47919 36136
rect 21449 36078 47919 36080
rect 21449 36075 21515 36078
rect 47853 36075 47919 36078
rect 48037 36138 48103 36141
rect 49200 36138 50000 36168
rect 48037 36136 50000 36138
rect 48037 36080 48042 36136
rect 48098 36080 50000 36136
rect 48037 36078 50000 36080
rect 48037 36075 48103 36078
rect 49200 36048 50000 36078
rect 20437 36004 20503 36005
rect 20437 36002 20484 36004
rect 20392 36000 20484 36002
rect 20392 35944 20442 36000
rect 20392 35942 20484 35944
rect 20437 35940 20484 35942
rect 20548 35940 20554 36004
rect 20437 35939 20503 35940
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 23013 35866 23079 35869
rect 25262 35866 25268 35868
rect 23013 35864 25268 35866
rect 23013 35808 23018 35864
rect 23074 35808 25268 35864
rect 23013 35806 25268 35808
rect 23013 35803 23079 35806
rect 25262 35804 25268 35806
rect 25332 35804 25338 35868
rect 25405 35866 25471 35869
rect 27889 35866 27955 35869
rect 25405 35864 27955 35866
rect 25405 35808 25410 35864
rect 25466 35808 27894 35864
rect 27950 35808 27955 35864
rect 25405 35806 27955 35808
rect 25405 35803 25471 35806
rect 27889 35803 27955 35806
rect 34145 35866 34211 35869
rect 39297 35866 39363 35869
rect 34145 35864 39363 35866
rect 34145 35808 34150 35864
rect 34206 35808 39302 35864
rect 39358 35808 39363 35864
rect 34145 35806 39363 35808
rect 34145 35803 34211 35806
rect 39297 35803 39363 35806
rect 18781 35730 18847 35733
rect 45461 35730 45527 35733
rect 18781 35728 45527 35730
rect 18781 35672 18786 35728
rect 18842 35672 45466 35728
rect 45522 35672 45527 35728
rect 18781 35670 45527 35672
rect 18781 35667 18847 35670
rect 45461 35667 45527 35670
rect 24485 35594 24551 35597
rect 25865 35594 25931 35597
rect 24485 35592 25931 35594
rect 24485 35536 24490 35592
rect 24546 35536 25870 35592
rect 25926 35536 25931 35592
rect 24485 35534 25931 35536
rect 24485 35531 24551 35534
rect 25865 35531 25931 35534
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 30005 35186 30071 35189
rect 35525 35186 35591 35189
rect 30005 35184 35591 35186
rect 30005 35128 30010 35184
rect 30066 35128 35530 35184
rect 35586 35128 35591 35184
rect 30005 35126 35591 35128
rect 30005 35123 30071 35126
rect 35525 35123 35591 35126
rect 32397 35050 32463 35053
rect 39941 35050 40007 35053
rect 32397 35048 40007 35050
rect 32397 34992 32402 35048
rect 32458 34992 39946 35048
rect 40002 34992 40007 35048
rect 32397 34990 40007 34992
rect 32397 34987 32463 34990
rect 39941 34987 40007 34990
rect 27061 34914 27127 34917
rect 27889 34914 27955 34917
rect 28165 34914 28231 34917
rect 30925 34914 30991 34917
rect 32213 34914 32279 34917
rect 34789 34914 34855 34917
rect 27061 34912 34855 34914
rect 27061 34856 27066 34912
rect 27122 34856 27894 34912
rect 27950 34856 28170 34912
rect 28226 34856 30930 34912
rect 30986 34856 32218 34912
rect 32274 34856 34794 34912
rect 34850 34856 34855 34912
rect 27061 34854 34855 34856
rect 27061 34851 27127 34854
rect 27889 34851 27955 34854
rect 28165 34851 28231 34854
rect 30925 34851 30991 34854
rect 32213 34851 32279 34854
rect 34789 34851 34855 34854
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 29913 34778 29979 34781
rect 33409 34780 33475 34781
rect 30414 34778 30420 34780
rect 29913 34776 30420 34778
rect 29913 34720 29918 34776
rect 29974 34720 30420 34776
rect 29913 34718 30420 34720
rect 29913 34715 29979 34718
rect 30414 34716 30420 34718
rect 30484 34716 30490 34780
rect 33358 34716 33364 34780
rect 33428 34778 33475 34780
rect 33428 34776 33520 34778
rect 33470 34720 33520 34776
rect 33428 34718 33520 34720
rect 33428 34716 33475 34718
rect 33409 34715 33475 34716
rect 25037 34642 25103 34645
rect 30046 34642 30052 34644
rect 25037 34640 30052 34642
rect 25037 34584 25042 34640
rect 25098 34584 30052 34640
rect 25037 34582 30052 34584
rect 25037 34579 25103 34582
rect 30046 34580 30052 34582
rect 30116 34580 30122 34644
rect 30741 34642 30807 34645
rect 31201 34642 31267 34645
rect 36997 34642 37063 34645
rect 30741 34640 37063 34642
rect 30741 34584 30746 34640
rect 30802 34584 31206 34640
rect 31262 34584 37002 34640
rect 37058 34584 37063 34640
rect 30741 34582 37063 34584
rect 30741 34579 30807 34582
rect 31201 34579 31267 34582
rect 36997 34579 37063 34582
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 32397 34234 32463 34237
rect 33041 34234 33107 34237
rect 33174 34234 33180 34236
rect 32397 34232 33180 34234
rect 32397 34176 32402 34232
rect 32458 34176 33046 34232
rect 33102 34176 33180 34232
rect 32397 34174 33180 34176
rect 32397 34171 32463 34174
rect 33041 34171 33107 34174
rect 33174 34172 33180 34174
rect 33244 34172 33250 34236
rect 0 34098 800 34128
rect 1577 34098 1643 34101
rect 0 34096 1643 34098
rect 0 34040 1582 34096
rect 1638 34040 1643 34096
rect 0 34038 1643 34040
rect 0 34008 800 34038
rect 1577 34035 1643 34038
rect 8017 34098 8083 34101
rect 39941 34098 40007 34101
rect 40769 34098 40835 34101
rect 8017 34096 40835 34098
rect 8017 34040 8022 34096
rect 8078 34040 39946 34096
rect 40002 34040 40774 34096
rect 40830 34040 40835 34096
rect 8017 34038 40835 34040
rect 8017 34035 8083 34038
rect 39941 34035 40007 34038
rect 40769 34035 40835 34038
rect 48129 34098 48195 34101
rect 49200 34098 50000 34128
rect 48129 34096 50000 34098
rect 48129 34040 48134 34096
rect 48190 34040 50000 34096
rect 48129 34038 50000 34040
rect 48129 34035 48195 34038
rect 49200 34008 50000 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 1669 33554 1735 33557
rect 37733 33554 37799 33557
rect 1669 33552 37799 33554
rect 1669 33496 1674 33552
rect 1730 33496 37738 33552
rect 37794 33496 37799 33552
rect 1669 33494 37799 33496
rect 1669 33491 1735 33494
rect 37733 33491 37799 33494
rect 18413 33282 18479 33285
rect 21909 33282 21975 33285
rect 18413 33280 21975 33282
rect 18413 33224 18418 33280
rect 18474 33224 21914 33280
rect 21970 33224 21975 33280
rect 18413 33222 21975 33224
rect 18413 33219 18479 33222
rect 21909 33219 21975 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 0 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1577 32058 1643 32061
rect 0 32056 1643 32058
rect 0 32000 1582 32056
rect 1638 32000 1643 32056
rect 0 31998 1643 32000
rect 0 31968 800 31998
rect 1577 31995 1643 31998
rect 48037 32058 48103 32061
rect 49200 32058 50000 32088
rect 48037 32056 50000 32058
rect 48037 32000 48042 32056
rect 48098 32000 50000 32056
rect 48037 31998 50000 32000
rect 48037 31995 48103 31998
rect 49200 31968 50000 31998
rect 11789 31786 11855 31789
rect 15377 31786 15443 31789
rect 11789 31784 15443 31786
rect 11789 31728 11794 31784
rect 11850 31728 15382 31784
rect 15438 31728 15443 31784
rect 11789 31726 15443 31728
rect 11789 31723 11855 31726
rect 15377 31723 15443 31726
rect 19006 31724 19012 31788
rect 19076 31786 19082 31788
rect 20161 31786 20227 31789
rect 19076 31784 20227 31786
rect 19076 31728 20166 31784
rect 20222 31728 20227 31784
rect 19076 31726 20227 31728
rect 19076 31724 19082 31726
rect 20161 31723 20227 31726
rect 19006 31588 19012 31652
rect 19076 31650 19082 31652
rect 19333 31650 19399 31653
rect 19076 31648 19399 31650
rect 19076 31592 19338 31648
rect 19394 31592 19399 31648
rect 19076 31590 19399 31592
rect 19076 31588 19082 31590
rect 19333 31587 19399 31590
rect 31293 31650 31359 31653
rect 36077 31650 36143 31653
rect 31293 31648 36143 31650
rect 31293 31592 31298 31648
rect 31354 31592 36082 31648
rect 36138 31592 36143 31648
rect 31293 31590 36143 31592
rect 31293 31587 31359 31590
rect 36077 31587 36143 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 22001 31242 22067 31245
rect 23013 31242 23079 31245
rect 46749 31242 46815 31245
rect 22001 31240 46815 31242
rect 22001 31184 22006 31240
rect 22062 31184 23018 31240
rect 23074 31184 46754 31240
rect 46810 31184 46815 31240
rect 22001 31182 46815 31184
rect 22001 31179 22067 31182
rect 23013 31179 23079 31182
rect 46749 31179 46815 31182
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 0 30018 800 30048
rect 1577 30018 1643 30021
rect 0 30016 1643 30018
rect 0 29960 1582 30016
rect 1638 29960 1643 30016
rect 0 29958 1643 29960
rect 0 29928 800 29958
rect 1577 29955 1643 29958
rect 48129 30018 48195 30021
rect 49200 30018 50000 30048
rect 48129 30016 50000 30018
rect 48129 29960 48134 30016
rect 48190 29960 50000 30016
rect 48129 29958 50000 29960
rect 48129 29955 48195 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 49200 29928 50000 29958
rect 34930 29887 35246 29888
rect 20621 29610 20687 29613
rect 34646 29610 34652 29612
rect 20621 29608 34652 29610
rect 20621 29552 20626 29608
rect 20682 29552 34652 29608
rect 20621 29550 34652 29552
rect 20621 29547 20687 29550
rect 34646 29548 34652 29550
rect 34716 29548 34722 29612
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 2865 28114 2931 28117
rect 20989 28114 21055 28117
rect 22277 28114 22343 28117
rect 2865 28112 22343 28114
rect 2865 28056 2870 28112
rect 2926 28056 20994 28112
rect 21050 28056 22282 28112
rect 22338 28056 22343 28112
rect 2865 28054 22343 28056
rect 2865 28051 2931 28054
rect 20989 28051 21055 28054
rect 22277 28051 22343 28054
rect 30230 28052 30236 28116
rect 30300 28114 30306 28116
rect 30833 28114 30899 28117
rect 30300 28112 30899 28114
rect 30300 28056 30838 28112
rect 30894 28056 30899 28112
rect 30300 28054 30899 28056
rect 30300 28052 30306 28054
rect 30833 28051 30899 28054
rect 0 27978 800 28008
rect 1485 27978 1551 27981
rect 0 27976 1551 27978
rect 0 27920 1490 27976
rect 1546 27920 1551 27976
rect 0 27918 1551 27920
rect 0 27888 800 27918
rect 1485 27915 1551 27918
rect 48129 27978 48195 27981
rect 49200 27978 50000 28008
rect 48129 27976 50000 27978
rect 48129 27920 48134 27976
rect 48190 27920 50000 27976
rect 48129 27918 50000 27920
rect 48129 27915 48195 27918
rect 49200 27888 50000 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 20345 27162 20411 27165
rect 20478 27162 20484 27164
rect 20345 27160 20484 27162
rect 20345 27104 20350 27160
rect 20406 27104 20484 27160
rect 20345 27102 20484 27104
rect 20345 27099 20411 27102
rect 20478 27100 20484 27102
rect 20548 27100 20554 27164
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 0 25938 800 25968
rect 1577 25938 1643 25941
rect 0 25936 1643 25938
rect 0 25880 1582 25936
rect 1638 25880 1643 25936
rect 0 25878 1643 25880
rect 0 25848 800 25878
rect 1577 25875 1643 25878
rect 48129 25938 48195 25941
rect 49200 25938 50000 25968
rect 48129 25936 50000 25938
rect 48129 25880 48134 25936
rect 48190 25880 50000 25936
rect 48129 25878 50000 25880
rect 48129 25875 48195 25878
rect 49200 25848 50000 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 0 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 1485 23898 1551 23901
rect 0 23896 1551 23898
rect 0 23840 1490 23896
rect 1546 23840 1551 23896
rect 0 23838 1551 23840
rect 0 23808 800 23838
rect 1485 23835 1551 23838
rect 48129 23898 48195 23901
rect 49200 23898 50000 23928
rect 48129 23896 50000 23898
rect 48129 23840 48134 23896
rect 48190 23840 50000 23896
rect 48129 23838 50000 23840
rect 48129 23835 48195 23838
rect 49200 23808 50000 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 0 21858 800 21888
rect 1577 21858 1643 21861
rect 0 21856 1643 21858
rect 0 21800 1582 21856
rect 1638 21800 1643 21856
rect 0 21798 1643 21800
rect 0 21768 800 21798
rect 1577 21795 1643 21798
rect 48037 21858 48103 21861
rect 49200 21858 50000 21888
rect 48037 21856 50000 21858
rect 48037 21800 48042 21856
rect 48098 21800 50000 21856
rect 48037 21798 50000 21800
rect 48037 21795 48103 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 49200 21768 50000 21798
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 0 19818 800 19848
rect 1853 19818 1919 19821
rect 0 19816 1919 19818
rect 0 19760 1858 19816
rect 1914 19760 1919 19816
rect 0 19758 1919 19760
rect 0 19728 800 19758
rect 1853 19755 1919 19758
rect 48037 19818 48103 19821
rect 49200 19818 50000 19848
rect 48037 19816 50000 19818
rect 48037 19760 48042 19816
rect 48098 19760 50000 19816
rect 48037 19758 50000 19760
rect 48037 19755 48103 19758
rect 49200 19728 50000 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 0 17778 800 17808
rect 1577 17778 1643 17781
rect 0 17776 1643 17778
rect 0 17720 1582 17776
rect 1638 17720 1643 17776
rect 0 17718 1643 17720
rect 0 17688 800 17718
rect 1577 17715 1643 17718
rect 48037 17778 48103 17781
rect 49200 17778 50000 17808
rect 48037 17776 50000 17778
rect 48037 17720 48042 17776
rect 48098 17720 50000 17776
rect 48037 17718 50000 17720
rect 48037 17715 48103 17718
rect 49200 17688 50000 17718
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 0 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1577 15738 1643 15741
rect 0 15736 1643 15738
rect 0 15680 1582 15736
rect 1638 15680 1643 15736
rect 0 15678 1643 15680
rect 0 15648 800 15678
rect 1577 15675 1643 15678
rect 48129 15738 48195 15741
rect 49200 15738 50000 15768
rect 48129 15736 50000 15738
rect 48129 15680 48134 15736
rect 48190 15680 50000 15736
rect 48129 15678 50000 15680
rect 48129 15675 48195 15678
rect 49200 15648 50000 15678
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 30966 13908 30972 13972
rect 31036 13970 31042 13972
rect 47853 13970 47919 13973
rect 31036 13968 47919 13970
rect 31036 13912 47858 13968
rect 47914 13912 47919 13968
rect 31036 13910 47919 13912
rect 31036 13908 31042 13910
rect 47853 13907 47919 13910
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 48037 13698 48103 13701
rect 49200 13698 50000 13728
rect 48037 13696 50000 13698
rect 48037 13640 48042 13696
rect 48098 13640 50000 13696
rect 48037 13638 50000 13640
rect 48037 13635 48103 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 49200 13608 50000 13638
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 0 11658 800 11688
rect 1485 11658 1551 11661
rect 0 11656 1551 11658
rect 0 11600 1490 11656
rect 1546 11600 1551 11656
rect 0 11598 1551 11600
rect 0 11568 800 11598
rect 1485 11595 1551 11598
rect 48129 11658 48195 11661
rect 49200 11658 50000 11688
rect 48129 11656 50000 11658
rect 48129 11600 48134 11656
rect 48190 11600 50000 11656
rect 48129 11598 50000 11600
rect 48129 11595 48195 11598
rect 49200 11568 50000 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 0 9618 800 9648
rect 1577 9618 1643 9621
rect 0 9616 1643 9618
rect 0 9560 1582 9616
rect 1638 9560 1643 9616
rect 0 9558 1643 9560
rect 0 9528 800 9558
rect 1577 9555 1643 9558
rect 48037 9618 48103 9621
rect 49200 9618 50000 9648
rect 48037 9616 50000 9618
rect 48037 9560 48042 9616
rect 48098 9560 50000 9616
rect 48037 9558 50000 9560
rect 48037 9555 48103 9558
rect 49200 9528 50000 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 0 7578 800 7608
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 1485 7578 1551 7581
rect 0 7576 1551 7578
rect 0 7520 1490 7576
rect 1546 7520 1551 7576
rect 0 7518 1551 7520
rect 0 7488 800 7518
rect 1485 7515 1551 7518
rect 48037 7578 48103 7581
rect 49200 7578 50000 7608
rect 48037 7576 50000 7578
rect 48037 7520 48042 7576
rect 48098 7520 50000 7576
rect 48037 7518 50000 7520
rect 48037 7515 48103 7518
rect 49200 7488 50000 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 0 5538 800 5568
rect 1577 5538 1643 5541
rect 0 5536 1643 5538
rect 0 5480 1582 5536
rect 1638 5480 1643 5536
rect 0 5478 1643 5480
rect 0 5448 800 5478
rect 1577 5475 1643 5478
rect 48037 5538 48103 5541
rect 49200 5538 50000 5568
rect 48037 5536 50000 5538
rect 48037 5480 48042 5536
rect 48098 5480 50000 5536
rect 48037 5478 50000 5480
rect 48037 5475 48103 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 49200 5448 50000 5478
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 28758 3572 28764 3636
rect 28828 3634 28834 3636
rect 47301 3634 47367 3637
rect 28828 3632 47367 3634
rect 28828 3576 47306 3632
rect 47362 3576 47367 3632
rect 28828 3574 47367 3576
rect 28828 3572 28834 3574
rect 47301 3571 47367 3574
rect 0 3498 800 3528
rect 1485 3498 1551 3501
rect 0 3496 1551 3498
rect 0 3440 1490 3496
rect 1546 3440 1551 3496
rect 0 3438 1551 3440
rect 0 3408 800 3438
rect 1485 3435 1551 3438
rect 48037 3498 48103 3501
rect 49200 3498 50000 3528
rect 48037 3496 50000 3498
rect 48037 3440 48042 3496
rect 48098 3440 50000 3496
rect 48037 3438 50000 3440
rect 48037 3435 48103 3438
rect 49200 3408 50000 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 11973 2954 12039 2957
rect 26734 2954 26740 2956
rect 11973 2952 26740 2954
rect 11973 2896 11978 2952
rect 12034 2896 26740 2952
rect 11973 2894 26740 2896
rect 11973 2891 12039 2894
rect 26734 2892 26740 2894
rect 26804 2892 26810 2956
rect 35382 2892 35388 2956
rect 35452 2954 35458 2956
rect 46565 2954 46631 2957
rect 35452 2952 46631 2954
rect 35452 2896 46570 2952
rect 46626 2896 46631 2952
rect 35452 2894 46631 2896
rect 35452 2892 35458 2894
rect 46565 2891 46631 2894
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 14958 2484 14964 2548
rect 15028 2546 15034 2548
rect 15193 2546 15259 2549
rect 15028 2544 15259 2546
rect 15028 2488 15198 2544
rect 15254 2488 15259 2544
rect 15028 2486 15259 2488
rect 15028 2484 15034 2486
rect 15193 2483 15259 2486
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 0 1458 800 1488
rect 1393 1458 1459 1461
rect 0 1456 1459 1458
rect 0 1400 1398 1456
rect 1454 1400 1459 1456
rect 0 1398 1459 1400
rect 0 1368 800 1398
rect 1393 1395 1459 1398
rect 46841 1458 46907 1461
rect 49200 1458 50000 1488
rect 46841 1456 50000 1458
rect 46841 1400 46846 1456
rect 46902 1400 50000 1456
rect 46841 1398 50000 1400
rect 46841 1395 46907 1398
rect 49200 1368 50000 1398
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 30972 46956 31036 47020
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 34652 45928 34716 45932
rect 34652 45872 34702 45928
rect 34702 45872 34716 45928
rect 34652 45868 34716 45872
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 25268 45656 25332 45660
rect 25268 45600 25282 45656
rect 25282 45600 25332 45656
rect 25268 45596 25332 45600
rect 30052 45596 30116 45660
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 26740 41788 26804 41852
rect 28764 41652 28828 41716
rect 30420 41712 30484 41716
rect 30420 41656 30434 41712
rect 30434 41656 30484 41712
rect 30420 41652 30484 41656
rect 28396 41516 28460 41580
rect 35388 41652 35452 41716
rect 19380 41440 19444 41444
rect 19380 41384 19430 41440
rect 19430 41384 19444 41440
rect 19380 41380 19444 41384
rect 33364 41516 33428 41580
rect 32444 41440 32508 41444
rect 32444 41384 32494 41440
rect 32494 41384 32508 41440
rect 32444 41380 32508 41384
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 14964 40488 15028 40492
rect 14964 40432 15014 40488
rect 15014 40432 15028 40488
rect 14964 40428 15028 40432
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 19380 40216 19444 40220
rect 19380 40160 19394 40216
rect 19394 40160 19444 40216
rect 19380 40156 19444 40160
rect 33180 40020 33244 40084
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 26740 39068 26804 39132
rect 35388 38720 35452 38724
rect 35388 38664 35438 38720
rect 35438 38664 35452 38720
rect 35388 38660 35452 38664
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 28396 37768 28460 37772
rect 28396 37712 28446 37768
rect 28446 37712 28460 37768
rect 28396 37708 28460 37712
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 28396 37164 28460 37228
rect 30236 37164 30300 37228
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 32444 36620 32508 36684
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 20484 36000 20548 36004
rect 20484 35944 20498 36000
rect 20498 35944 20548 36000
rect 20484 35940 20548 35944
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 25268 35804 25332 35868
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 30420 34716 30484 34780
rect 33364 34776 33428 34780
rect 33364 34720 33414 34776
rect 33414 34720 33428 34776
rect 33364 34716 33428 34720
rect 30052 34580 30116 34644
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 33180 34172 33244 34236
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19012 31724 19076 31788
rect 19012 31588 19076 31652
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 34652 29548 34716 29612
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 30236 28052 30300 28116
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 20484 27100 20548 27164
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 30972 13908 31036 13972
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 28764 3572 28828 3636
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 26740 2892 26804 2956
rect 35388 2892 35452 2956
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 14964 2484 15028 2548
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 19568 46816 19888 47376
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 30971 47020 31037 47021
rect 30971 46956 30972 47020
rect 31036 46956 31037 47020
rect 30971 46955 31037 46956
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 25267 45660 25333 45661
rect 25267 45596 25268 45660
rect 25332 45596 25333 45660
rect 25267 45595 25333 45596
rect 30051 45660 30117 45661
rect 30051 45596 30052 45660
rect 30116 45596 30117 45660
rect 30051 45595 30117 45596
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19379 41444 19445 41445
rect 19379 41380 19380 41444
rect 19444 41380 19445 41444
rect 19379 41379 19445 41380
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 14963 40492 15029 40493
rect 14963 40428 14964 40492
rect 15028 40428 15029 40492
rect 14963 40427 15029 40428
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 14966 2549 15026 40427
rect 19382 40221 19442 41379
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19379 40220 19445 40221
rect 19379 40156 19380 40220
rect 19444 40156 19445 40220
rect 19379 40155 19445 40156
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 20483 36004 20549 36005
rect 20483 35940 20484 36004
rect 20548 35940 20549 36004
rect 20483 35939 20549 35940
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19011 31788 19077 31789
rect 19011 31724 19012 31788
rect 19076 31724 19077 31788
rect 19011 31723 19077 31724
rect 19014 31653 19074 31723
rect 19011 31652 19077 31653
rect 19011 31588 19012 31652
rect 19076 31588 19077 31652
rect 19011 31587 19077 31588
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 20486 27165 20546 35939
rect 25270 35869 25330 45595
rect 26739 41852 26805 41853
rect 26739 41788 26740 41852
rect 26804 41788 26805 41852
rect 26739 41787 26805 41788
rect 26742 39133 26802 41787
rect 28763 41716 28829 41717
rect 28763 41652 28764 41716
rect 28828 41652 28829 41716
rect 28763 41651 28829 41652
rect 28395 41580 28461 41581
rect 28395 41516 28396 41580
rect 28460 41516 28461 41580
rect 28395 41515 28461 41516
rect 26739 39132 26805 39133
rect 26739 39068 26740 39132
rect 26804 39068 26805 39132
rect 26739 39067 26805 39068
rect 25267 35868 25333 35869
rect 25267 35804 25268 35868
rect 25332 35804 25333 35868
rect 25267 35803 25333 35804
rect 20483 27164 20549 27165
rect 20483 27100 20484 27164
rect 20548 27100 20549 27164
rect 20483 27099 20549 27100
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 14963 2548 15029 2549
rect 14963 2484 14964 2548
rect 15028 2484 15029 2548
rect 14963 2483 15029 2484
rect 19568 2208 19888 3232
rect 26742 2957 26802 39067
rect 28398 37773 28458 41515
rect 28395 37772 28461 37773
rect 28395 37708 28396 37772
rect 28460 37708 28461 37772
rect 28395 37707 28461 37708
rect 28398 37229 28458 37707
rect 28395 37228 28461 37229
rect 28395 37164 28396 37228
rect 28460 37164 28461 37228
rect 28395 37163 28461 37164
rect 28766 3637 28826 41651
rect 30054 34645 30114 45595
rect 30419 41716 30485 41717
rect 30419 41652 30420 41716
rect 30484 41652 30485 41716
rect 30419 41651 30485 41652
rect 30235 37228 30301 37229
rect 30235 37164 30236 37228
rect 30300 37164 30301 37228
rect 30235 37163 30301 37164
rect 30051 34644 30117 34645
rect 30051 34580 30052 34644
rect 30116 34580 30117 34644
rect 30051 34579 30117 34580
rect 30238 28117 30298 37163
rect 30422 34781 30482 41651
rect 30419 34780 30485 34781
rect 30419 34716 30420 34780
rect 30484 34716 30485 34780
rect 30419 34715 30485 34716
rect 30235 28116 30301 28117
rect 30235 28052 30236 28116
rect 30300 28052 30301 28116
rect 30235 28051 30301 28052
rect 30974 13973 31034 46955
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34651 45932 34717 45933
rect 34651 45868 34652 45932
rect 34716 45868 34717 45932
rect 34651 45867 34717 45868
rect 33363 41580 33429 41581
rect 33363 41516 33364 41580
rect 33428 41516 33429 41580
rect 33363 41515 33429 41516
rect 32443 41444 32509 41445
rect 32443 41380 32444 41444
rect 32508 41380 32509 41444
rect 32443 41379 32509 41380
rect 32446 36685 32506 41379
rect 33179 40084 33245 40085
rect 33179 40020 33180 40084
rect 33244 40020 33245 40084
rect 33179 40019 33245 40020
rect 32443 36684 32509 36685
rect 32443 36620 32444 36684
rect 32508 36620 32509 36684
rect 32443 36619 32509 36620
rect 33182 34237 33242 40019
rect 33366 34781 33426 41515
rect 33363 34780 33429 34781
rect 33363 34716 33364 34780
rect 33428 34716 33429 34780
rect 33363 34715 33429 34716
rect 33179 34236 33245 34237
rect 33179 34172 33180 34236
rect 33244 34172 33245 34236
rect 33179 34171 33245 34172
rect 34654 29613 34714 45867
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 35387 41716 35453 41717
rect 35387 41652 35388 41716
rect 35452 41652 35453 41716
rect 35387 41651 35453 41652
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 35390 38725 35450 41651
rect 35387 38724 35453 38725
rect 35387 38660 35388 38724
rect 35452 38660 35453 38724
rect 35387 38659 35453 38660
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34651 29612 34717 29613
rect 34651 29548 34652 29612
rect 34716 29548 34717 29612
rect 34651 29547 34717 29548
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 30971 13972 31037 13973
rect 30971 13908 30972 13972
rect 31036 13908 31037 13972
rect 30971 13907 31037 13908
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 28763 3636 28829 3637
rect 28763 3572 28764 3636
rect 28828 3572 28829 3636
rect 28763 3571 28829 3572
rect 26739 2956 26805 2957
rect 26739 2892 26740 2956
rect 26804 2892 26805 2956
rect 26739 2891 26805 2892
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2752 35248 3776
rect 35390 2957 35450 38659
rect 35387 2956 35453 2957
rect 35387 2892 35388 2956
rect 35452 2892 35453 2956
rect 35387 2891 35453 2892
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__A dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10212 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__B
timestamp 1649977179
transform -1 0 9936 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__A
timestamp 1649977179
transform 1 0 10304 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__B
timestamp 1649977179
transform -1 0 9660 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A
timestamp 1649977179
transform -1 0 11960 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__A
timestamp 1649977179
transform 1 0 10856 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__B
timestamp 1649977179
transform 1 0 11224 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__A1
timestamp 1649977179
transform -1 0 10764 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__A2
timestamp 1649977179
transform 1 0 10304 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__A
timestamp 1649977179
transform -1 0 10488 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__B
timestamp 1649977179
transform 1 0 9660 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A
timestamp 1649977179
transform 1 0 9752 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__B
timestamp 1649977179
transform 1 0 9200 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__A
timestamp 1649977179
transform 1 0 39744 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__B
timestamp 1649977179
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__A
timestamp 1649977179
transform 1 0 11776 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A
timestamp 1649977179
transform 1 0 10856 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__B
timestamp 1649977179
transform 1 0 11132 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A
timestamp 1649977179
transform 1 0 10764 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__B
timestamp 1649977179
transform 1 0 10212 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__B
timestamp 1649977179
transform -1 0 11316 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A
timestamp 1649977179
transform 1 0 40756 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__A
timestamp 1649977179
transform -1 0 48208 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__A
timestamp 1649977179
transform 1 0 35604 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__B1
timestamp 1649977179
transform -1 0 12052 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A
timestamp 1649977179
transform -1 0 42596 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__A
timestamp 1649977179
transform 1 0 41308 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__B
timestamp 1649977179
transform 1 0 12880 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__C1
timestamp 1649977179
transform -1 0 12512 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__A2
timestamp 1649977179
transform -1 0 11868 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__B
timestamp 1649977179
transform -1 0 9752 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__B
timestamp 1649977179
transform 1 0 10120 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A
timestamp 1649977179
transform 1 0 9752 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A
timestamp 1649977179
transform 1 0 40848 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__A
timestamp 1649977179
transform -1 0 38732 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__B
timestamp 1649977179
transform 1 0 11684 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__B
timestamp 1649977179
transform 1 0 10856 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__B
timestamp 1649977179
transform 1 0 12052 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__A
timestamp 1649977179
transform 1 0 41676 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__A1
timestamp 1649977179
transform 1 0 12604 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__B2
timestamp 1649977179
transform -1 0 12604 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__C1
timestamp 1649977179
transform -1 0 12512 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__A1
timestamp 1649977179
transform 1 0 11868 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__A
timestamp 1649977179
transform -1 0 20424 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__A
timestamp 1649977179
transform 1 0 30360 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__A2
timestamp 1649977179
transform 1 0 10580 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__B1
timestamp 1649977179
transform -1 0 11040 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__C1
timestamp 1649977179
transform -1 0 10212 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__A
timestamp 1649977179
transform -1 0 11408 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__A
timestamp 1649977179
transform -1 0 10856 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__A
timestamp 1649977179
transform -1 0 9384 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__A
timestamp 1649977179
transform -1 0 11960 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__B
timestamp 1649977179
transform 1 0 12420 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__A
timestamp 1649977179
transform 1 0 14720 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__B
timestamp 1649977179
transform 1 0 14076 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A2
timestamp 1649977179
transform 1 0 14260 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__B1
timestamp 1649977179
transform 1 0 13984 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__B
timestamp 1649977179
transform 1 0 13432 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__C
timestamp 1649977179
transform 1 0 15456 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A1
timestamp 1649977179
transform 1 0 14536 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__B2
timestamp 1649977179
transform 1 0 13432 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__C1
timestamp 1649977179
transform 1 0 12972 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A1
timestamp 1649977179
transform -1 0 11960 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__A
timestamp 1649977179
transform -1 0 12880 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__B
timestamp 1649977179
transform 1 0 11776 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A
timestamp 1649977179
transform -1 0 12604 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__B
timestamp 1649977179
transform 1 0 12880 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A
timestamp 1649977179
transform -1 0 20516 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__A
timestamp 1649977179
transform 1 0 23736 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__B1
timestamp 1649977179
transform 1 0 17480 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A
timestamp 1649977179
transform 1 0 17480 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__B
timestamp 1649977179
transform 1 0 18584 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__A
timestamp 1649977179
transform 1 0 14352 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__B
timestamp 1649977179
transform 1 0 15732 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__A
timestamp 1649977179
transform 1 0 47104 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__A
timestamp 1649977179
transform 1 0 42136 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__B
timestamp 1649977179
transform 1 0 13524 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__C
timestamp 1649977179
transform 1 0 13708 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__D
timestamp 1649977179
transform 1 0 12880 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A
timestamp 1649977179
transform 1 0 14168 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__A1
timestamp 1649977179
transform 1 0 14812 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A1
timestamp 1649977179
transform 1 0 14628 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A
timestamp 1649977179
transform 1 0 31464 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__B1
timestamp 1649977179
transform -1 0 29716 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A
timestamp 1649977179
transform 1 0 12328 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__A
timestamp 1649977179
transform 1 0 23184 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A
timestamp 1649977179
transform -1 0 23368 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__A
timestamp 1649977179
transform 1 0 14444 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__B
timestamp 1649977179
transform -1 0 16560 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__A
timestamp 1649977179
transform 1 0 17296 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__B
timestamp 1649977179
transform 1 0 18584 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__A
timestamp 1649977179
transform 1 0 21252 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__A1
timestamp 1649977179
transform 1 0 25392 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__B2
timestamp 1649977179
transform -1 0 26128 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__C1
timestamp 1649977179
transform 1 0 21160 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__A1
timestamp 1649977179
transform 1 0 26128 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A
timestamp 1649977179
transform -1 0 15916 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__B
timestamp 1649977179
transform -1 0 16100 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__B2
timestamp 1649977179
transform 1 0 13432 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A
timestamp 1649977179
transform 1 0 34040 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__A
timestamp 1649977179
transform -1 0 35420 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A
timestamp 1649977179
transform 1 0 33672 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__A
timestamp 1649977179
transform 1 0 13432 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A
timestamp 1649977179
transform 1 0 20332 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__B
timestamp 1649977179
transform 1 0 19964 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A
timestamp 1649977179
transform 1 0 16928 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__B
timestamp 1649977179
transform 1 0 18032 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__A1
timestamp 1649977179
transform 1 0 27508 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__B1
timestamp 1649977179
transform 1 0 26772 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A
timestamp 1649977179
transform 1 0 26128 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__B
timestamp 1649977179
transform 1 0 26956 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__A
timestamp 1649977179
transform 1 0 26680 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A1
timestamp 1649977179
transform -1 0 25760 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__B1
timestamp 1649977179
transform -1 0 30360 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__A1
timestamp 1649977179
transform 1 0 12236 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__B1
timestamp 1649977179
transform -1 0 13616 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__B2
timestamp 1649977179
transform -1 0 17112 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A1
timestamp 1649977179
transform 1 0 16008 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A2
timestamp 1649977179
transform 1 0 17480 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__A
timestamp 1649977179
transform -1 0 38364 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__B
timestamp 1649977179
transform -1 0 41676 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A
timestamp 1649977179
transform 1 0 40848 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__B
timestamp 1649977179
transform 1 0 40020 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__A
timestamp 1649977179
transform 1 0 42412 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__A
timestamp 1649977179
transform 1 0 39652 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__A
timestamp 1649977179
transform 1 0 36064 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__B1
timestamp 1649977179
transform 1 0 36616 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__A
timestamp 1649977179
transform 1 0 38364 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__B
timestamp 1649977179
transform 1 0 38916 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__A
timestamp 1649977179
transform 1 0 37260 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__B
timestamp 1649977179
transform 1 0 37812 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__A
timestamp 1649977179
transform 1 0 15088 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__B
timestamp 1649977179
transform 1 0 17848 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__A
timestamp 1649977179
transform 1 0 39100 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A
timestamp 1649977179
transform 1 0 39928 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__A1
timestamp 1649977179
transform 1 0 38732 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__B2
timestamp 1649977179
transform -1 0 35696 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__C1
timestamp 1649977179
transform -1 0 36248 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__A
timestamp 1649977179
transform 1 0 39836 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__B
timestamp 1649977179
transform -1 0 40756 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__A
timestamp 1649977179
transform 1 0 41952 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__B
timestamp 1649977179
transform -1 0 38916 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A1
timestamp 1649977179
transform 1 0 41952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A
timestamp 1649977179
transform 1 0 42964 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__A
timestamp 1649977179
transform 1 0 42964 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__A
timestamp 1649977179
transform 1 0 40756 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__A
timestamp 1649977179
transform 1 0 39836 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__A
timestamp 1649977179
transform -1 0 39192 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__B
timestamp 1649977179
transform 1 0 40204 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A
timestamp 1649977179
transform -1 0 40296 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__B
timestamp 1649977179
transform 1 0 39560 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__B2
timestamp 1649977179
transform -1 0 40020 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__A1
timestamp 1649977179
transform -1 0 40848 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A
timestamp 1649977179
transform 1 0 40480 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__A
timestamp 1649977179
transform 1 0 41584 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__B
timestamp 1649977179
transform 1 0 41032 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A
timestamp 1649977179
transform 1 0 42412 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__B
timestamp 1649977179
transform 1 0 41492 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__A
timestamp 1649977179
transform 1 0 40940 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__B
timestamp 1649977179
transform 1 0 39836 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A1
timestamp 1649977179
transform 1 0 40388 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A2
timestamp 1649977179
transform 1 0 40756 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A
timestamp 1649977179
transform -1 0 32200 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__B
timestamp 1649977179
transform 1 0 39100 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A1
timestamp 1649977179
transform 1 0 40388 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__B1
timestamp 1649977179
transform -1 0 39836 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__B1
timestamp 1649977179
transform -1 0 40388 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__A1
timestamp 1649977179
transform -1 0 42596 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__A2
timestamp 1649977179
transform 1 0 41400 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__B1
timestamp 1649977179
transform 1 0 40388 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__B2
timestamp 1649977179
transform 1 0 39284 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__A1
timestamp 1649977179
transform -1 0 43148 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0944__A
timestamp 1649977179
transform -1 0 43240 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__A
timestamp 1649977179
transform 1 0 41124 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__B
timestamp 1649977179
transform 1 0 39836 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__B1
timestamp 1649977179
transform -1 0 43700 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A
timestamp 1649977179
transform 1 0 42504 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__A1
timestamp 1649977179
transform -1 0 33304 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__D1
timestamp 1649977179
transform 1 0 40388 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__A
timestamp 1649977179
transform -1 0 37444 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A
timestamp 1649977179
transform 1 0 43056 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__B
timestamp 1649977179
transform -1 0 42688 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A1
timestamp 1649977179
transform 1 0 42964 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__A
timestamp 1649977179
transform 1 0 43148 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A
timestamp 1649977179
transform 1 0 42964 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__B1
timestamp 1649977179
transform -1 0 41768 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__B1
timestamp 1649977179
transform 1 0 40940 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A1
timestamp 1649977179
transform -1 0 41216 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__B2
timestamp 1649977179
transform 1 0 33948 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__A
timestamp 1649977179
transform -1 0 37444 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__B
timestamp 1649977179
transform -1 0 36708 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A
timestamp 1649977179
transform 1 0 37076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__B
timestamp 1649977179
transform -1 0 37812 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A1
timestamp 1649977179
transform 1 0 43516 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A2
timestamp 1649977179
transform -1 0 42688 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__B1
timestamp 1649977179
transform 1 0 41676 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A1
timestamp 1649977179
transform 1 0 40940 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A2
timestamp 1649977179
transform -1 0 40572 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A1
timestamp 1649977179
transform -1 0 38916 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A
timestamp 1649977179
transform -1 0 43148 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A
timestamp 1649977179
transform 1 0 43240 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A
timestamp 1649977179
transform 1 0 42044 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__B
timestamp 1649977179
transform 1 0 41216 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A
timestamp 1649977179
transform 1 0 42412 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__B
timestamp 1649977179
transform 1 0 42688 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A
timestamp 1649977179
transform -1 0 42228 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__B
timestamp 1649977179
transform 1 0 43240 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__A1
timestamp 1649977179
transform -1 0 41492 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__B1
timestamp 1649977179
transform 1 0 41492 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__B
timestamp 1649977179
transform 1 0 41584 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A1
timestamp 1649977179
transform 1 0 40480 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__C1
timestamp 1649977179
transform -1 0 40020 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__A
timestamp 1649977179
transform -1 0 23368 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__A
timestamp 1649977179
transform -1 0 34684 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__B
timestamp 1649977179
transform 1 0 33948 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__A
timestamp 1649977179
transform -1 0 35236 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__B
timestamp 1649977179
transform -1 0 36432 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A
timestamp 1649977179
transform 1 0 39468 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A
timestamp 1649977179
transform 1 0 38732 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__B1
timestamp 1649977179
transform 1 0 41400 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__A
timestamp 1649977179
transform 1 0 41860 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__A1
timestamp 1649977179
transform 1 0 41952 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__A
timestamp 1649977179
transform 1 0 43516 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__B
timestamp 1649977179
transform 1 0 42596 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__A
timestamp 1649977179
transform 1 0 43792 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__B
timestamp 1649977179
transform 1 0 42688 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__B2
timestamp 1649977179
transform -1 0 41124 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__A
timestamp 1649977179
transform 1 0 34592 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__B
timestamp 1649977179
transform -1 0 33764 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A
timestamp 1649977179
transform 1 0 38180 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__A
timestamp 1649977179
transform -1 0 31556 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__B
timestamp 1649977179
transform 1 0 37076 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A
timestamp 1649977179
transform -1 0 31004 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__B
timestamp 1649977179
transform 1 0 31096 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__A
timestamp 1649977179
transform -1 0 43148 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__B
timestamp 1649977179
transform 1 0 42412 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__A1
timestamp 1649977179
transform 1 0 42136 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__A2
timestamp 1649977179
transform 1 0 41768 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__A
timestamp 1649977179
transform 1 0 42412 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__B
timestamp 1649977179
transform 1 0 34040 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__A
timestamp 1649977179
transform 1 0 42412 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__A1
timestamp 1649977179
transform -1 0 40572 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__B2
timestamp 1649977179
transform 1 0 34684 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__C1
timestamp 1649977179
transform -1 0 41308 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A1
timestamp 1649977179
transform 1 0 39836 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__A
timestamp 1649977179
transform -1 0 26496 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A
timestamp 1649977179
transform 1 0 30452 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__B
timestamp 1649977179
transform 1 0 31924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A
timestamp 1649977179
transform 1 0 31464 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__B
timestamp 1649977179
transform -1 0 29808 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A
timestamp 1649977179
transform 1 0 32660 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__B
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__A1
timestamp 1649977179
transform 1 0 38088 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__C1
timestamp 1649977179
transform 1 0 38640 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__A1
timestamp 1649977179
transform 1 0 38916 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A1
timestamp 1649977179
transform 1 0 28060 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__A1
timestamp 1649977179
transform 1 0 39192 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__A
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__B
timestamp 1649977179
transform -1 0 33672 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__A
timestamp 1649977179
transform 1 0 10856 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__B
timestamp 1649977179
transform 1 0 11224 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__A
timestamp 1649977179
transform 1 0 11776 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__B
timestamp 1649977179
transform -1 0 12144 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__A1
timestamp 1649977179
transform -1 0 13800 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__A2
timestamp 1649977179
transform 1 0 14352 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A
timestamp 1649977179
transform -1 0 15364 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__B
timestamp 1649977179
transform -1 0 11960 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A
timestamp 1649977179
transform -1 0 36156 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A
timestamp 1649977179
transform 1 0 34684 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__A
timestamp 1649977179
transform 1 0 28336 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__A
timestamp 1649977179
transform 1 0 12236 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__B
timestamp 1649977179
transform 1 0 12788 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__A
timestamp 1649977179
transform -1 0 12420 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__B
timestamp 1649977179
transform 1 0 11684 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__A1
timestamp 1649977179
transform -1 0 37444 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__B1
timestamp 1649977179
transform -1 0 39376 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__C1
timestamp 1649977179
transform 1 0 37812 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__A1
timestamp 1649977179
transform -1 0 31464 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__A2
timestamp 1649977179
transform -1 0 37444 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__B2
timestamp 1649977179
transform 1 0 28244 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__C1
timestamp 1649977179
transform 1 0 30820 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A
timestamp 1649977179
transform 1 0 12236 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__B
timestamp 1649977179
transform 1 0 12880 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__A
timestamp 1649977179
transform -1 0 12512 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__B
timestamp 1649977179
transform 1 0 11408 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__B1
timestamp 1649977179
transform 1 0 13340 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__A
timestamp 1649977179
transform 1 0 10672 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__B
timestamp 1649977179
transform -1 0 13248 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__A
timestamp 1649977179
transform -1 0 10488 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__B
timestamp 1649977179
transform -1 0 11132 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__A
timestamp 1649977179
transform -1 0 11408 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__B1
timestamp 1649977179
transform 1 0 11776 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__A
timestamp 1649977179
transform 1 0 13432 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__B
timestamp 1649977179
transform 1 0 31372 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__C
timestamp 1649977179
transform 1 0 35052 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__A2
timestamp 1649977179
transform 1 0 30360 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__B1
timestamp 1649977179
transform 1 0 27692 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__B
timestamp 1649977179
transform 1 0 30728 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__B1
timestamp 1649977179
transform 1 0 26312 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__A1
timestamp 1649977179
transform -1 0 26220 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__B1
timestamp 1649977179
transform 1 0 26128 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__A1
timestamp 1649977179
transform -1 0 25668 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__A
timestamp 1649977179
transform 1 0 11224 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__B
timestamp 1649977179
transform 1 0 10856 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__A
timestamp 1649977179
transform 1 0 11132 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__B
timestamp 1649977179
transform 1 0 11684 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__A1
timestamp 1649977179
transform 1 0 11960 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__A2
timestamp 1649977179
transform 1 0 12788 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__A
timestamp 1649977179
transform 1 0 10396 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__B
timestamp 1649977179
transform 1 0 10856 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__A
timestamp 1649977179
transform 1 0 10304 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__B
timestamp 1649977179
transform 1 0 9752 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__A1
timestamp 1649977179
transform -1 0 12696 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__A2
timestamp 1649977179
transform 1 0 10120 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__A
timestamp 1649977179
transform 1 0 10304 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__A
timestamp 1649977179
transform 1 0 10856 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__A1
timestamp 1649977179
transform 1 0 12788 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__B2
timestamp 1649977179
transform 1 0 13156 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__A
timestamp 1649977179
transform -1 0 11040 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__B
timestamp 1649977179
transform 1 0 11776 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__A
timestamp 1649977179
transform 1 0 10304 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__B
timestamp 1649977179
transform 1 0 10856 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__A
timestamp 1649977179
transform 1 0 20516 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__A
timestamp 1649977179
transform 1 0 23736 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__B
timestamp 1649977179
transform 1 0 23828 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__A1
timestamp 1649977179
transform 1 0 26956 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__B1
timestamp 1649977179
transform 1 0 26128 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__A
timestamp 1649977179
transform 1 0 9660 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__B
timestamp 1649977179
transform 1 0 10304 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__A
timestamp 1649977179
transform 1 0 9752 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__B
timestamp 1649977179
transform -1 0 9292 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__B1
timestamp 1649977179
transform 1 0 10672 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__A
timestamp 1649977179
transform -1 0 10304 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__A1
timestamp 1649977179
transform -1 0 10396 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__A1
timestamp 1649977179
transform 1 0 24932 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__B2
timestamp 1649977179
transform 1 0 21344 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__A1
timestamp 1649977179
transform 1 0 14904 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__A2
timestamp 1649977179
transform 1 0 14168 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__A
timestamp 1649977179
transform 1 0 16468 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__B
timestamp 1649977179
transform 1 0 15364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__A
timestamp 1649977179
transform 1 0 15732 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__B
timestamp 1649977179
transform 1 0 14812 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__A
timestamp 1649977179
transform 1 0 10856 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__A
timestamp 1649977179
transform 1 0 23736 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__A
timestamp 1649977179
transform 1 0 19228 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__B
timestamp 1649977179
transform 1 0 23276 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__C
timestamp 1649977179
transform 1 0 19780 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__A
timestamp 1649977179
transform 1 0 11776 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__B
timestamp 1649977179
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__A
timestamp 1649977179
transform -1 0 11960 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__B
timestamp 1649977179
transform 1 0 11224 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__A
timestamp 1649977179
transform -1 0 11868 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__B
timestamp 1649977179
transform 1 0 10856 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__B2
timestamp 1649977179
transform 1 0 19780 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__C1
timestamp 1649977179
transform 1 0 22908 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__A1
timestamp 1649977179
transform 1 0 19228 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__A1
timestamp 1649977179
transform 1 0 23000 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__A
timestamp 1649977179
transform -1 0 11408 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__B
timestamp 1649977179
transform -1 0 12236 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__A
timestamp 1649977179
transform 1 0 13708 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__B
timestamp 1649977179
transform 1 0 14904 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__A
timestamp 1649977179
transform 1 0 14260 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__B
timestamp 1649977179
transform -1 0 17020 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__A
timestamp 1649977179
transform 1 0 17388 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__B
timestamp 1649977179
transform 1 0 18676 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__A
timestamp 1649977179
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__B1
timestamp 1649977179
transform 1 0 14812 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__A1
timestamp 1649977179
transform 1 0 11960 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__A
timestamp 1649977179
transform 1 0 14260 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__A1
timestamp 1649977179
transform 1 0 13156 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__B2
timestamp 1649977179
transform 1 0 12604 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__A
timestamp 1649977179
transform -1 0 12512 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__B
timestamp 1649977179
transform 1 0 12880 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__A
timestamp 1649977179
transform 1 0 16928 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__B
timestamp 1649977179
transform 1 0 19412 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__A
timestamp 1649977179
transform -1 0 12512 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__B
timestamp 1649977179
transform 1 0 12880 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__A1
timestamp 1649977179
transform 1 0 17204 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__B1
timestamp 1649977179
transform 1 0 20700 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__A
timestamp 1649977179
transform 1 0 17756 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__B
timestamp 1649977179
transform 1 0 22632 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__A
timestamp 1649977179
transform -1 0 17848 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__B
timestamp 1649977179
transform -1 0 14904 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__A
timestamp 1649977179
transform 1 0 17020 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__B
timestamp 1649977179
transform 1 0 17756 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__A
timestamp 1649977179
transform -1 0 18952 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1240__B1
timestamp 1649977179
transform 1 0 18584 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__A1
timestamp 1649977179
transform 1 0 14168 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__A1
timestamp 1649977179
transform 1 0 19964 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__A
timestamp 1649977179
transform 1 0 16008 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__B
timestamp 1649977179
transform 1 0 16836 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__A
timestamp 1649977179
transform -1 0 14536 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__B
timestamp 1649977179
transform 1 0 18400 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__B1
timestamp 1649977179
transform 1 0 16008 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__A
timestamp 1649977179
transform 1 0 18032 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__A1
timestamp 1649977179
transform 1 0 21160 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__A
timestamp 1649977179
transform 1 0 19596 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__B
timestamp 1649977179
transform -1 0 20608 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__A
timestamp 1649977179
transform 1 0 19504 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__B
timestamp 1649977179
transform 1 0 20516 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__A
timestamp 1649977179
transform 1 0 17480 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1262__B1
timestamp 1649977179
transform 1 0 15456 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__B2
timestamp 1649977179
transform 1 0 18584 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__B1
timestamp 1649977179
transform 1 0 17480 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__A
timestamp 1649977179
transform 1 0 22264 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__B
timestamp 1649977179
transform 1 0 22908 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__A
timestamp 1649977179
transform 1 0 19964 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__B
timestamp 1649977179
transform 1 0 21896 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__A
timestamp 1649977179
transform -1 0 18768 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__A
timestamp 1649977179
transform 1 0 16836 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__B
timestamp 1649977179
transform 1 0 22264 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__A
timestamp 1649977179
transform -1 0 20424 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__B
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__A1
timestamp 1649977179
transform 1 0 16008 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__A2
timestamp 1649977179
transform 1 0 16744 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__A
timestamp 1649977179
transform 1 0 19872 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__A1
timestamp 1649977179
transform -1 0 23552 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__B2
timestamp 1649977179
transform 1 0 23736 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__C1
timestamp 1649977179
transform 1 0 23920 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__A1
timestamp 1649977179
transform 1 0 21436 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__A1
timestamp 1649977179
transform 1 0 26128 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__B1
timestamp 1649977179
transform 1 0 25576 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__A
timestamp 1649977179
transform 1 0 25576 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__B
timestamp 1649977179
transform 1 0 25300 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__A1
timestamp 1649977179
transform 1 0 18584 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__B2
timestamp 1649977179
transform 1 0 19872 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__A1
timestamp 1649977179
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__A
timestamp 1649977179
transform -1 0 21988 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__B
timestamp 1649977179
transform 1 0 22448 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__A
timestamp 1649977179
transform 1 0 20792 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__B
timestamp 1649977179
transform 1 0 21344 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__A
timestamp 1649977179
transform 1 0 23092 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__B1
timestamp 1649977179
transform 1 0 23736 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1319__A
timestamp 1649977179
transform 1 0 16560 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1319__B
timestamp 1649977179
transform 1 0 18584 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1320__A
timestamp 1649977179
transform 1 0 18584 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1320__B
timestamp 1649977179
transform 1 0 21988 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__A
timestamp 1649977179
transform 1 0 24472 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__C1
timestamp 1649977179
transform 1 0 25944 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1326__A
timestamp 1649977179
transform 1 0 23552 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1326__B
timestamp 1649977179
transform 1 0 25760 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__A
timestamp 1649977179
transform 1 0 24104 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__B
timestamp 1649977179
transform 1 0 25116 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1331__A
timestamp 1649977179
transform 1 0 23736 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__A
timestamp 1649977179
transform 1 0 23276 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__B
timestamp 1649977179
transform 1 0 22264 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__A
timestamp 1649977179
transform -1 0 21344 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__B
timestamp 1649977179
transform -1 0 21160 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1338__A
timestamp 1649977179
transform 1 0 24288 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1341__A
timestamp 1649977179
transform 1 0 26956 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__A1
timestamp 1649977179
transform -1 0 23920 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1343__A1
timestamp 1649977179
transform 1 0 26404 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__A
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__B
timestamp 1649977179
transform 1 0 25944 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__A
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__B
timestamp 1649977179
transform 1 0 28336 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__A
timestamp 1649977179
transform 1 0 27692 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1353__A
timestamp 1649977179
transform 1 0 26128 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1353__B
timestamp 1649977179
transform 1 0 27048 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__A
timestamp 1649977179
transform 1 0 25392 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__B
timestamp 1649977179
transform -1 0 24564 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1358__A
timestamp 1649977179
transform -1 0 26680 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__B1
timestamp 1649977179
transform 1 0 26312 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1363__A1
timestamp 1649977179
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1364__A1
timestamp 1649977179
transform 1 0 25944 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1368__A1
timestamp 1649977179
transform 1 0 27324 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1369__A1
timestamp 1649977179
transform 1 0 27876 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1371__A
timestamp 1649977179
transform 1 0 25024 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1371__B
timestamp 1649977179
transform 1 0 23736 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1372__A
timestamp 1649977179
transform 1 0 23184 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1372__B
timestamp 1649977179
transform -1 0 23552 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1374__A
timestamp 1649977179
transform -1 0 24656 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1374__B
timestamp 1649977179
transform -1 0 25852 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1377__A
timestamp 1649977179
transform 1 0 27692 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__B1
timestamp 1649977179
transform -1 0 29164 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1386__A
timestamp 1649977179
transform -1 0 26496 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1386__B
timestamp 1649977179
transform 1 0 28152 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1387__A
timestamp 1649977179
transform -1 0 29072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1387__B
timestamp 1649977179
transform 1 0 28888 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__A
timestamp 1649977179
transform 1 0 32660 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__B
timestamp 1649977179
transform -1 0 34960 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1392__A1
timestamp 1649977179
transform 1 0 28244 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1392__A2
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1392__B1
timestamp 1649977179
transform 1 0 32108 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__A1
timestamp 1649977179
transform 1 0 28704 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__A
timestamp 1649977179
transform 1 0 35972 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__B
timestamp 1649977179
transform 1 0 29624 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1398__A
timestamp 1649977179
transform -1 0 31372 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1398__B
timestamp 1649977179
transform 1 0 31372 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__B1
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1403__A
timestamp 1649977179
transform 1 0 28244 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1403__B
timestamp 1649977179
transform -1 0 28796 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__A
timestamp 1649977179
transform 1 0 27600 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__B
timestamp 1649977179
transform 1 0 26956 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1408__A
timestamp 1649977179
transform 1 0 29072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__A1
timestamp 1649977179
transform 1 0 28704 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1410__A1
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__A
timestamp 1649977179
transform 1 0 33580 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1417__A1
timestamp 1649977179
transform -1 0 35604 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1420__A
timestamp 1649977179
transform 1 0 28796 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1422__A
timestamp 1649977179
transform -1 0 31464 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1422__B
timestamp 1649977179
transform -1 0 32016 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1423__A
timestamp 1649977179
transform 1 0 32476 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1423__B
timestamp 1649977179
transform 1 0 33028 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1425__A
timestamp 1649977179
transform 1 0 28704 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1425__B
timestamp 1649977179
transform 1 0 26312 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1428__A
timestamp 1649977179
transform 1 0 34040 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1429__A
timestamp 1649977179
transform 1 0 31924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1431__B1
timestamp 1649977179
transform 1 0 30176 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1433__A
timestamp 1649977179
transform 1 0 36708 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__A
timestamp 1649977179
transform 1 0 36156 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1435__A
timestamp 1649977179
transform -1 0 33212 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1435__B
timestamp 1649977179
transform 1 0 32292 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__A
timestamp 1649977179
transform 1 0 36524 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__B
timestamp 1649977179
transform 1 0 31740 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1440__B1
timestamp 1649977179
transform -1 0 33028 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1441__A1
timestamp 1649977179
transform -1 0 35788 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1442__B1
timestamp 1649977179
transform 1 0 34684 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1443__B
timestamp 1649977179
transform -1 0 33580 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__A
timestamp 1649977179
transform 1 0 36984 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__A
timestamp 1649977179
transform 1 0 28244 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1454__A
timestamp 1649977179
transform 1 0 34040 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1455__C1
timestamp 1649977179
transform 1 0 39192 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1459__A
timestamp 1649977179
transform 1 0 12236 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1460__A2
timestamp 1649977179
transform -1 0 12328 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1460__C1
timestamp 1649977179
transform 1 0 13432 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__A1
timestamp 1649977179
transform 1 0 11868 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__A1
timestamp 1649977179
transform 1 0 10856 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__A2
timestamp 1649977179
transform -1 0 10488 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__B1
timestamp 1649977179
transform 1 0 11684 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1463__A2
timestamp 1649977179
transform -1 0 11500 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1463__C1
timestamp 1649977179
transform -1 0 11776 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1489__D
timestamp 1649977179
transform -1 0 35972 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1649977179
transform -1 0 31096 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 47472 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 47564 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 48208 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 1748 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 43516 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 2668 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 48208 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 35788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 1748 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 1748 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 12604 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 1748 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 4876 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 1748 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 1748 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 48208 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 34224 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 41952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 1748 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 1748 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 1748 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 28428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 19596 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 46920 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 2852 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 48208 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 31648 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 10488 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 46736 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 20700 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 1748 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 48208 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 11040 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 48208 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 48208 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 12512 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 40020 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 48208 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 7452 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 1748 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 24748 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 2300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 29992 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 9752 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 30636 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 1748 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 3220 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 6808 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 3036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 45356 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 35052 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 22264 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 47288 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 47472 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 2668 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 48208 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 9292 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 17020 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 1748 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform -1 0 48208 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1649977179
transform -1 0 26496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1649977179
transform -1 0 40296 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1649977179
transform -1 0 38364 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1649977179
transform -1 0 4784 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1649977179
transform -1 0 9200 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1649977179
transform -1 0 34224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1649977179
transform -1 0 1564 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1649977179
transform -1 0 1564 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1649977179
transform -1 0 48208 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output70_A
timestamp 1649977179
transform -1 0 8832 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output71_A
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output72_A
timestamp 1649977179
transform 1 0 11868 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output73_A
timestamp 1649977179
transform 1 0 47288 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output74_A
timestamp 1649977179
transform 1 0 47564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output75_A
timestamp 1649977179
transform 1 0 47288 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output76_A
timestamp 1649977179
transform -1 0 36800 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output77_A
timestamp 1649977179
transform -1 0 9384 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output78_A
timestamp 1649977179
transform 1 0 46552 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output79_A
timestamp 1649977179
transform 1 0 47288 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output80_A
timestamp 1649977179
transform 1 0 46184 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output82_A
timestamp 1649977179
transform 1 0 2116 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output83_A
timestamp 1649977179
transform 1 0 47288 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output84_A
timestamp 1649977179
transform 1 0 2116 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output85_A
timestamp 1649977179
transform 1 0 2116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output86_A
timestamp 1649977179
transform -1 0 34224 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output87_A
timestamp 1649977179
transform 1 0 2116 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output88_A
timestamp 1649977179
transform 1 0 37536 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output89_A
timestamp 1649977179
transform 1 0 42412 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output90_A
timestamp 1649977179
transform -1 0 2300 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output91_A
timestamp 1649977179
transform 1 0 4140 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output92_A
timestamp 1649977179
transform 1 0 15640 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output93_A
timestamp 1649977179
transform 1 0 45264 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output94_A
timestamp 1649977179
transform 1 0 47288 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output95_A
timestamp 1649977179
transform -1 0 47840 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output96_A
timestamp 1649977179
transform 1 0 2116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output97_A
timestamp 1649977179
transform 1 0 2116 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output98_A
timestamp 1649977179
transform 1 0 47288 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output99_A
timestamp 1649977179
transform 1 0 6716 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output100_A
timestamp 1649977179
transform -1 0 47840 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output101_A
timestamp 1649977179
transform -1 0 47840 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater102_A
timestamp 1649977179
transform 1 0 28796 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater103_A
timestamp 1649977179
transform 1 0 31648 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33
timestamp 1649977179
transform 1 0 4140 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49
timestamp 1649977179
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1649977179
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62
timestamp 1649977179
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7544 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93
timestamp 1649977179
transform 1 0 9660 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105
timestamp 1649977179
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1649977179
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117
timestamp 1649977179
transform 1 0 11868 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_133
timestamp 1649977179
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1649977179
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149
timestamp 1649977179
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_154
timestamp 1649977179
transform 1 0 15272 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_160
timestamp 1649977179
transform 1 0 15824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_177
timestamp 1649977179
transform 1 0 17388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189
timestamp 1649977179
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1649977179
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_205
timestamp 1649977179
transform 1 0 19964 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217
timestamp 1649977179
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1649977179
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1649977179
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_244
timestamp 1649977179
transform 1 0 23552 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_253
timestamp 1649977179
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_261
timestamp 1649977179
transform 1 0 25116 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_273
timestamp 1649977179
transform 1 0 26220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1649977179
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_291
timestamp 1649977179
transform 1 0 27876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1649977179
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1649977179
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_314
timestamp 1649977179
transform 1 0 29992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_328
timestamp 1649977179
transform 1 0 31280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_343
timestamp 1649977179
transform 1 0 32660 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_355
timestamp 1649977179
transform 1 0 33764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1649977179
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_369
timestamp 1649977179
transform 1 0 35052 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 1649977179
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_387
timestamp 1649977179
transform 1 0 36708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1649977179
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_393
timestamp 1649977179
transform 1 0 37260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_398
timestamp 1649977179
transform 1 0 37720 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_406
timestamp 1649977179
transform 1 0 38456 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_418
timestamp 1649977179
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1649977179
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_427
timestamp 1649977179
transform 1 0 40388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_439
timestamp 1649977179
transform 1 0 41492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_444
timestamp 1649977179
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_453
timestamp 1649977179
transform 1 0 42780 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_461
timestamp 1649977179
transform 1 0 43516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_471
timestamp 1649977179
transform 1 0 44436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1649977179
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_477
timestamp 1649977179
transform 1 0 44988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_482
timestamp 1649977179
transform 1 0 45448 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_490
timestamp 1649977179
transform 1 0 46184 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1649977179
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1649977179
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_511
timestamp 1649977179
transform 1 0 48116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_515
timestamp 1649977179
transform 1 0 48484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_7
timestamp 1649977179
transform 1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1649977179
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_19
timestamp 1649977179
transform 1 0 2852 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_31
timestamp 1649977179
transform 1 0 3956 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_35
timestamp 1649977179
transform 1 0 4324 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_47
timestamp 1649977179
transform 1 0 5428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_89
timestamp 1649977179
transform 1 0 9292 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_101
timestamp 1649977179
transform 1 0 10396 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_109
timestamp 1649977179
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_119
timestamp 1649977179
transform 1 0 12052 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_131
timestamp 1649977179
transform 1 0 13156 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_143
timestamp 1649977179
transform 1 0 14260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_155
timestamp 1649977179
transform 1 0 15364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_173
timestamp 1649977179
transform 1 0 17020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_185
timestamp 1649977179
transform 1 0 18124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_197
timestamp 1649977179
transform 1 0 19228 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_201
timestamp 1649977179
transform 1 0 19596 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_209
timestamp 1649977179
transform 1 0 20332 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_213
timestamp 1649977179
transform 1 0 20700 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_221
timestamp 1649977179
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1649977179
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_249
timestamp 1649977179
transform 1 0 24012 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_257
timestamp 1649977179
transform 1 0 24748 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_269
timestamp 1649977179
transform 1 0 25852 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_277
timestamp 1649977179
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_293
timestamp 1649977179
transform 1 0 28060 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_297
timestamp 1649977179
transform 1 0 28428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_309
timestamp 1649977179
transform 1 0 29532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_321
timestamp 1649977179
transform 1 0 30636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_333
timestamp 1649977179
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_339
timestamp 1649977179
transform 1 0 32292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_351
timestamp 1649977179
transform 1 0 33396 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_363
timestamp 1649977179
transform 1 0 34500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_375
timestamp 1649977179
transform 1 0 35604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_387
timestamp 1649977179
transform 1 0 36708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1649977179
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1649977179
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1649977179
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_417
timestamp 1649977179
transform 1 0 39468 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_423
timestamp 1649977179
transform 1 0 40020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_435
timestamp 1649977179
transform 1 0 41124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1649977179
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1649977179
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1649977179
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1649977179
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_485
timestamp 1649977179
transform 1 0 45724 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_493
timestamp 1649977179
transform 1 0 46460 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_496
timestamp 1649977179
transform 1 0 46736 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_505
timestamp 1649977179
transform 1 0 47564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_512
timestamp 1649977179
transform 1 0 48208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_7
timestamp 1649977179
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_13
timestamp 1649977179
transform 1 0 2300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_25
timestamp 1649977179
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1649977179
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1649977179
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1649977179
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1649977179
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1649977179
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1649977179
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1649977179
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1649977179
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1649977179
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1649977179
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1649977179
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1649977179
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1649977179
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1649977179
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1649977179
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1649977179
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1649977179
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1649977179
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1649977179
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1649977179
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1649977179
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1649977179
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1649977179
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1649977179
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1649977179
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_489
timestamp 1649977179
transform 1 0 46092 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_495
timestamp 1649977179
transform 1 0 46644 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_498
timestamp 1649977179
transform 1 0 46920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_504
timestamp 1649977179
transform 1 0 47472 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1649977179
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1649977179
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1649977179
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1649977179
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1649977179
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1649977179
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1649977179
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1649977179
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1649977179
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1649977179
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1649977179
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1649977179
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1649977179
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1649977179
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1649977179
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1649977179
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1649977179
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1649977179
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1649977179
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1649977179
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1649977179
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1649977179
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1649977179
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1649977179
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_507
timestamp 1649977179
transform 1 0 47748 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_515
timestamp 1649977179
transform 1 0 48484 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1649977179
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1649977179
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1649977179
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1649977179
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1649977179
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1649977179
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1649977179
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1649977179
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1649977179
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1649977179
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1649977179
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1649977179
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1649977179
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1649977179
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1649977179
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1649977179
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1649977179
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1649977179
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1649977179
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1649977179
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1649977179
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1649977179
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1649977179
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1649977179
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1649977179
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1649977179
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_513
timestamp 1649977179
transform 1 0 48300 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7
timestamp 1649977179
transform 1 0 1748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_19
timestamp 1649977179
transform 1 0 2852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_31
timestamp 1649977179
transform 1 0 3956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_43
timestamp 1649977179
transform 1 0 5060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1649977179
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1649977179
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1649977179
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1649977179
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1649977179
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1649977179
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1649977179
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1649977179
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1649977179
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1649977179
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1649977179
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1649977179
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1649977179
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1649977179
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1649977179
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1649977179
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1649977179
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1649977179
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1649977179
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1649977179
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1649977179
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1649977179
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1649977179
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1649977179
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_505
timestamp 1649977179
transform 1 0 47564 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_513
timestamp 1649977179
transform 1 0 48300 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_11
timestamp 1649977179
transform 1 0 2116 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1649977179
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1649977179
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1649977179
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1649977179
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1649977179
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1649977179
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1649977179
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1649977179
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1649977179
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1649977179
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1649977179
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1649977179
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1649977179
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1649977179
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1649977179
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1649977179
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1649977179
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1649977179
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1649977179
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1649977179
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1649977179
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1649977179
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1649977179
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_501
timestamp 1649977179
transform 1 0 47196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_504
timestamp 1649977179
transform 1 0 47472 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_512
timestamp 1649977179
transform 1 0 48208 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1649977179
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1649977179
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1649977179
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1649977179
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1649977179
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1649977179
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1649977179
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1649977179
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1649977179
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1649977179
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1649977179
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1649977179
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1649977179
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1649977179
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1649977179
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1649977179
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1649977179
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1649977179
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1649977179
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_505
timestamp 1649977179
transform 1 0 47564 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_513
timestamp 1649977179
transform 1 0 48300 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1649977179
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1649977179
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1649977179
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1649977179
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1649977179
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1649977179
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1649977179
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1649977179
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1649977179
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1649977179
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1649977179
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1649977179
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1649977179
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1649977179
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1649977179
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1649977179
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1649977179
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1649977179
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1649977179
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1649977179
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1649977179
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1649977179
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1649977179
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1649977179
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1649977179
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1649977179
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_513
timestamp 1649977179
transform 1 0 48300 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1649977179
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1649977179
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1649977179
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1649977179
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1649977179
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1649977179
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1649977179
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1649977179
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1649977179
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1649977179
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1649977179
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1649977179
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1649977179
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1649977179
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1649977179
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1649977179
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1649977179
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1649977179
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1649977179
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1649977179
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1649977179
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1649977179
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1649977179
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1649977179
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_505
timestamp 1649977179
transform 1 0 47564 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_513
timestamp 1649977179
transform 1 0 48300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_7
timestamp 1649977179
transform 1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_13
timestamp 1649977179
transform 1 0 2300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1649977179
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1649977179
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1649977179
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1649977179
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1649977179
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1649977179
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1649977179
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1649977179
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1649977179
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1649977179
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1649977179
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1649977179
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1649977179
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1649977179
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1649977179
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1649977179
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1649977179
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1649977179
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1649977179
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1649977179
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1649977179
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1649977179
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1649977179
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1649977179
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1649977179
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1649977179
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1649977179
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_501
timestamp 1649977179
transform 1 0 47196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_504
timestamp 1649977179
transform 1 0 47472 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_512
timestamp 1649977179
transform 1 0 48208 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1649977179
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1649977179
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1649977179
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1649977179
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1649977179
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1649977179
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1649977179
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1649977179
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1649977179
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1649977179
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1649977179
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1649977179
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1649977179
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1649977179
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1649977179
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1649977179
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1649977179
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1649977179
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1649977179
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1649977179
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1649977179
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1649977179
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1649977179
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1649977179
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_505
timestamp 1649977179
transform 1 0 47564 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_513
timestamp 1649977179
transform 1 0 48300 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1649977179
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1649977179
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1649977179
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1649977179
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1649977179
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1649977179
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1649977179
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1649977179
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1649977179
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1649977179
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1649977179
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1649977179
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1649977179
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1649977179
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1649977179
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1649977179
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1649977179
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1649977179
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1649977179
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1649977179
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1649977179
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1649977179
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1649977179
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1649977179
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1649977179
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1649977179
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_513
timestamp 1649977179
transform 1 0 48300 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_7
timestamp 1649977179
transform 1 0 1748 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_19
timestamp 1649977179
transform 1 0 2852 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_31
timestamp 1649977179
transform 1 0 3956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_43
timestamp 1649977179
transform 1 0 5060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1649977179
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1649977179
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1649977179
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1649977179
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1649977179
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1649977179
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1649977179
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1649977179
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1649977179
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1649977179
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1649977179
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1649977179
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1649977179
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1649977179
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1649977179
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1649977179
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1649977179
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1649977179
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1649977179
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1649977179
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1649977179
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1649977179
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1649977179
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_505
timestamp 1649977179
transform 1 0 47564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_513
timestamp 1649977179
transform 1 0 48300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_13
timestamp 1649977179
transform 1 0 2300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 1649977179
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1649977179
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1649977179
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1649977179
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1649977179
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1649977179
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1649977179
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1649977179
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1649977179
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1649977179
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1649977179
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1649977179
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1649977179
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1649977179
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1649977179
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1649977179
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1649977179
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1649977179
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1649977179
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1649977179
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1649977179
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1649977179
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1649977179
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1649977179
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1649977179
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1649977179
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_501
timestamp 1649977179
transform 1 0 47196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_504
timestamp 1649977179
transform 1 0 47472 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_512
timestamp 1649977179
transform 1 0 48208 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1649977179
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1649977179
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1649977179
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1649977179
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1649977179
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1649977179
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1649977179
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1649977179
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1649977179
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1649977179
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1649977179
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1649977179
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1649977179
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1649977179
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1649977179
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1649977179
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1649977179
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1649977179
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1649977179
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1649977179
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1649977179
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1649977179
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1649977179
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1649977179
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1649977179
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1649977179
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_505
timestamp 1649977179
transform 1 0 47564 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_513
timestamp 1649977179
transform 1 0 48300 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1649977179
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1649977179
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1649977179
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1649977179
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1649977179
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1649977179
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1649977179
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1649977179
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1649977179
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1649977179
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1649977179
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1649977179
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1649977179
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1649977179
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1649977179
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1649977179
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1649977179
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1649977179
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1649977179
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1649977179
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1649977179
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1649977179
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1649977179
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1649977179
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1649977179
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1649977179
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_501
timestamp 1649977179
transform 1 0 47196 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_509
timestamp 1649977179
transform 1 0 47932 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_512
timestamp 1649977179
transform 1 0 48208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_7
timestamp 1649977179
transform 1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_13
timestamp 1649977179
transform 1 0 2300 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_25
timestamp 1649977179
transform 1 0 3404 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_37
timestamp 1649977179
transform 1 0 4508 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_49
timestamp 1649977179
transform 1 0 5612 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1649977179
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1649977179
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1649977179
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1649977179
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1649977179
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1649977179
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1649977179
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1649977179
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1649977179
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1649977179
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1649977179
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1649977179
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1649977179
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1649977179
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1649977179
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1649977179
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1649977179
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1649977179
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1649977179
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1649977179
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1649977179
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1649977179
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1649977179
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_505
timestamp 1649977179
transform 1 0 47564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_512
timestamp 1649977179
transform 1 0 48208 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1649977179
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1649977179
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1649977179
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1649977179
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1649977179
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1649977179
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1649977179
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1649977179
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1649977179
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1649977179
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1649977179
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1649977179
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1649977179
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1649977179
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1649977179
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1649977179
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1649977179
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1649977179
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1649977179
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1649977179
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1649977179
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1649977179
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1649977179
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1649977179
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1649977179
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_513
timestamp 1649977179
transform 1 0 48300 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1649977179
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1649977179
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1649977179
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1649977179
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1649977179
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1649977179
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1649977179
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1649977179
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1649977179
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1649977179
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1649977179
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1649977179
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1649977179
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1649977179
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1649977179
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1649977179
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1649977179
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1649977179
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1649977179
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1649977179
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1649977179
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1649977179
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1649977179
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1649977179
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1649977179
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1649977179
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_505
timestamp 1649977179
transform 1 0 47564 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_513
timestamp 1649977179
transform 1 0 48300 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_5
timestamp 1649977179
transform 1 0 1564 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_17
timestamp 1649977179
transform 1 0 2668 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_25
timestamp 1649977179
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1649977179
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1649977179
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1649977179
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1649977179
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1649977179
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1649977179
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1649977179
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1649977179
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1649977179
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1649977179
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1649977179
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1649977179
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1649977179
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1649977179
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1649977179
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1649977179
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1649977179
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1649977179
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1649977179
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1649977179
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1649977179
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1649977179
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1649977179
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1649977179
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1649977179
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1649977179
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_501
timestamp 1649977179
transform 1 0 47196 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_505
timestamp 1649977179
transform 1 0 47564 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_508
timestamp 1649977179
transform 1 0 47840 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_7
timestamp 1649977179
transform 1 0 1748 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_19
timestamp 1649977179
transform 1 0 2852 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_31
timestamp 1649977179
transform 1 0 3956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_43
timestamp 1649977179
transform 1 0 5060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1649977179
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1649977179
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1649977179
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1649977179
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1649977179
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1649977179
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1649977179
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1649977179
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1649977179
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1649977179
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1649977179
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1649977179
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1649977179
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1649977179
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1649977179
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1649977179
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1649977179
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1649977179
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1649977179
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1649977179
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1649977179
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1649977179
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1649977179
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1649977179
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1649977179
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1649977179
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_505
timestamp 1649977179
transform 1 0 47564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_512
timestamp 1649977179
transform 1 0 48208 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1649977179
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1649977179
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1649977179
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1649977179
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1649977179
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1649977179
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1649977179
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1649977179
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1649977179
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1649977179
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1649977179
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1649977179
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1649977179
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1649977179
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1649977179
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1649977179
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1649977179
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1649977179
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1649977179
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1649977179
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1649977179
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1649977179
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1649977179
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1649977179
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1649977179
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1649977179
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_513
timestamp 1649977179
transform 1 0 48300 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1649977179
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1649977179
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1649977179
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1649977179
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1649977179
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1649977179
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1649977179
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1649977179
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1649977179
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1649977179
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1649977179
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1649977179
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1649977179
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1649977179
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1649977179
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1649977179
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1649977179
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1649977179
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1649977179
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1649977179
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1649977179
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1649977179
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1649977179
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1649977179
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1649977179
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_505
timestamp 1649977179
transform 1 0 47564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_513
timestamp 1649977179
transform 1 0 48300 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_7
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_19
timestamp 1649977179
transform 1 0 2852 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1649977179
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1649977179
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1649977179
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1649977179
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1649977179
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1649977179
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1649977179
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1649977179
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1649977179
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1649977179
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1649977179
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1649977179
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1649977179
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1649977179
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1649977179
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1649977179
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1649977179
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1649977179
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1649977179
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1649977179
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1649977179
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1649977179
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1649977179
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1649977179
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1649977179
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_501
timestamp 1649977179
transform 1 0 47196 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_509
timestamp 1649977179
transform 1 0 47932 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_512
timestamp 1649977179
transform 1 0 48208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_13
timestamp 1649977179
transform 1 0 2300 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_25
timestamp 1649977179
transform 1 0 3404 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_37
timestamp 1649977179
transform 1 0 4508 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_49
timestamp 1649977179
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1649977179
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1649977179
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1649977179
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1649977179
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1649977179
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1649977179
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1649977179
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1649977179
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1649977179
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1649977179
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1649977179
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1649977179
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1649977179
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1649977179
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1649977179
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1649977179
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1649977179
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1649977179
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1649977179
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1649977179
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1649977179
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1649977179
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1649977179
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1649977179
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1649977179
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1649977179
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_505
timestamp 1649977179
transform 1 0 47564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_512
timestamp 1649977179
transform 1 0 48208 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1649977179
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1649977179
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1649977179
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1649977179
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1649977179
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1649977179
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1649977179
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1649977179
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1649977179
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1649977179
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1649977179
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1649977179
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1649977179
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1649977179
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1649977179
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1649977179
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1649977179
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1649977179
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1649977179
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1649977179
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1649977179
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1649977179
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1649977179
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1649977179
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1649977179
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1649977179
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_513
timestamp 1649977179
transform 1 0 48300 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1649977179
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1649977179
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1649977179
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1649977179
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1649977179
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1649977179
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1649977179
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1649977179
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1649977179
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1649977179
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1649977179
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1649977179
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1649977179
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1649977179
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1649977179
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1649977179
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1649977179
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1649977179
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1649977179
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1649977179
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1649977179
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1649977179
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1649977179
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1649977179
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1649977179
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1649977179
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1649977179
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_505
timestamp 1649977179
transform 1 0 47564 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_513
timestamp 1649977179
transform 1 0 48300 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_7
timestamp 1649977179
transform 1 0 1748 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_19
timestamp 1649977179
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1649977179
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1649977179
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1649977179
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1649977179
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1649977179
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1649977179
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1649977179
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1649977179
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1649977179
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1649977179
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1649977179
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1649977179
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1649977179
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1649977179
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1649977179
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1649977179
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1649977179
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1649977179
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1649977179
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1649977179
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1649977179
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1649977179
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1649977179
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1649977179
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1649977179
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1649977179
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1649977179
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_501
timestamp 1649977179
transform 1 0 47196 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_505
timestamp 1649977179
transform 1 0 47564 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_508
timestamp 1649977179
transform 1 0 47840 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_11
timestamp 1649977179
transform 1 0 2116 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_23
timestamp 1649977179
transform 1 0 3220 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_35
timestamp 1649977179
transform 1 0 4324 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_47
timestamp 1649977179
transform 1 0 5428 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1649977179
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1649977179
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1649977179
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1649977179
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1649977179
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1649977179
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1649977179
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1649977179
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1649977179
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1649977179
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1649977179
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1649977179
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1649977179
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1649977179
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1649977179
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1649977179
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1649977179
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1649977179
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1649977179
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1649977179
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1649977179
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1649977179
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1649977179
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1649977179
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1649977179
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_505
timestamp 1649977179
transform 1 0 47564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_512
timestamp 1649977179
transform 1 0 48208 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1649977179
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1649977179
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1649977179
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1649977179
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1649977179
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1649977179
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1649977179
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1649977179
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1649977179
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1649977179
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1649977179
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1649977179
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1649977179
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1649977179
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1649977179
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1649977179
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1649977179
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1649977179
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1649977179
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1649977179
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1649977179
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1649977179
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1649977179
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1649977179
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1649977179
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1649977179
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1649977179
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_513
timestamp 1649977179
transform 1 0 48300 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_7
timestamp 1649977179
transform 1 0 1748 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_19
timestamp 1649977179
transform 1 0 2852 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_31
timestamp 1649977179
transform 1 0 3956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_43
timestamp 1649977179
transform 1 0 5060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1649977179
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1649977179
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1649977179
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1649977179
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1649977179
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1649977179
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1649977179
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1649977179
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1649977179
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1649977179
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1649977179
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1649977179
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1649977179
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1649977179
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1649977179
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1649977179
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1649977179
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1649977179
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1649977179
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1649977179
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1649977179
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1649977179
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1649977179
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1649977179
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1649977179
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_505
timestamp 1649977179
transform 1 0 47564 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_513
timestamp 1649977179
transform 1 0 48300 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_13
timestamp 1649977179
transform 1 0 2300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_25
timestamp 1649977179
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1649977179
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1649977179
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1649977179
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1649977179
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1649977179
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1649977179
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1649977179
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1649977179
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1649977179
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1649977179
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1649977179
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1649977179
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1649977179
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1649977179
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1649977179
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1649977179
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1649977179
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1649977179
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1649977179
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1649977179
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1649977179
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1649977179
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1649977179
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1649977179
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1649977179
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1649977179
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1649977179
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_501
timestamp 1649977179
transform 1 0 47196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_504
timestamp 1649977179
transform 1 0 47472 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_512
timestamp 1649977179
transform 1 0 48208 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1649977179
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1649977179
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1649977179
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1649977179
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1649977179
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1649977179
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1649977179
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1649977179
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1649977179
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1649977179
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1649977179
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1649977179
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1649977179
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1649977179
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1649977179
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1649977179
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1649977179
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1649977179
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1649977179
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1649977179
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1649977179
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1649977179
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1649977179
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1649977179
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1649977179
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1649977179
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1649977179
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1649977179
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1649977179
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_505
timestamp 1649977179
transform 1 0 47564 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_513
timestamp 1649977179
transform 1 0 48300 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1649977179
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1649977179
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1649977179
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1649977179
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1649977179
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1649977179
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1649977179
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1649977179
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1649977179
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1649977179
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1649977179
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1649977179
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1649977179
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1649977179
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1649977179
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1649977179
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1649977179
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1649977179
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1649977179
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1649977179
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1649977179
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1649977179
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1649977179
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1649977179
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1649977179
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1649977179
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1649977179
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1649977179
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1649977179
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1649977179
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1649977179
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1649977179
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1649977179
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1649977179
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1649977179
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1649977179
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1649977179
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1649977179
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1649977179
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1649977179
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_513
timestamp 1649977179
transform 1 0 48300 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_7
timestamp 1649977179
transform 1 0 1748 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_19
timestamp 1649977179
transform 1 0 2852 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_31
timestamp 1649977179
transform 1 0 3956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_43
timestamp 1649977179
transform 1 0 5060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1649977179
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1649977179
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1649977179
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1649977179
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1649977179
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1649977179
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1649977179
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1649977179
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1649977179
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1649977179
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1649977179
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1649977179
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1649977179
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1649977179
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1649977179
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1649977179
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1649977179
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1649977179
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1649977179
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1649977179
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1649977179
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1649977179
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1649977179
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1649977179
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1649977179
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1649977179
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1649977179
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1649977179
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1649977179
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1649977179
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1649977179
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1649977179
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1649977179
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1649977179
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1649977179
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1649977179
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1649977179
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_505
timestamp 1649977179
transform 1 0 47564 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_513
timestamp 1649977179
transform 1 0 48300 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_11
timestamp 1649977179
transform 1 0 2116 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_23
timestamp 1649977179
transform 1 0 3220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1649977179
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1649977179
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1649977179
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1649977179
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1649977179
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1649977179
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1649977179
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1649977179
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1649977179
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1649977179
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1649977179
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1649977179
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1649977179
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1649977179
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1649977179
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1649977179
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1649977179
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1649977179
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1649977179
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1649977179
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1649977179
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1649977179
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1649977179
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1649977179
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1649977179
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1649977179
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1649977179
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1649977179
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1649977179
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1649977179
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1649977179
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1649977179
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1649977179
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1649977179
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1649977179
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1649977179
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1649977179
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1649977179
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1649977179
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_501
timestamp 1649977179
transform 1 0 47196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_504
timestamp 1649977179
transform 1 0 47472 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_512
timestamp 1649977179
transform 1 0 48208 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1649977179
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1649977179
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1649977179
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1649977179
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1649977179
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1649977179
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1649977179
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1649977179
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1649977179
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1649977179
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1649977179
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1649977179
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1649977179
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1649977179
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1649977179
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1649977179
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1649977179
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1649977179
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1649977179
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1649977179
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1649977179
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1649977179
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1649977179
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1649977179
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1649977179
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1649977179
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1649977179
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1649977179
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1649977179
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1649977179
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1649977179
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1649977179
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1649977179
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1649977179
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1649977179
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1649977179
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1649977179
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1649977179
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1649977179
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1649977179
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1649977179
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1649977179
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1649977179
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1649977179
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_505
timestamp 1649977179
transform 1 0 47564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_513
timestamp 1649977179
transform 1 0 48300 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1649977179
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1649977179
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1649977179
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1649977179
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1649977179
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1649977179
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1649977179
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1649977179
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1649977179
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1649977179
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1649977179
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1649977179
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1649977179
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1649977179
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1649977179
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1649977179
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1649977179
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1649977179
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1649977179
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1649977179
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1649977179
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1649977179
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1649977179
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1649977179
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1649977179
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1649977179
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1649977179
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1649977179
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1649977179
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1649977179
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1649977179
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1649977179
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1649977179
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1649977179
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1649977179
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1649977179
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1649977179
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1649977179
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1649977179
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1649977179
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1649977179
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1649977179
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_513
timestamp 1649977179
transform 1 0 48300 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1649977179
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1649977179
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1649977179
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1649977179
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1649977179
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1649977179
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1649977179
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1649977179
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1649977179
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1649977179
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1649977179
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1649977179
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1649977179
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1649977179
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1649977179
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1649977179
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1649977179
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1649977179
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1649977179
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1649977179
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1649977179
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1649977179
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1649977179
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1649977179
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1649977179
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1649977179
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1649977179
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1649977179
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1649977179
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1649977179
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1649977179
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1649977179
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1649977179
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1649977179
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1649977179
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1649977179
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1649977179
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1649977179
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1649977179
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1649977179
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1649977179
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1649977179
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1649977179
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1649977179
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_505
timestamp 1649977179
transform 1 0 47564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_509
timestamp 1649977179
transform 1 0 47932 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_512
timestamp 1649977179
transform 1 0 48208 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_7
timestamp 1649977179
transform 1 0 1748 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_13
timestamp 1649977179
transform 1 0 2300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_25
timestamp 1649977179
transform 1 0 3404 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1649977179
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1649977179
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1649977179
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1649977179
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1649977179
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1649977179
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1649977179
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1649977179
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1649977179
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1649977179
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1649977179
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1649977179
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1649977179
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1649977179
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1649977179
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1649977179
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_245
timestamp 1649977179
transform 1 0 23644 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1649977179
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_256
timestamp 1649977179
transform 1 0 24656 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_262
timestamp 1649977179
transform 1 0 25208 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_274
timestamp 1649977179
transform 1 0 26312 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_280
timestamp 1649977179
transform 1 0 26864 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_283
timestamp 1649977179
transform 1 0 27140 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_287
timestamp 1649977179
transform 1 0 27508 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_290
timestamp 1649977179
transform 1 0 27784 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_294
timestamp 1649977179
transform 1 0 28152 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_297
timestamp 1649977179
transform 1 0 28428 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_305
timestamp 1649977179
transform 1 0 29164 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1649977179
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1649977179
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1649977179
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1649977179
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1649977179
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1649977179
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1649977179
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1649977179
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1649977179
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1649977179
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1649977179
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1649977179
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1649977179
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1649977179
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1649977179
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1649977179
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1649977179
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1649977179
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_501
timestamp 1649977179
transform 1 0 47196 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_505
timestamp 1649977179
transform 1 0 47564 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_512
timestamp 1649977179
transform 1 0 48208 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1649977179
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1649977179
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1649977179
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1649977179
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1649977179
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1649977179
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1649977179
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1649977179
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1649977179
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1649977179
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1649977179
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1649977179
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1649977179
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1649977179
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1649977179
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1649977179
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1649977179
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1649977179
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1649977179
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_237
timestamp 1649977179
transform 1 0 22908 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_242
timestamp 1649977179
transform 1 0 23368 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_251
timestamp 1649977179
transform 1 0 24196 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1649977179
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_273
timestamp 1649977179
transform 1 0 26220 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1649977179
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_288
timestamp 1649977179
transform 1 0 27600 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_295
timestamp 1649977179
transform 1 0 28244 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_301
timestamp 1649977179
transform 1 0 28796 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_313
timestamp 1649977179
transform 1 0 29900 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_325
timestamp 1649977179
transform 1 0 31004 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_333
timestamp 1649977179
transform 1 0 31740 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1649977179
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1649977179
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1649977179
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1649977179
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1649977179
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1649977179
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1649977179
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1649977179
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1649977179
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1649977179
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1649977179
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1649977179
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1649977179
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1649977179
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1649977179
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1649977179
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_505
timestamp 1649977179
transform 1 0 47564 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_513
timestamp 1649977179
transform 1 0 48300 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1649977179
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1649977179
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1649977179
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1649977179
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1649977179
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1649977179
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1649977179
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1649977179
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1649977179
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1649977179
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1649977179
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1649977179
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1649977179
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1649977179
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1649977179
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1649977179
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1649977179
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_233
timestamp 1649977179
transform 1 0 22540 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_241
timestamp 1649977179
transform 1 0 23276 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_244
timestamp 1649977179
transform 1 0 23552 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_263
timestamp 1649977179
transform 1 0 25300 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_269
timestamp 1649977179
transform 1 0 25852 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_277
timestamp 1649977179
transform 1 0 26588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_281
timestamp 1649977179
transform 1 0 26956 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_289
timestamp 1649977179
transform 1 0 27692 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_296
timestamp 1649977179
transform 1 0 28336 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_302
timestamp 1649977179
transform 1 0 28888 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_321
timestamp 1649977179
transform 1 0 30636 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_327
timestamp 1649977179
transform 1 0 31188 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_330
timestamp 1649977179
transform 1 0 31464 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_336
timestamp 1649977179
transform 1 0 32016 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_348
timestamp 1649977179
transform 1 0 33120 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_360
timestamp 1649977179
transform 1 0 34224 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1649977179
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1649977179
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1649977179
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1649977179
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1649977179
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1649977179
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1649977179
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1649977179
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1649977179
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1649977179
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1649977179
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1649977179
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1649977179
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1649977179
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_513
timestamp 1649977179
transform 1 0 48300 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_7
timestamp 1649977179
transform 1 0 1748 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_19
timestamp 1649977179
transform 1 0 2852 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_31
timestamp 1649977179
transform 1 0 3956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_43
timestamp 1649977179
transform 1 0 5060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1649977179
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1649977179
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1649977179
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1649977179
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1649977179
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1649977179
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1649977179
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1649977179
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1649977179
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1649977179
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1649977179
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1649977179
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1649977179
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_205
timestamp 1649977179
transform 1 0 19964 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_213
timestamp 1649977179
transform 1 0 20700 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_221
timestamp 1649977179
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_227
timestamp 1649977179
transform 1 0 21988 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_231
timestamp 1649977179
transform 1 0 22356 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_234
timestamp 1649977179
transform 1 0 22632 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_246
timestamp 1649977179
transform 1 0 23736 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_254
timestamp 1649977179
transform 1 0 24472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_258
timestamp 1649977179
transform 1 0 24840 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_266
timestamp 1649977179
transform 1 0 25576 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_274
timestamp 1649977179
transform 1 0 26312 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_281
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_289
timestamp 1649977179
transform 1 0 27692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_301
timestamp 1649977179
transform 1 0 28796 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_309
timestamp 1649977179
transform 1 0 29532 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_318
timestamp 1649977179
transform 1 0 30360 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_324
timestamp 1649977179
transform 1 0 30912 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_328
timestamp 1649977179
transform 1 0 31280 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_339
timestamp 1649977179
transform 1 0 32292 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_345
timestamp 1649977179
transform 1 0 32844 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_357
timestamp 1649977179
transform 1 0 33948 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_369
timestamp 1649977179
transform 1 0 35052 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_381
timestamp 1649977179
transform 1 0 36156 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_389
timestamp 1649977179
transform 1 0 36892 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1649977179
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1649977179
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1649977179
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1649977179
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1649977179
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1649977179
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1649977179
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1649977179
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1649977179
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1649977179
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1649977179
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_505
timestamp 1649977179
transform 1 0 47564 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_509
timestamp 1649977179
transform 1 0 47932 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_512
timestamp 1649977179
transform 1 0 48208 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_11
timestamp 1649977179
transform 1 0 2116 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_23
timestamp 1649977179
transform 1 0 3220 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1649977179
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1649977179
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1649977179
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1649977179
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1649977179
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1649977179
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1649977179
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1649977179
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1649977179
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1649977179
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1649977179
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1649977179
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1649977179
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1649977179
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1649977179
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_197
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_202
timestamp 1649977179
transform 1 0 19688 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_209
timestamp 1649977179
transform 1 0 20332 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_213
timestamp 1649977179
transform 1 0 20700 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_216
timestamp 1649977179
transform 1 0 20976 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_222
timestamp 1649977179
transform 1 0 21528 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_226
timestamp 1649977179
transform 1 0 21896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_232
timestamp 1649977179
transform 1 0 22448 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_240
timestamp 1649977179
transform 1 0 23184 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_256
timestamp 1649977179
transform 1 0 24656 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_265
timestamp 1649977179
transform 1 0 25484 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_272
timestamp 1649977179
transform 1 0 26128 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_278
timestamp 1649977179
transform 1 0 26680 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_284
timestamp 1649977179
transform 1 0 27232 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_288
timestamp 1649977179
transform 1 0 27600 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_291
timestamp 1649977179
transform 1 0 27876 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_297
timestamp 1649977179
transform 1 0 28428 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_305
timestamp 1649977179
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_309
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_320
timestamp 1649977179
transform 1 0 30544 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_331
timestamp 1649977179
transform 1 0 31556 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_337
timestamp 1649977179
transform 1 0 32108 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_343
timestamp 1649977179
transform 1 0 32660 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_349
timestamp 1649977179
transform 1 0 33212 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_355
timestamp 1649977179
transform 1 0 33764 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1649977179
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1649977179
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1649977179
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1649977179
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1649977179
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1649977179
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1649977179
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1649977179
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1649977179
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1649977179
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1649977179
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1649977179
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1649977179
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1649977179
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_501
timestamp 1649977179
transform 1 0 47196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_512
timestamp 1649977179
transform 1 0 48208 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1649977179
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1649977179
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1649977179
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1649977179
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1649977179
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1649977179
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1649977179
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1649977179
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1649977179
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1649977179
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1649977179
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1649977179
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1649977179
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1649977179
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1649977179
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_181
timestamp 1649977179
transform 1 0 17756 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_189
timestamp 1649977179
transform 1 0 18492 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_194
timestamp 1649977179
transform 1 0 18952 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_200
timestamp 1649977179
transform 1 0 19504 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_203
timestamp 1649977179
transform 1 0 19780 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_212
timestamp 1649977179
transform 1 0 20608 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_216
timestamp 1649977179
transform 1 0 20976 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1649977179
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_231
timestamp 1649977179
transform 1 0 22356 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_235
timestamp 1649977179
transform 1 0 22724 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_243
timestamp 1649977179
transform 1 0 23460 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_252
timestamp 1649977179
transform 1 0 24288 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_263
timestamp 1649977179
transform 1 0 25300 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_272
timestamp 1649977179
transform 1 0 26128 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_289
timestamp 1649977179
transform 1 0 27692 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_302
timestamp 1649977179
transform 1 0 28888 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_313
timestamp 1649977179
transform 1 0 29900 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_320
timestamp 1649977179
transform 1 0 30544 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_327
timestamp 1649977179
transform 1 0 31188 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1649977179
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_342
timestamp 1649977179
transform 1 0 32568 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_346
timestamp 1649977179
transform 1 0 32936 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_360
timestamp 1649977179
transform 1 0 34224 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_366
timestamp 1649977179
transform 1 0 34776 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_378
timestamp 1649977179
transform 1 0 35880 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_390
timestamp 1649977179
transform 1 0 36984 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1649977179
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1649977179
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1649977179
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1649977179
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1649977179
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1649977179
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1649977179
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1649977179
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1649977179
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1649977179
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1649977179
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_505
timestamp 1649977179
transform 1 0 47564 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_509
timestamp 1649977179
transform 1 0 47932 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_512
timestamp 1649977179
transform 1 0 48208 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1649977179
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1649977179
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1649977179
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1649977179
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1649977179
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1649977179
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1649977179
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1649977179
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1649977179
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1649977179
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1649977179
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1649977179
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1649977179
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1649977179
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_189
timestamp 1649977179
transform 1 0 18492 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1649977179
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_201
timestamp 1649977179
transform 1 0 19596 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_205
timestamp 1649977179
transform 1 0 19964 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_209
timestamp 1649977179
transform 1 0 20332 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_212
timestamp 1649977179
transform 1 0 20608 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_218
timestamp 1649977179
transform 1 0 21160 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_228
timestamp 1649977179
transform 1 0 22080 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_240
timestamp 1649977179
transform 1 0 23184 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_247
timestamp 1649977179
transform 1 0 23828 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1649977179
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_255
timestamp 1649977179
transform 1 0 24564 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_264
timestamp 1649977179
transform 1 0 25392 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_270
timestamp 1649977179
transform 1 0 25944 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_276
timestamp 1649977179
transform 1 0 26496 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_288
timestamp 1649977179
transform 1 0 27600 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_296
timestamp 1649977179
transform 1 0 28336 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_302
timestamp 1649977179
transform 1 0 28888 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_311
timestamp 1649977179
transform 1 0 29716 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_321
timestamp 1649977179
transform 1 0 30636 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_330
timestamp 1649977179
transform 1 0 31464 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_336
timestamp 1649977179
transform 1 0 32016 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_340
timestamp 1649977179
transform 1 0 32384 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_344
timestamp 1649977179
transform 1 0 32752 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_353
timestamp 1649977179
transform 1 0 33580 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_359
timestamp 1649977179
transform 1 0 34132 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1649977179
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1649977179
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1649977179
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1649977179
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1649977179
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1649977179
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1649977179
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1649977179
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1649977179
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1649977179
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1649977179
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1649977179
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1649977179
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1649977179
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_501
timestamp 1649977179
transform 1 0 47196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_512
timestamp 1649977179
transform 1 0 48208 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_7
timestamp 1649977179
transform 1 0 1748 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_13
timestamp 1649977179
transform 1 0 2300 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_25
timestamp 1649977179
transform 1 0 3404 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_37
timestamp 1649977179
transform 1 0 4508 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_49
timestamp 1649977179
transform 1 0 5612 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1649977179
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1649977179
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1649977179
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1649977179
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1649977179
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1649977179
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1649977179
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1649977179
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1649977179
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1649977179
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1649977179
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1649977179
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_169
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_177
timestamp 1649977179
transform 1 0 17388 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_182
timestamp 1649977179
transform 1 0 17848 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_190
timestamp 1649977179
transform 1 0 18584 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_194
timestamp 1649977179
transform 1 0 18952 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_203
timestamp 1649977179
transform 1 0 19780 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_213
timestamp 1649977179
transform 1 0 20700 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_217
timestamp 1649977179
transform 1 0 21068 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1649977179
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_229
timestamp 1649977179
transform 1 0 22172 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_232
timestamp 1649977179
transform 1 0 22448 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_239
timestamp 1649977179
transform 1 0 23092 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_248
timestamp 1649977179
transform 1 0 23920 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_254
timestamp 1649977179
transform 1 0 24472 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_262
timestamp 1649977179
transform 1 0 25208 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_47_274
timestamp 1649977179
transform 1 0 26312 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_281
timestamp 1649977179
transform 1 0 26956 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_285
timestamp 1649977179
transform 1 0 27324 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_293
timestamp 1649977179
transform 1 0 28060 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_300
timestamp 1649977179
transform 1 0 28704 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_306
timestamp 1649977179
transform 1 0 29256 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_312
timestamp 1649977179
transform 1 0 29808 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_319
timestamp 1649977179
transform 1 0 30452 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_326
timestamp 1649977179
transform 1 0 31096 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1649977179
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_337
timestamp 1649977179
transform 1 0 32108 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_351
timestamp 1649977179
transform 1 0 33396 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_359
timestamp 1649977179
transform 1 0 34132 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_365
timestamp 1649977179
transform 1 0 34684 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_371
timestamp 1649977179
transform 1 0 35236 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_383
timestamp 1649977179
transform 1 0 36340 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1649977179
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1649977179
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1649977179
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1649977179
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1649977179
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1649977179
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1649977179
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1649977179
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1649977179
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1649977179
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1649977179
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1649977179
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_505
timestamp 1649977179
transform 1 0 47564 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_513
timestamp 1649977179
transform 1 0 48300 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1649977179
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1649977179
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1649977179
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1649977179
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1649977179
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1649977179
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1649977179
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1649977179
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1649977179
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1649977179
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1649977179
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1649977179
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_155
timestamp 1649977179
transform 1 0 15364 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_161
timestamp 1649977179
transform 1 0 15916 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_169
timestamp 1649977179
transform 1 0 16652 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_175
timestamp 1649977179
transform 1 0 17204 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_185
timestamp 1649977179
transform 1 0 18124 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_189
timestamp 1649977179
transform 1 0 18492 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1649977179
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_197
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_201
timestamp 1649977179
transform 1 0 19596 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_207
timestamp 1649977179
transform 1 0 20148 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_218
timestamp 1649977179
transform 1 0 21160 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_222
timestamp 1649977179
transform 1 0 21528 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_228
timestamp 1649977179
transform 1 0 22080 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_237
timestamp 1649977179
transform 1 0 22908 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_243
timestamp 1649977179
transform 1 0 23460 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1649977179
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_253
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_261
timestamp 1649977179
transform 1 0 25116 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_269
timestamp 1649977179
transform 1 0 25852 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_275
timestamp 1649977179
transform 1 0 26404 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_284
timestamp 1649977179
transform 1 0 27232 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_297
timestamp 1649977179
transform 1 0 28428 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_303
timestamp 1649977179
transform 1 0 28980 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1649977179
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_312
timestamp 1649977179
transform 1 0 29808 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_316
timestamp 1649977179
transform 1 0 30176 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_322
timestamp 1649977179
transform 1 0 30728 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_338
timestamp 1649977179
transform 1 0 32200 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_348
timestamp 1649977179
transform 1 0 33120 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_354
timestamp 1649977179
transform 1 0 33672 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_360
timestamp 1649977179
transform 1 0 34224 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_372
timestamp 1649977179
transform 1 0 35328 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_379
timestamp 1649977179
transform 1 0 35972 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_391
timestamp 1649977179
transform 1 0 37076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_403
timestamp 1649977179
transform 1 0 38180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_415
timestamp 1649977179
transform 1 0 39284 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1649977179
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1649977179
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1649977179
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1649977179
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1649977179
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1649977179
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1649977179
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1649977179
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1649977179
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1649977179
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_513
timestamp 1649977179
transform 1 0 48300 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1649977179
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1649977179
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1649977179
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1649977179
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1649977179
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1649977179
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1649977179
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1649977179
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1649977179
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1649977179
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1649977179
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1649977179
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1649977179
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_151
timestamp 1649977179
transform 1 0 14996 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_157
timestamp 1649977179
transform 1 0 15548 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1649977179
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_174
timestamp 1649977179
transform 1 0 17112 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_178
timestamp 1649977179
transform 1 0 17480 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_188
timestamp 1649977179
transform 1 0 18400 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_198
timestamp 1649977179
transform 1 0 19320 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_206
timestamp 1649977179
transform 1 0 20056 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1649977179
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1649977179
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_225
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_234
timestamp 1649977179
transform 1 0 22632 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_242
timestamp 1649977179
transform 1 0 23368 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_249
timestamp 1649977179
transform 1 0 24012 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_253
timestamp 1649977179
transform 1 0 24380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_260
timestamp 1649977179
transform 1 0 25024 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_268
timestamp 1649977179
transform 1 0 25760 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_276
timestamp 1649977179
transform 1 0 26496 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_287
timestamp 1649977179
transform 1 0 27508 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_298
timestamp 1649977179
transform 1 0 28520 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_306
timestamp 1649977179
transform 1 0 29256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_311
timestamp 1649977179
transform 1 0 29716 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_320
timestamp 1649977179
transform 1 0 30544 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_328
timestamp 1649977179
transform 1 0 31280 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_49_339
timestamp 1649977179
transform 1 0 32292 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_350
timestamp 1649977179
transform 1 0 33304 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_358
timestamp 1649977179
transform 1 0 34040 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_366
timestamp 1649977179
transform 1 0 34776 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_378
timestamp 1649977179
transform 1 0 35880 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_384
timestamp 1649977179
transform 1 0 36432 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1649977179
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1649977179
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1649977179
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1649977179
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1649977179
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1649977179
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1649977179
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1649977179
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1649977179
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1649977179
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1649977179
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1649977179
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_505
timestamp 1649977179
transform 1 0 47564 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_509
timestamp 1649977179
transform 1 0 47932 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_512
timestamp 1649977179
transform 1 0 48208 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1649977179
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_7
timestamp 1649977179
transform 1 0 1748 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_19
timestamp 1649977179
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1649977179
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1649977179
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1649977179
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1649977179
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1649977179
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1649977179
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1649977179
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1649977179
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1649977179
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1649977179
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1649977179
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_146
timestamp 1649977179
transform 1 0 14536 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_152
timestamp 1649977179
transform 1 0 15088 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_158
timestamp 1649977179
transform 1 0 15640 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_167
timestamp 1649977179
transform 1 0 16468 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_174
timestamp 1649977179
transform 1 0 17112 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_180
timestamp 1649977179
transform 1 0 17664 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_183
timestamp 1649977179
transform 1 0 17940 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_192
timestamp 1649977179
transform 1 0 18768 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_197
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_204
timestamp 1649977179
transform 1 0 19872 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_213
timestamp 1649977179
transform 1 0 20700 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_217
timestamp 1649977179
transform 1 0 21068 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_221
timestamp 1649977179
transform 1 0 21436 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_228
timestamp 1649977179
transform 1 0 22080 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_239
timestamp 1649977179
transform 1 0 23092 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_247
timestamp 1649977179
transform 1 0 23828 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1649977179
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_255
timestamp 1649977179
transform 1 0 24564 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_266
timestamp 1649977179
transform 1 0 25576 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_272
timestamp 1649977179
transform 1 0 26128 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_285
timestamp 1649977179
transform 1 0 27324 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_297
timestamp 1649977179
transform 1 0 28428 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_304
timestamp 1649977179
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_313
timestamp 1649977179
transform 1 0 29900 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_322
timestamp 1649977179
transform 1 0 30728 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_331
timestamp 1649977179
transform 1 0 31556 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_337
timestamp 1649977179
transform 1 0 32108 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_344
timestamp 1649977179
transform 1 0 32752 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_354
timestamp 1649977179
transform 1 0 33672 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_360
timestamp 1649977179
transform 1 0 34224 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_367
timestamp 1649977179
transform 1 0 34868 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_381
timestamp 1649977179
transform 1 0 36156 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_390
timestamp 1649977179
transform 1 0 36984 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_402
timestamp 1649977179
transform 1 0 38088 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_414
timestamp 1649977179
transform 1 0 39192 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1649977179
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1649977179
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1649977179
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1649977179
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1649977179
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1649977179
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1649977179
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1649977179
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_501
timestamp 1649977179
transform 1 0 47196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_512
timestamp 1649977179
transform 1 0 48208 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_11
timestamp 1649977179
transform 1 0 2116 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_23
timestamp 1649977179
transform 1 0 3220 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_35
timestamp 1649977179
transform 1 0 4324 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_47
timestamp 1649977179
transform 1 0 5428 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1649977179
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1649977179
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1649977179
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1649977179
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1649977179
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1649977179
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_113
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_117
timestamp 1649977179
transform 1 0 11868 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_120
timestamp 1649977179
transform 1 0 12144 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_126
timestamp 1649977179
transform 1 0 12696 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_132
timestamp 1649977179
transform 1 0 13248 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_138
timestamp 1649977179
transform 1 0 13800 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_144
timestamp 1649977179
transform 1 0 14352 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_150
timestamp 1649977179
transform 1 0 14904 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_160
timestamp 1649977179
transform 1 0 15824 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_175
timestamp 1649977179
transform 1 0 17204 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_184
timestamp 1649977179
transform 1 0 18032 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_192
timestamp 1649977179
transform 1 0 18768 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_196
timestamp 1649977179
transform 1 0 19136 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_204
timestamp 1649977179
transform 1 0 19872 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_220
timestamp 1649977179
transform 1 0 21344 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_225
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_229
timestamp 1649977179
transform 1 0 22172 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_232
timestamp 1649977179
transform 1 0 22448 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_236
timestamp 1649977179
transform 1 0 22816 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_239
timestamp 1649977179
transform 1 0 23092 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_254
timestamp 1649977179
transform 1 0 24472 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_264
timestamp 1649977179
transform 1 0 25392 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_271
timestamp 1649977179
transform 1 0 26036 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1649977179
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_283
timestamp 1649977179
transform 1 0 27140 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_291
timestamp 1649977179
transform 1 0 27876 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_299
timestamp 1649977179
transform 1 0 28612 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_305
timestamp 1649977179
transform 1 0 29164 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_313
timestamp 1649977179
transform 1 0 29900 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_320
timestamp 1649977179
transform 1 0 30544 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_326
timestamp 1649977179
transform 1 0 31096 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_332
timestamp 1649977179
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_337
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_344
timestamp 1649977179
transform 1 0 32752 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_350
timestamp 1649977179
transform 1 0 33304 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_354
timestamp 1649977179
transform 1 0 33672 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_361
timestamp 1649977179
transform 1 0 34316 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_372
timestamp 1649977179
transform 1 0 35328 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_380
timestamp 1649977179
transform 1 0 36064 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_388
timestamp 1649977179
transform 1 0 36800 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_395
timestamp 1649977179
transform 1 0 37444 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_407
timestamp 1649977179
transform 1 0 38548 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_419
timestamp 1649977179
transform 1 0 39652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_431
timestamp 1649977179
transform 1 0 40756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_443
timestamp 1649977179
transform 1 0 41860 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1649977179
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1649977179
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1649977179
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1649977179
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1649977179
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1649977179
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1649977179
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1649977179
transform 1 0 47564 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_513
timestamp 1649977179
transform 1 0 48300 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1649977179
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1649977179
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1649977179
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1649977179
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1649977179
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1649977179
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1649977179
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1649977179
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1649977179
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_109
timestamp 1649977179
transform 1 0 11132 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_112
timestamp 1649977179
transform 1 0 11408 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_118
timestamp 1649977179
transform 1 0 11960 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_125
timestamp 1649977179
transform 1 0 12604 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_132
timestamp 1649977179
transform 1 0 13248 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_52_146
timestamp 1649977179
transform 1 0 14536 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_152
timestamp 1649977179
transform 1 0 15088 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_159
timestamp 1649977179
transform 1 0 15732 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_169
timestamp 1649977179
transform 1 0 16652 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_181
timestamp 1649977179
transform 1 0 17756 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_189
timestamp 1649977179
transform 1 0 18492 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp 1649977179
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_197
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_201
timestamp 1649977179
transform 1 0 19596 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_206
timestamp 1649977179
transform 1 0 20056 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_215
timestamp 1649977179
transform 1 0 20884 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_226
timestamp 1649977179
transform 1 0 21896 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_234
timestamp 1649977179
transform 1 0 22632 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_238
timestamp 1649977179
transform 1 0 23000 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_241
timestamp 1649977179
transform 1 0 23276 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_245
timestamp 1649977179
transform 1 0 23644 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1649977179
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_256
timestamp 1649977179
transform 1 0 24656 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_260
timestamp 1649977179
transform 1 0 25024 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_263
timestamp 1649977179
transform 1 0 25300 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_269
timestamp 1649977179
transform 1 0 25852 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_272
timestamp 1649977179
transform 1 0 26128 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_278
timestamp 1649977179
transform 1 0 26680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_282
timestamp 1649977179
transform 1 0 27048 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_286
timestamp 1649977179
transform 1 0 27416 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_292
timestamp 1649977179
transform 1 0 27968 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_298
timestamp 1649977179
transform 1 0 28520 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_304
timestamp 1649977179
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_312
timestamp 1649977179
transform 1 0 29808 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_318
timestamp 1649977179
transform 1 0 30360 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_327
timestamp 1649977179
transform 1 0 31188 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_348
timestamp 1649977179
transform 1 0 33120 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_355
timestamp 1649977179
transform 1 0 33764 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1649977179
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_365
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_369
timestamp 1649977179
transform 1 0 35052 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_375
timestamp 1649977179
transform 1 0 35604 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_381
timestamp 1649977179
transform 1 0 36156 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_387
timestamp 1649977179
transform 1 0 36708 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_393
timestamp 1649977179
transform 1 0 37260 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_399
timestamp 1649977179
transform 1 0 37812 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_405
timestamp 1649977179
transform 1 0 38364 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_411
timestamp 1649977179
transform 1 0 38916 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1649977179
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1649977179
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1649977179
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1649977179
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1649977179
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1649977179
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1649977179
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1649977179
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1649977179
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1649977179
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_513
timestamp 1649977179
transform 1 0 48300 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1649977179
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1649977179
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1649977179
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1649977179
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1649977179
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1649977179
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1649977179
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1649977179
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_105
timestamp 1649977179
transform 1 0 10764 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_108
timestamp 1649977179
transform 1 0 11040 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_118
timestamp 1649977179
transform 1 0 11960 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_127
timestamp 1649977179
transform 1 0 12788 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_133
timestamp 1649977179
transform 1 0 13340 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_140
timestamp 1649977179
transform 1 0 13984 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_148
timestamp 1649977179
transform 1 0 14720 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_153
timestamp 1649977179
transform 1 0 15180 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_162
timestamp 1649977179
transform 1 0 16008 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1649977179
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_173
timestamp 1649977179
transform 1 0 17020 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_183
timestamp 1649977179
transform 1 0 17940 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_191
timestamp 1649977179
transform 1 0 18676 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_198
timestamp 1649977179
transform 1 0 19320 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_205
timestamp 1649977179
transform 1 0 19964 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_211
timestamp 1649977179
transform 1 0 20516 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_218
timestamp 1649977179
transform 1 0 21160 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_225
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_228
timestamp 1649977179
transform 1 0 22080 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_237
timestamp 1649977179
transform 1 0 22908 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_244
timestamp 1649977179
transform 1 0 23552 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_252
timestamp 1649977179
transform 1 0 24288 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_261
timestamp 1649977179
transform 1 0 25116 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_268
timestamp 1649977179
transform 1 0 25760 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_275
timestamp 1649977179
transform 1 0 26404 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1649977179
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_283
timestamp 1649977179
transform 1 0 27140 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_291
timestamp 1649977179
transform 1 0 27876 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_298
timestamp 1649977179
transform 1 0 28520 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_304
timestamp 1649977179
transform 1 0 29072 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_314
timestamp 1649977179
transform 1 0 29992 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_321
timestamp 1649977179
transform 1 0 30636 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_328
timestamp 1649977179
transform 1 0 31280 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_337
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_347
timestamp 1649977179
transform 1 0 33028 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_354
timestamp 1649977179
transform 1 0 33672 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_364
timestamp 1649977179
transform 1 0 34592 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_375
timestamp 1649977179
transform 1 0 35604 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_381
timestamp 1649977179
transform 1 0 36156 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_387
timestamp 1649977179
transform 1 0 36708 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1649977179
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_399
timestamp 1649977179
transform 1 0 37812 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_405
timestamp 1649977179
transform 1 0 38364 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_411
timestamp 1649977179
transform 1 0 38916 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_417
timestamp 1649977179
transform 1 0 39468 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_423
timestamp 1649977179
transform 1 0 40020 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1649977179
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1649977179
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1649977179
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1649977179
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1649977179
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1649977179
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1649977179
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1649977179
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1649977179
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1649977179
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1649977179
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1649977179
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_7
timestamp 1649977179
transform 1 0 1748 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_19
timestamp 1649977179
transform 1 0 2852 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1649977179
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1649977179
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1649977179
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1649977179
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1649977179
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_97
timestamp 1649977179
transform 1 0 10028 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_100
timestamp 1649977179
transform 1 0 10304 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_106
timestamp 1649977179
transform 1 0 10856 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_112
timestamp 1649977179
transform 1 0 11408 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_118
timestamp 1649977179
transform 1 0 11960 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_126
timestamp 1649977179
transform 1 0 12696 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_130
timestamp 1649977179
transform 1 0 13064 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_136
timestamp 1649977179
transform 1 0 13616 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_145
timestamp 1649977179
transform 1 0 14444 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_154
timestamp 1649977179
transform 1 0 15272 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_162
timestamp 1649977179
transform 1 0 16008 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_170
timestamp 1649977179
transform 1 0 16744 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_178
timestamp 1649977179
transform 1 0 17480 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_190
timestamp 1649977179
transform 1 0 18584 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_200
timestamp 1649977179
transform 1 0 19504 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_206
timestamp 1649977179
transform 1 0 20056 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_218
timestamp 1649977179
transform 1 0 21160 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_222
timestamp 1649977179
transform 1 0 21528 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_228
timestamp 1649977179
transform 1 0 22080 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_237
timestamp 1649977179
transform 1 0 22908 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_248
timestamp 1649977179
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_262
timestamp 1649977179
transform 1 0 25208 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_271
timestamp 1649977179
transform 1 0 26036 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_284
timestamp 1649977179
transform 1 0 27232 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_292
timestamp 1649977179
transform 1 0 27968 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_296
timestamp 1649977179
transform 1 0 28336 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1649977179
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_316
timestamp 1649977179
transform 1 0 30176 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_323
timestamp 1649977179
transform 1 0 30820 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_329
timestamp 1649977179
transform 1 0 31372 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_340
timestamp 1649977179
transform 1 0 32384 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_349
timestamp 1649977179
transform 1 0 33212 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_355
timestamp 1649977179
transform 1 0 33764 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_360
timestamp 1649977179
transform 1 0 34224 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_365
timestamp 1649977179
transform 1 0 34684 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_374
timestamp 1649977179
transform 1 0 35512 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_380
timestamp 1649977179
transform 1 0 36064 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_398
timestamp 1649977179
transform 1 0 37720 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_404
timestamp 1649977179
transform 1 0 38272 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_410
timestamp 1649977179
transform 1 0 38824 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_416
timestamp 1649977179
transform 1 0 39376 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_423
timestamp 1649977179
transform 1 0 40020 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_429
timestamp 1649977179
transform 1 0 40572 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_435
timestamp 1649977179
transform 1 0 41124 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_447
timestamp 1649977179
transform 1 0 42228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_459
timestamp 1649977179
transform 1 0 43332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_471
timestamp 1649977179
transform 1 0 44436 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1649977179
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1649977179
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1649977179
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_501
timestamp 1649977179
transform 1 0 47196 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_505
timestamp 1649977179
transform 1 0 47564 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_508
timestamp 1649977179
transform 1 0 47840 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_3
timestamp 1649977179
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_11
timestamp 1649977179
transform 1 0 2116 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_23
timestamp 1649977179
transform 1 0 3220 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_35
timestamp 1649977179
transform 1 0 4324 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_47
timestamp 1649977179
transform 1 0 5428 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1649977179
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1649977179
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1649977179
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_93
timestamp 1649977179
transform 1 0 9660 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_99
timestamp 1649977179
transform 1 0 10212 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_102
timestamp 1649977179
transform 1 0 10488 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_108
timestamp 1649977179
transform 1 0 11040 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_117
timestamp 1649977179
transform 1 0 11868 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_120
timestamp 1649977179
transform 1 0 12144 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_131
timestamp 1649977179
transform 1 0 13156 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_140
timestamp 1649977179
transform 1 0 13984 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_147
timestamp 1649977179
transform 1 0 14628 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_164
timestamp 1649977179
transform 1 0 16192 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_174
timestamp 1649977179
transform 1 0 17112 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_180
timestamp 1649977179
transform 1 0 17664 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_189
timestamp 1649977179
transform 1 0 18492 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_198
timestamp 1649977179
transform 1 0 19320 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_207
timestamp 1649977179
transform 1 0 20148 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1649977179
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_227
timestamp 1649977179
transform 1 0 21988 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_234
timestamp 1649977179
transform 1 0 22632 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_246
timestamp 1649977179
transform 1 0 23736 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_254
timestamp 1649977179
transform 1 0 24472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_259
timestamp 1649977179
transform 1 0 24932 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_266
timestamp 1649977179
transform 1 0 25576 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1649977179
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1649977179
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_284
timestamp 1649977179
transform 1 0 27232 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_295
timestamp 1649977179
transform 1 0 28244 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_305
timestamp 1649977179
transform 1 0 29164 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_317
timestamp 1649977179
transform 1 0 30268 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_325
timestamp 1649977179
transform 1 0 31004 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_331
timestamp 1649977179
transform 1 0 31556 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1649977179
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_337
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_349
timestamp 1649977179
transform 1 0 33212 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_359
timestamp 1649977179
transform 1 0 34132 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_363
timestamp 1649977179
transform 1 0 34500 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_370
timestamp 1649977179
transform 1 0 35144 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_379
timestamp 1649977179
transform 1 0 35972 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_386
timestamp 1649977179
transform 1 0 36616 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_398
timestamp 1649977179
transform 1 0 37720 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_407
timestamp 1649977179
transform 1 0 38548 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_413
timestamp 1649977179
transform 1 0 39100 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_419
timestamp 1649977179
transform 1 0 39652 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_425
timestamp 1649977179
transform 1 0 40204 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_431
timestamp 1649977179
transform 1 0 40756 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_437
timestamp 1649977179
transform 1 0 41308 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_443
timestamp 1649977179
transform 1 0 41860 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1649977179
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1649977179
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1649977179
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1649977179
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1649977179
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1649977179
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1649977179
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_505
timestamp 1649977179
transform 1 0 47564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_512
timestamp 1649977179
transform 1 0 48208 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1649977179
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1649977179
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1649977179
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1649977179
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1649977179
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1649977179
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1649977179
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_97
timestamp 1649977179
transform 1 0 10028 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_103
timestamp 1649977179
transform 1 0 10580 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_109
timestamp 1649977179
transform 1 0 11132 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_116
timestamp 1649977179
transform 1 0 11776 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_124
timestamp 1649977179
transform 1 0 12512 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_132
timestamp 1649977179
transform 1 0 13248 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_141
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_145
timestamp 1649977179
transform 1 0 14444 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_151
timestamp 1649977179
transform 1 0 14996 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_167
timestamp 1649977179
transform 1 0 16468 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_179
timestamp 1649977179
transform 1 0 17572 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_186
timestamp 1649977179
transform 1 0 18216 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1649977179
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_199
timestamp 1649977179
transform 1 0 19412 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_208
timestamp 1649977179
transform 1 0 20240 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_212
timestamp 1649977179
transform 1 0 20608 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_216
timestamp 1649977179
transform 1 0 20976 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_227
timestamp 1649977179
transform 1 0 21988 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_237
timestamp 1649977179
transform 1 0 22908 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_244
timestamp 1649977179
transform 1 0 23552 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_253
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_260
timestamp 1649977179
transform 1 0 25024 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_271
timestamp 1649977179
transform 1 0 26036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_277
timestamp 1649977179
transform 1 0 26588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_281
timestamp 1649977179
transform 1 0 26956 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_290
timestamp 1649977179
transform 1 0 27784 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1649977179
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1649977179
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_311
timestamp 1649977179
transform 1 0 29716 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_322
timestamp 1649977179
transform 1 0 30728 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_326
timestamp 1649977179
transform 1 0 31096 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_334
timestamp 1649977179
transform 1 0 31832 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_346
timestamp 1649977179
transform 1 0 32936 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_355
timestamp 1649977179
transform 1 0 33764 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1649977179
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_371
timestamp 1649977179
transform 1 0 35236 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_377
timestamp 1649977179
transform 1 0 35788 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_383
timestamp 1649977179
transform 1 0 36340 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_389
timestamp 1649977179
transform 1 0 36892 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_398
timestamp 1649977179
transform 1 0 37720 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_405
timestamp 1649977179
transform 1 0 38364 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_411
timestamp 1649977179
transform 1 0 38916 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1649977179
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_428
timestamp 1649977179
transform 1 0 40480 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_434
timestamp 1649977179
transform 1 0 41032 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_440
timestamp 1649977179
transform 1 0 41584 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_446
timestamp 1649977179
transform 1 0 42136 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_452
timestamp 1649977179
transform 1 0 42688 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_464
timestamp 1649977179
transform 1 0 43792 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1649977179
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1649977179
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1649977179
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_513
timestamp 1649977179
transform 1 0 48300 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1649977179
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1649977179
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1649977179
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1649977179
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1649977179
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1649977179
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1649977179
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1649977179
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_93
timestamp 1649977179
transform 1 0 9660 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_96
timestamp 1649977179
transform 1 0 9936 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_102
timestamp 1649977179
transform 1 0 10488 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_108
timestamp 1649977179
transform 1 0 11040 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_118
timestamp 1649977179
transform 1 0 11960 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_131
timestamp 1649977179
transform 1 0 13156 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_139
timestamp 1649977179
transform 1 0 13892 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_145
timestamp 1649977179
transform 1 0 14444 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_152
timestamp 1649977179
transform 1 0 15088 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_159
timestamp 1649977179
transform 1 0 15732 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1649977179
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_173
timestamp 1649977179
transform 1 0 17020 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_179
timestamp 1649977179
transform 1 0 17572 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_186
timestamp 1649977179
transform 1 0 18216 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_198
timestamp 1649977179
transform 1 0 19320 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_210
timestamp 1649977179
transform 1 0 20424 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_219
timestamp 1649977179
transform 1 0 21252 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1649977179
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_225
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_229
timestamp 1649977179
transform 1 0 22172 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_232
timestamp 1649977179
transform 1 0 22448 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_239
timestamp 1649977179
transform 1 0 23092 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_243
timestamp 1649977179
transform 1 0 23460 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_246
timestamp 1649977179
transform 1 0 23736 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_254
timestamp 1649977179
transform 1 0 24472 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_262
timestamp 1649977179
transform 1 0 25208 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_269
timestamp 1649977179
transform 1 0 25852 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_273
timestamp 1649977179
transform 1 0 26220 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_276
timestamp 1649977179
transform 1 0 26496 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_290
timestamp 1649977179
transform 1 0 27784 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_296
timestamp 1649977179
transform 1 0 28336 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_302
timestamp 1649977179
transform 1 0 28888 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_312
timestamp 1649977179
transform 1 0 29808 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_323
timestamp 1649977179
transform 1 0 30820 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_330
timestamp 1649977179
transform 1 0 31464 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_337
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_343
timestamp 1649977179
transform 1 0 32660 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_349
timestamp 1649977179
transform 1 0 33212 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_355
timestamp 1649977179
transform 1 0 33764 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_359
timestamp 1649977179
transform 1 0 34132 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_365
timestamp 1649977179
transform 1 0 34684 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_376
timestamp 1649977179
transform 1 0 35696 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_383
timestamp 1649977179
transform 1 0 36340 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1649977179
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_400
timestamp 1649977179
transform 1 0 37904 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_409
timestamp 1649977179
transform 1 0 38732 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_423
timestamp 1649977179
transform 1 0 40020 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_435
timestamp 1649977179
transform 1 0 41124 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1649977179
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1649977179
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_451
timestamp 1649977179
transform 1 0 42596 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_457
timestamp 1649977179
transform 1 0 43148 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_463
timestamp 1649977179
transform 1 0 43700 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_475
timestamp 1649977179
transform 1 0 44804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_487
timestamp 1649977179
transform 1 0 45908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_499
timestamp 1649977179
transform 1 0 47012 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1649977179
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_505
timestamp 1649977179
transform 1 0 47564 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_509
timestamp 1649977179
transform 1 0 47932 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_512
timestamp 1649977179
transform 1 0 48208 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_3
timestamp 1649977179
transform 1 0 1380 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_7
timestamp 1649977179
transform 1 0 1748 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_19
timestamp 1649977179
transform 1 0 2852 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1649977179
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1649977179
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1649977179
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1649977179
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1649977179
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1649977179
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_85
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_93
timestamp 1649977179
transform 1 0 9660 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_96
timestamp 1649977179
transform 1 0 9936 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_102
timestamp 1649977179
transform 1 0 10488 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_109
timestamp 1649977179
transform 1 0 11132 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_121
timestamp 1649977179
transform 1 0 12236 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_136
timestamp 1649977179
transform 1 0 13616 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_141
timestamp 1649977179
transform 1 0 14076 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_148
timestamp 1649977179
transform 1 0 14720 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_156
timestamp 1649977179
transform 1 0 15456 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_165
timestamp 1649977179
transform 1 0 16284 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_175
timestamp 1649977179
transform 1 0 17204 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_184
timestamp 1649977179
transform 1 0 18032 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_192
timestamp 1649977179
transform 1 0 18768 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_204
timestamp 1649977179
transform 1 0 19872 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_210
timestamp 1649977179
transform 1 0 20424 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_215
timestamp 1649977179
transform 1 0 20884 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_58_226
timestamp 1649977179
transform 1 0 21896 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_241
timestamp 1649977179
transform 1 0 23276 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_245
timestamp 1649977179
transform 1 0 23644 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_248
timestamp 1649977179
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_253
timestamp 1649977179
transform 1 0 24380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_264
timestamp 1649977179
transform 1 0 25392 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_270
timestamp 1649977179
transform 1 0 25944 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_278
timestamp 1649977179
transform 1 0 26680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_282
timestamp 1649977179
transform 1 0 27048 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_293
timestamp 1649977179
transform 1 0 28060 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1649977179
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1649977179
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_309
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_320
timestamp 1649977179
transform 1 0 30544 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_329
timestamp 1649977179
transform 1 0 31372 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_335
timestamp 1649977179
transform 1 0 31924 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_341
timestamp 1649977179
transform 1 0 32476 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_347
timestamp 1649977179
transform 1 0 33028 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_351
timestamp 1649977179
transform 1 0 33396 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_358
timestamp 1649977179
transform 1 0 34040 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_370
timestamp 1649977179
transform 1 0 35144 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_378
timestamp 1649977179
transform 1 0 35880 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_385
timestamp 1649977179
transform 1 0 36524 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_391
timestamp 1649977179
transform 1 0 37076 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_399
timestamp 1649977179
transform 1 0 37812 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_411
timestamp 1649977179
transform 1 0 38916 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1649977179
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_423
timestamp 1649977179
transform 1 0 40020 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_440
timestamp 1649977179
transform 1 0 41584 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_446
timestamp 1649977179
transform 1 0 42136 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_452
timestamp 1649977179
transform 1 0 42688 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_458
timestamp 1649977179
transform 1 0 43240 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_470
timestamp 1649977179
transform 1 0 44344 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1649977179
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1649977179
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_501
timestamp 1649977179
transform 1 0 47196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_512
timestamp 1649977179
transform 1 0 48208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_3
timestamp 1649977179
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_11
timestamp 1649977179
transform 1 0 2116 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_23
timestamp 1649977179
transform 1 0 3220 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_35
timestamp 1649977179
transform 1 0 4324 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_47
timestamp 1649977179
transform 1 0 5428 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1649977179
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1649977179
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_81
timestamp 1649977179
transform 1 0 8556 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_89
timestamp 1649977179
transform 1 0 9292 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_95
timestamp 1649977179
transform 1 0 9844 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_101
timestamp 1649977179
transform 1 0 10396 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_108
timestamp 1649977179
transform 1 0 11040 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_118
timestamp 1649977179
transform 1 0 11960 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_122
timestamp 1649977179
transform 1 0 12328 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_129
timestamp 1649977179
transform 1 0 12972 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_137
timestamp 1649977179
transform 1 0 13708 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_142
timestamp 1649977179
transform 1 0 14168 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_151
timestamp 1649977179
transform 1 0 14996 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_162
timestamp 1649977179
transform 1 0 16008 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_59_176
timestamp 1649977179
transform 1 0 17296 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_187
timestamp 1649977179
transform 1 0 18308 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_193
timestamp 1649977179
transform 1 0 18860 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_203
timestamp 1649977179
transform 1 0 19780 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_207
timestamp 1649977179
transform 1 0 20148 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_210
timestamp 1649977179
transform 1 0 20424 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_219
timestamp 1649977179
transform 1 0 21252 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1649977179
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_225
timestamp 1649977179
transform 1 0 21804 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_235
timestamp 1649977179
transform 1 0 22724 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_247
timestamp 1649977179
transform 1 0 23828 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_254
timestamp 1649977179
transform 1 0 24472 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_264
timestamp 1649977179
transform 1 0 25392 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_275
timestamp 1649977179
transform 1 0 26404 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1649977179
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_288
timestamp 1649977179
transform 1 0 27600 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_296
timestamp 1649977179
transform 1 0 28336 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_305
timestamp 1649977179
transform 1 0 29164 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_314
timestamp 1649977179
transform 1 0 29992 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_325
timestamp 1649977179
transform 1 0 31004 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_332
timestamp 1649977179
transform 1 0 31648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_339
timestamp 1649977179
transform 1 0 32292 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_345
timestamp 1649977179
transform 1 0 32844 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_349
timestamp 1649977179
transform 1 0 33212 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_355
timestamp 1649977179
transform 1 0 33764 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_363
timestamp 1649977179
transform 1 0 34500 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_371
timestamp 1649977179
transform 1 0 35236 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_379
timestamp 1649977179
transform 1 0 35972 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_387
timestamp 1649977179
transform 1 0 36708 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1649977179
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_399
timestamp 1649977179
transform 1 0 37812 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_409
timestamp 1649977179
transform 1 0 38732 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_416
timestamp 1649977179
transform 1 0 39376 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_422
timestamp 1649977179
transform 1 0 39928 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_439
timestamp 1649977179
transform 1 0 41492 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1649977179
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_451
timestamp 1649977179
transform 1 0 42596 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_457
timestamp 1649977179
transform 1 0 43148 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_469
timestamp 1649977179
transform 1 0 44252 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_481
timestamp 1649977179
transform 1 0 45356 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_493
timestamp 1649977179
transform 1 0 46460 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_501
timestamp 1649977179
transform 1 0 47196 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_505
timestamp 1649977179
transform 1 0 47564 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_513
timestamp 1649977179
transform 1 0 48300 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1649977179
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1649977179
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1649977179
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1649977179
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1649977179
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1649977179
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1649977179
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1649977179
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_97
timestamp 1649977179
transform 1 0 10028 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_100
timestamp 1649977179
transform 1 0 10304 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_106
timestamp 1649977179
transform 1 0 10856 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_112
timestamp 1649977179
transform 1 0 11408 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_119
timestamp 1649977179
transform 1 0 12052 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_123
timestamp 1649977179
transform 1 0 12420 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_128
timestamp 1649977179
transform 1 0 12880 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_136
timestamp 1649977179
transform 1 0 13616 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_147
timestamp 1649977179
transform 1 0 14628 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_151
timestamp 1649977179
transform 1 0 14996 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_158
timestamp 1649977179
transform 1 0 15640 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_167
timestamp 1649977179
transform 1 0 16468 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_173
timestamp 1649977179
transform 1 0 17020 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_182
timestamp 1649977179
transform 1 0 17848 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_192
timestamp 1649977179
transform 1 0 18768 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_199
timestamp 1649977179
transform 1 0 19412 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_207
timestamp 1649977179
transform 1 0 20148 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_218
timestamp 1649977179
transform 1 0 21160 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_226
timestamp 1649977179
transform 1 0 21896 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_230
timestamp 1649977179
transform 1 0 22264 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_241
timestamp 1649977179
transform 1 0 23276 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_245
timestamp 1649977179
transform 1 0 23644 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_248
timestamp 1649977179
transform 1 0 23920 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_253
timestamp 1649977179
transform 1 0 24380 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_257
timestamp 1649977179
transform 1 0 24748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_261
timestamp 1649977179
transform 1 0 25116 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_266
timestamp 1649977179
transform 1 0 25576 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_275
timestamp 1649977179
transform 1 0 26404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_287
timestamp 1649977179
transform 1 0 27508 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_296
timestamp 1649977179
transform 1 0 28336 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_304
timestamp 1649977179
transform 1 0 29072 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_311
timestamp 1649977179
transform 1 0 29716 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_317
timestamp 1649977179
transform 1 0 30268 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_326
timestamp 1649977179
transform 1 0 31096 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_335
timestamp 1649977179
transform 1 0 31924 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_345
timestamp 1649977179
transform 1 0 32844 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_356
timestamp 1649977179
transform 1 0 33856 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_369
timestamp 1649977179
transform 1 0 35052 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_375
timestamp 1649977179
transform 1 0 35604 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_386
timestamp 1649977179
transform 1 0 36616 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_392
timestamp 1649977179
transform 1 0 37168 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_403
timestamp 1649977179
transform 1 0 38180 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_410
timestamp 1649977179
transform 1 0 38824 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_416
timestamp 1649977179
transform 1 0 39376 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_428
timestamp 1649977179
transform 1 0 40480 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_434
timestamp 1649977179
transform 1 0 41032 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_440
timestamp 1649977179
transform 1 0 41584 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_446
timestamp 1649977179
transform 1 0 42136 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_452
timestamp 1649977179
transform 1 0 42688 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_458
timestamp 1649977179
transform 1 0 43240 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_470
timestamp 1649977179
transform 1 0 44344 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1649977179
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1649977179
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1649977179
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_513
timestamp 1649977179
transform 1 0 48300 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1649977179
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1649977179
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1649977179
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1649977179
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1649977179
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1649977179
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1649977179
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1649977179
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1649977179
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_93
timestamp 1649977179
transform 1 0 9660 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_99
timestamp 1649977179
transform 1 0 10212 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_102
timestamp 1649977179
transform 1 0 10488 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_108
timestamp 1649977179
transform 1 0 11040 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_115
timestamp 1649977179
transform 1 0 11684 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_121
timestamp 1649977179
transform 1 0 12236 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_127
timestamp 1649977179
transform 1 0 12788 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_133
timestamp 1649977179
transform 1 0 13340 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_139
timestamp 1649977179
transform 1 0 13892 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_146
timestamp 1649977179
transform 1 0 14536 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_152
timestamp 1649977179
transform 1 0 15088 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_160
timestamp 1649977179
transform 1 0 15824 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_61_174
timestamp 1649977179
transform 1 0 17112 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_186
timestamp 1649977179
transform 1 0 18216 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_198
timestamp 1649977179
transform 1 0 19320 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_205
timestamp 1649977179
transform 1 0 19964 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1649977179
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1649977179
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_225
timestamp 1649977179
transform 1 0 21804 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_235
timestamp 1649977179
transform 1 0 22724 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_241
timestamp 1649977179
transform 1 0 23276 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_244
timestamp 1649977179
transform 1 0 23552 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_250
timestamp 1649977179
transform 1 0 24104 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_262
timestamp 1649977179
transform 1 0 25208 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1649977179
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1649977179
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_285
timestamp 1649977179
transform 1 0 27324 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_291
timestamp 1649977179
transform 1 0 27876 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_297
timestamp 1649977179
transform 1 0 28428 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_61_311
timestamp 1649977179
transform 1 0 29716 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_317
timestamp 1649977179
transform 1 0 30268 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_327
timestamp 1649977179
transform 1 0 31188 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1649977179
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_342
timestamp 1649977179
transform 1 0 32568 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_348
timestamp 1649977179
transform 1 0 33120 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_354
timestamp 1649977179
transform 1 0 33672 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_362
timestamp 1649977179
transform 1 0 34408 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_368
timestamp 1649977179
transform 1 0 34960 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_372
timestamp 1649977179
transform 1 0 35328 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_376
timestamp 1649977179
transform 1 0 35696 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_383
timestamp 1649977179
transform 1 0 36340 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1649977179
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_396
timestamp 1649977179
transform 1 0 37536 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_407
timestamp 1649977179
transform 1 0 38548 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_415
timestamp 1649977179
transform 1 0 39284 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_421
timestamp 1649977179
transform 1 0 39836 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_427
timestamp 1649977179
transform 1 0 40388 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_433
timestamp 1649977179
transform 1 0 40940 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_439
timestamp 1649977179
transform 1 0 41492 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1649977179
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_451
timestamp 1649977179
transform 1 0 42596 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_457
timestamp 1649977179
transform 1 0 43148 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_463
timestamp 1649977179
transform 1 0 43700 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_475
timestamp 1649977179
transform 1 0 44804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_487
timestamp 1649977179
transform 1 0 45908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_499
timestamp 1649977179
transform 1 0 47012 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1649977179
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_505
timestamp 1649977179
transform 1 0 47564 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_509
timestamp 1649977179
transform 1 0 47932 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_512
timestamp 1649977179
transform 1 0 48208 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_7
timestamp 1649977179
transform 1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_13
timestamp 1649977179
transform 1 0 2300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_25
timestamp 1649977179
transform 1 0 3404 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1649977179
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1649977179
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1649977179
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1649977179
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1649977179
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1649977179
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_109
timestamp 1649977179
transform 1 0 11132 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_112
timestamp 1649977179
transform 1 0 11408 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_118
timestamp 1649977179
transform 1 0 11960 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_124
timestamp 1649977179
transform 1 0 12512 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_130
timestamp 1649977179
transform 1 0 13064 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_136
timestamp 1649977179
transform 1 0 13616 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_141
timestamp 1649977179
transform 1 0 14076 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_146
timestamp 1649977179
transform 1 0 14536 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_152
timestamp 1649977179
transform 1 0 15088 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_163
timestamp 1649977179
transform 1 0 16100 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_170
timestamp 1649977179
transform 1 0 16744 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_174
timestamp 1649977179
transform 1 0 17112 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_181
timestamp 1649977179
transform 1 0 17756 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_185
timestamp 1649977179
transform 1 0 18124 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_191
timestamp 1649977179
transform 1 0 18676 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1649977179
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_200
timestamp 1649977179
transform 1 0 19504 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_206
timestamp 1649977179
transform 1 0 20056 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_213
timestamp 1649977179
transform 1 0 20700 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_223
timestamp 1649977179
transform 1 0 21620 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_229
timestamp 1649977179
transform 1 0 22172 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_240
timestamp 1649977179
transform 1 0 23184 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_248
timestamp 1649977179
transform 1 0 23920 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_253
timestamp 1649977179
transform 1 0 24380 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_256
timestamp 1649977179
transform 1 0 24656 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_264
timestamp 1649977179
transform 1 0 25392 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_271
timestamp 1649977179
transform 1 0 26036 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_277
timestamp 1649977179
transform 1 0 26588 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_283
timestamp 1649977179
transform 1 0 27140 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_292
timestamp 1649977179
transform 1 0 27968 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_303
timestamp 1649977179
transform 1 0 28980 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1649977179
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_309
timestamp 1649977179
transform 1 0 29532 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_313
timestamp 1649977179
transform 1 0 29900 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_323
timestamp 1649977179
transform 1 0 30820 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_336
timestamp 1649977179
transform 1 0 32016 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_344
timestamp 1649977179
transform 1 0 32752 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_350
timestamp 1649977179
transform 1 0 33304 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1649977179
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1649977179
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_367
timestamp 1649977179
transform 1 0 34868 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_376
timestamp 1649977179
transform 1 0 35696 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_384
timestamp 1649977179
transform 1 0 36432 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_393
timestamp 1649977179
transform 1 0 37260 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_407
timestamp 1649977179
transform 1 0 38548 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_414
timestamp 1649977179
transform 1 0 39192 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_429
timestamp 1649977179
transform 1 0 40572 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_439
timestamp 1649977179
transform 1 0 41492 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_445
timestamp 1649977179
transform 1 0 42044 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_451
timestamp 1649977179
transform 1 0 42596 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1649977179
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1649977179
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1649977179
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1649977179
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_489
timestamp 1649977179
transform 1 0 46092 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_497
timestamp 1649977179
transform 1 0 46828 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_502
timestamp 1649977179
transform 1 0 47288 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_512
timestamp 1649977179
transform 1 0 48208 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1649977179
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1649977179
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1649977179
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1649977179
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1649977179
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1649977179
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1649977179
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1649977179
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1649977179
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1649977179
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_105
timestamp 1649977179
transform 1 0 10764 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_108
timestamp 1649977179
transform 1 0 11040 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_113
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_118
timestamp 1649977179
transform 1 0 11960 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_124
timestamp 1649977179
transform 1 0 12512 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_130
timestamp 1649977179
transform 1 0 13064 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_137
timestamp 1649977179
transform 1 0 13708 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_144
timestamp 1649977179
transform 1 0 14352 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_63_156
timestamp 1649977179
transform 1 0 15456 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_164
timestamp 1649977179
transform 1 0 16192 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1649977179
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_173
timestamp 1649977179
transform 1 0 17020 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_183
timestamp 1649977179
transform 1 0 17940 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_196
timestamp 1649977179
transform 1 0 19136 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_205
timestamp 1649977179
transform 1 0 19964 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_214
timestamp 1649977179
transform 1 0 20792 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_220
timestamp 1649977179
transform 1 0 21344 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_225
timestamp 1649977179
transform 1 0 21804 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_229
timestamp 1649977179
transform 1 0 22172 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_238
timestamp 1649977179
transform 1 0 23000 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_246
timestamp 1649977179
transform 1 0 23736 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_255
timestamp 1649977179
transform 1 0 24564 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_266
timestamp 1649977179
transform 1 0 25576 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_272
timestamp 1649977179
transform 1 0 26128 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_281
timestamp 1649977179
transform 1 0 26956 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_291
timestamp 1649977179
transform 1 0 27876 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_303
timestamp 1649977179
transform 1 0 28980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_313
timestamp 1649977179
transform 1 0 29900 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_317
timestamp 1649977179
transform 1 0 30268 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_321
timestamp 1649977179
transform 1 0 30636 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_330
timestamp 1649977179
transform 1 0 31464 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_337
timestamp 1649977179
transform 1 0 32108 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_349
timestamp 1649977179
transform 1 0 33212 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_358
timestamp 1649977179
transform 1 0 34040 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_367
timestamp 1649977179
transform 1 0 34868 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_373
timestamp 1649977179
transform 1 0 35420 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_381
timestamp 1649977179
transform 1 0 36156 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_388
timestamp 1649977179
transform 1 0 36800 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_395
timestamp 1649977179
transform 1 0 37444 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_399
timestamp 1649977179
transform 1 0 37812 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_406
timestamp 1649977179
transform 1 0 38456 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_412
timestamp 1649977179
transform 1 0 39008 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_416
timestamp 1649977179
transform 1 0 39376 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_426
timestamp 1649977179
transform 1 0 40296 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_430
timestamp 1649977179
transform 1 0 40664 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_444
timestamp 1649977179
transform 1 0 41952 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_451
timestamp 1649977179
transform 1 0 42596 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_457
timestamp 1649977179
transform 1 0 43148 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_469
timestamp 1649977179
transform 1 0 44252 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_481
timestamp 1649977179
transform 1 0 45356 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_493
timestamp 1649977179
transform 1 0 46460 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_500
timestamp 1649977179
transform 1 0 47104 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_510
timestamp 1649977179
transform 1 0 48024 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1649977179
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1649977179
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1649977179
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1649977179
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1649977179
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1649977179
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1649977179
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1649977179
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_97
timestamp 1649977179
transform 1 0 10028 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_102
timestamp 1649977179
transform 1 0 10488 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_108
timestamp 1649977179
transform 1 0 11040 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_114
timestamp 1649977179
transform 1 0 11592 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_120
timestamp 1649977179
transform 1 0 12144 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_127
timestamp 1649977179
transform 1 0 12788 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_136
timestamp 1649977179
transform 1 0 13616 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_141
timestamp 1649977179
transform 1 0 14076 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_145
timestamp 1649977179
transform 1 0 14444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_154
timestamp 1649977179
transform 1 0 15272 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_163
timestamp 1649977179
transform 1 0 16100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_169
timestamp 1649977179
transform 1 0 16652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_172
timestamp 1649977179
transform 1 0 16928 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_179
timestamp 1649977179
transform 1 0 17572 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_183
timestamp 1649977179
transform 1 0 17940 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_186
timestamp 1649977179
transform 1 0 18216 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_192
timestamp 1649977179
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1649977179
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_204
timestamp 1649977179
transform 1 0 19872 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_216
timestamp 1649977179
transform 1 0 20976 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_227
timestamp 1649977179
transform 1 0 21988 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_235
timestamp 1649977179
transform 1 0 22724 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_241
timestamp 1649977179
transform 1 0 23276 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_248
timestamp 1649977179
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_260
timestamp 1649977179
transform 1 0 25024 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_268
timestamp 1649977179
transform 1 0 25760 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_274
timestamp 1649977179
transform 1 0 26312 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_287
timestamp 1649977179
transform 1 0 27508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_293
timestamp 1649977179
transform 1 0 28060 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_300
timestamp 1649977179
transform 1 0 28704 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_309
timestamp 1649977179
transform 1 0 29532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_321
timestamp 1649977179
transform 1 0 30636 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_330
timestamp 1649977179
transform 1 0 31464 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_339
timestamp 1649977179
transform 1 0 32292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_348
timestamp 1649977179
transform 1 0 33120 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_360
timestamp 1649977179
transform 1 0 34224 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_368
timestamp 1649977179
transform 1 0 34960 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_374
timestamp 1649977179
transform 1 0 35512 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_380
timestamp 1649977179
transform 1 0 36064 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_389
timestamp 1649977179
transform 1 0 36892 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_395
timestamp 1649977179
transform 1 0 37444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_401
timestamp 1649977179
transform 1 0 37996 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_407
timestamp 1649977179
transform 1 0 38548 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_416
timestamp 1649977179
transform 1 0 39376 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_424
timestamp 1649977179
transform 1 0 40112 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_436
timestamp 1649977179
transform 1 0 41216 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_442
timestamp 1649977179
transform 1 0 41768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_448
timestamp 1649977179
transform 1 0 42320 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_454
timestamp 1649977179
transform 1 0 42872 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_460
timestamp 1649977179
transform 1 0 43424 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_472
timestamp 1649977179
transform 1 0 44528 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1649977179
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1649977179
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_501
timestamp 1649977179
transform 1 0 47196 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_509
timestamp 1649977179
transform 1 0 47932 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_512
timestamp 1649977179
transform 1 0 48208 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_3
timestamp 1649977179
transform 1 0 1380 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_7
timestamp 1649977179
transform 1 0 1748 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_19
timestamp 1649977179
transform 1 0 2852 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_31
timestamp 1649977179
transform 1 0 3956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_43
timestamp 1649977179
transform 1 0 5060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1649977179
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1649977179
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1649977179
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1649977179
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1649977179
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_105
timestamp 1649977179
transform 1 0 10764 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_108
timestamp 1649977179
transform 1 0 11040 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_113
timestamp 1649977179
transform 1 0 11500 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_117
timestamp 1649977179
transform 1 0 11868 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_123
timestamp 1649977179
transform 1 0 12420 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_129
timestamp 1649977179
transform 1 0 12972 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_135
timestamp 1649977179
transform 1 0 13524 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_147
timestamp 1649977179
transform 1 0 14628 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_157
timestamp 1649977179
transform 1 0 15548 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_161
timestamp 1649977179
transform 1 0 15916 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_164
timestamp 1649977179
transform 1 0 16192 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_173
timestamp 1649977179
transform 1 0 17020 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_179
timestamp 1649977179
transform 1 0 17572 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_187
timestamp 1649977179
transform 1 0 18308 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_195
timestamp 1649977179
transform 1 0 19044 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_205
timestamp 1649977179
transform 1 0 19964 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_215
timestamp 1649977179
transform 1 0 20884 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1649977179
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_231
timestamp 1649977179
transform 1 0 22356 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_239
timestamp 1649977179
transform 1 0 23092 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_247
timestamp 1649977179
transform 1 0 23828 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_259
timestamp 1649977179
transform 1 0 24932 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_265
timestamp 1649977179
transform 1 0 25484 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_276
timestamp 1649977179
transform 1 0 26496 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_288
timestamp 1649977179
transform 1 0 27600 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_299
timestamp 1649977179
transform 1 0 28612 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_311
timestamp 1649977179
transform 1 0 29716 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_320
timestamp 1649977179
transform 1 0 30544 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_327
timestamp 1649977179
transform 1 0 31188 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1649977179
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_345
timestamp 1649977179
transform 1 0 32844 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_65_358
timestamp 1649977179
transform 1 0 34040 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_366
timestamp 1649977179
transform 1 0 34776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_372
timestamp 1649977179
transform 1 0 35328 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_378
timestamp 1649977179
transform 1 0 35880 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1649977179
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1649977179
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_396
timestamp 1649977179
transform 1 0 37536 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_402
timestamp 1649977179
transform 1 0 38088 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_410
timestamp 1649977179
transform 1 0 38824 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_416
timestamp 1649977179
transform 1 0 39376 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_431
timestamp 1649977179
transform 1 0 40756 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_437
timestamp 1649977179
transform 1 0 41308 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_443
timestamp 1649977179
transform 1 0 41860 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1649977179
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_451
timestamp 1649977179
transform 1 0 42596 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_463
timestamp 1649977179
transform 1 0 43700 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_475
timestamp 1649977179
transform 1 0 44804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_487
timestamp 1649977179
transform 1 0 45908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_499
timestamp 1649977179
transform 1 0 47012 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1649977179
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_505
timestamp 1649977179
transform 1 0 47564 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_513
timestamp 1649977179
transform 1 0 48300 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_3
timestamp 1649977179
transform 1 0 1380 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_11
timestamp 1649977179
transform 1 0 2116 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_23
timestamp 1649977179
transform 1 0 3220 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1649977179
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1649977179
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1649977179
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1649977179
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1649977179
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1649977179
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1649977179
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1649977179
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1649977179
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_109
timestamp 1649977179
transform 1 0 11132 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_112
timestamp 1649977179
transform 1 0 11408 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_118
timestamp 1649977179
transform 1 0 11960 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_124
timestamp 1649977179
transform 1 0 12512 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_130
timestamp 1649977179
transform 1 0 13064 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_136
timestamp 1649977179
transform 1 0 13616 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_141
timestamp 1649977179
transform 1 0 14076 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_144
timestamp 1649977179
transform 1 0 14352 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_154
timestamp 1649977179
transform 1 0 15272 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_164
timestamp 1649977179
transform 1 0 16192 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_174
timestamp 1649977179
transform 1 0 17112 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_178
timestamp 1649977179
transform 1 0 17480 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_182
timestamp 1649977179
transform 1 0 17848 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_191
timestamp 1649977179
transform 1 0 18676 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1649977179
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_199
timestamp 1649977179
transform 1 0 19412 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_206
timestamp 1649977179
transform 1 0 20056 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_213
timestamp 1649977179
transform 1 0 20700 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_219
timestamp 1649977179
transform 1 0 21252 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_222
timestamp 1649977179
transform 1 0 21528 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_232
timestamp 1649977179
transform 1 0 22448 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_236
timestamp 1649977179
transform 1 0 22816 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_242
timestamp 1649977179
transform 1 0 23368 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_248
timestamp 1649977179
transform 1 0 23920 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_262
timestamp 1649977179
transform 1 0 25208 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_268
timestamp 1649977179
transform 1 0 25760 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_272
timestamp 1649977179
transform 1 0 26128 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_280
timestamp 1649977179
transform 1 0 26864 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_293
timestamp 1649977179
transform 1 0 28060 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_299
timestamp 1649977179
transform 1 0 28612 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_304
timestamp 1649977179
transform 1 0 29072 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_316
timestamp 1649977179
transform 1 0 30176 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_324
timestamp 1649977179
transform 1 0 30912 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_332
timestamp 1649977179
transform 1 0 31648 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_340
timestamp 1649977179
transform 1 0 32384 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_348
timestamp 1649977179
transform 1 0 33120 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_356
timestamp 1649977179
transform 1 0 33856 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_372
timestamp 1649977179
transform 1 0 35328 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_383
timestamp 1649977179
transform 1 0 36340 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_394
timestamp 1649977179
transform 1 0 37352 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_405
timestamp 1649977179
transform 1 0 38364 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_412
timestamp 1649977179
transform 1 0 39008 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_423
timestamp 1649977179
transform 1 0 40020 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_429
timestamp 1649977179
transform 1 0 40572 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_435
timestamp 1649977179
transform 1 0 41124 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_441
timestamp 1649977179
transform 1 0 41676 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_447
timestamp 1649977179
transform 1 0 42228 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_453
timestamp 1649977179
transform 1 0 42780 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_459
timestamp 1649977179
transform 1 0 43332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_471
timestamp 1649977179
transform 1 0 44436 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1649977179
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1649977179
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1649977179
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_501
timestamp 1649977179
transform 1 0 47196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_504
timestamp 1649977179
transform 1 0 47472 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_512
timestamp 1649977179
transform 1 0 48208 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1649977179
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1649977179
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1649977179
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1649977179
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1649977179
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1649977179
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1649977179
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1649977179
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1649977179
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1649977179
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_105
timestamp 1649977179
transform 1 0 10764 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_108
timestamp 1649977179
transform 1 0 11040 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_113
timestamp 1649977179
transform 1 0 11500 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_117
timestamp 1649977179
transform 1 0 11868 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_123
timestamp 1649977179
transform 1 0 12420 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_129
timestamp 1649977179
transform 1 0 12972 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_136
timestamp 1649977179
transform 1 0 13616 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_142
timestamp 1649977179
transform 1 0 14168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_147
timestamp 1649977179
transform 1 0 14628 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_151
timestamp 1649977179
transform 1 0 14996 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_155
timestamp 1649977179
transform 1 0 15364 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_164
timestamp 1649977179
transform 1 0 16192 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_174
timestamp 1649977179
transform 1 0 17112 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_180
timestamp 1649977179
transform 1 0 17664 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_183
timestamp 1649977179
transform 1 0 17940 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_193
timestamp 1649977179
transform 1 0 18860 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_202
timestamp 1649977179
transform 1 0 19688 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_211
timestamp 1649977179
transform 1 0 20516 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_218
timestamp 1649977179
transform 1 0 21160 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_230
timestamp 1649977179
transform 1 0 22264 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_234
timestamp 1649977179
transform 1 0 22632 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_239
timestamp 1649977179
transform 1 0 23092 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_243
timestamp 1649977179
transform 1 0 23460 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_248
timestamp 1649977179
transform 1 0 23920 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_259
timestamp 1649977179
transform 1 0 24932 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_267
timestamp 1649977179
transform 1 0 25668 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_273
timestamp 1649977179
transform 1 0 26220 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_276
timestamp 1649977179
transform 1 0 26496 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_281
timestamp 1649977179
transform 1 0 26956 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_287
timestamp 1649977179
transform 1 0 27508 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_295
timestamp 1649977179
transform 1 0 28244 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_303
timestamp 1649977179
transform 1 0 28980 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_314
timestamp 1649977179
transform 1 0 29992 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_320
timestamp 1649977179
transform 1 0 30544 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_330
timestamp 1649977179
transform 1 0 31464 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_337
timestamp 1649977179
transform 1 0 32108 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_347
timestamp 1649977179
transform 1 0 33028 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_357
timestamp 1649977179
transform 1 0 33948 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_365
timestamp 1649977179
transform 1 0 34684 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_371
timestamp 1649977179
transform 1 0 35236 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_377
timestamp 1649977179
transform 1 0 35788 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_384
timestamp 1649977179
transform 1 0 36432 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_393
timestamp 1649977179
transform 1 0 37260 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_399
timestamp 1649977179
transform 1 0 37812 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_408
timestamp 1649977179
transform 1 0 38640 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_417
timestamp 1649977179
transform 1 0 39468 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_426
timestamp 1649977179
transform 1 0 40296 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_432
timestamp 1649977179
transform 1 0 40848 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_438
timestamp 1649977179
transform 1 0 41400 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_444
timestamp 1649977179
transform 1 0 41952 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_451
timestamp 1649977179
transform 1 0 42596 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_457
timestamp 1649977179
transform 1 0 43148 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_463
timestamp 1649977179
transform 1 0 43700 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_475
timestamp 1649977179
transform 1 0 44804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_487
timestamp 1649977179
transform 1 0 45908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_499
timestamp 1649977179
transform 1 0 47012 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1649977179
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_505
timestamp 1649977179
transform 1 0 47564 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_513
timestamp 1649977179
transform 1 0 48300 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1649977179
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1649977179
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1649977179
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1649977179
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1649977179
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1649977179
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1649977179
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1649977179
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1649977179
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1649977179
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1649977179
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_111
timestamp 1649977179
transform 1 0 11316 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_117
timestamp 1649977179
transform 1 0 11868 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_123
timestamp 1649977179
transform 1 0 12420 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_129
timestamp 1649977179
transform 1 0 12972 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_136
timestamp 1649977179
transform 1 0 13616 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_146
timestamp 1649977179
transform 1 0 14536 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_150
timestamp 1649977179
transform 1 0 14904 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_158
timestamp 1649977179
transform 1 0 15640 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_68_167
timestamp 1649977179
transform 1 0 16468 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_177
timestamp 1649977179
transform 1 0 17388 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_188
timestamp 1649977179
transform 1 0 18400 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_199
timestamp 1649977179
transform 1 0 19412 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_205
timestamp 1649977179
transform 1 0 19964 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_216
timestamp 1649977179
transform 1 0 20976 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_224
timestamp 1649977179
transform 1 0 21712 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_231
timestamp 1649977179
transform 1 0 22356 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_239
timestamp 1649977179
transform 1 0 23092 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_248
timestamp 1649977179
transform 1 0 23920 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_253
timestamp 1649977179
transform 1 0 24380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_261
timestamp 1649977179
transform 1 0 25116 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_269
timestamp 1649977179
transform 1 0 25852 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_279
timestamp 1649977179
transform 1 0 26772 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_287
timestamp 1649977179
transform 1 0 27508 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_291
timestamp 1649977179
transform 1 0 27876 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_295
timestamp 1649977179
transform 1 0 28244 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_302
timestamp 1649977179
transform 1 0 28888 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_309
timestamp 1649977179
transform 1 0 29532 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_316
timestamp 1649977179
transform 1 0 30176 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_322
timestamp 1649977179
transform 1 0 30728 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_336
timestamp 1649977179
transform 1 0 32016 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_351
timestamp 1649977179
transform 1 0 33396 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_360
timestamp 1649977179
transform 1 0 34224 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_373
timestamp 1649977179
transform 1 0 35420 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_381
timestamp 1649977179
transform 1 0 36156 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_387
timestamp 1649977179
transform 1 0 36708 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_393
timestamp 1649977179
transform 1 0 37260 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_401
timestamp 1649977179
transform 1 0 37996 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_405
timestamp 1649977179
transform 1 0 38364 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_414
timestamp 1649977179
transform 1 0 39192 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_424
timestamp 1649977179
transform 1 0 40112 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_430
timestamp 1649977179
transform 1 0 40664 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_436
timestamp 1649977179
transform 1 0 41216 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_442
timestamp 1649977179
transform 1 0 41768 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_448
timestamp 1649977179
transform 1 0 42320 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_454
timestamp 1649977179
transform 1 0 42872 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_460
timestamp 1649977179
transform 1 0 43424 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_466
timestamp 1649977179
transform 1 0 43976 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_474
timestamp 1649977179
transform 1 0 44712 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1649977179
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1649977179
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1649977179
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_513
timestamp 1649977179
transform 1 0 48300 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_3
timestamp 1649977179
transform 1 0 1380 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_7
timestamp 1649977179
transform 1 0 1748 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_19
timestamp 1649977179
transform 1 0 2852 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_31
timestamp 1649977179
transform 1 0 3956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_43
timestamp 1649977179
transform 1 0 5060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1649977179
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1649977179
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1649977179
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1649977179
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1649977179
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1649977179
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1649977179
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_113
timestamp 1649977179
transform 1 0 11500 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_121
timestamp 1649977179
transform 1 0 12236 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_127
timestamp 1649977179
transform 1 0 12788 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_133
timestamp 1649977179
transform 1 0 13340 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_139
timestamp 1649977179
transform 1 0 13892 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_150
timestamp 1649977179
transform 1 0 14904 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_158
timestamp 1649977179
transform 1 0 15640 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_164
timestamp 1649977179
transform 1 0 16192 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_169
timestamp 1649977179
transform 1 0 16652 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_173
timestamp 1649977179
transform 1 0 17020 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_181
timestamp 1649977179
transform 1 0 17756 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_187
timestamp 1649977179
transform 1 0 18308 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_190
timestamp 1649977179
transform 1 0 18584 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_199
timestamp 1649977179
transform 1 0 19412 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_207
timestamp 1649977179
transform 1 0 20148 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_212
timestamp 1649977179
transform 1 0 20608 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_219
timestamp 1649977179
transform 1 0 21252 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1649977179
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_232
timestamp 1649977179
transform 1 0 22448 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_244
timestamp 1649977179
transform 1 0 23552 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_255
timestamp 1649977179
transform 1 0 24564 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_261
timestamp 1649977179
transform 1 0 25116 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_270
timestamp 1649977179
transform 1 0 25944 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_276
timestamp 1649977179
transform 1 0 26496 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_285
timestamp 1649977179
transform 1 0 27324 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_292
timestamp 1649977179
transform 1 0 27968 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_298
timestamp 1649977179
transform 1 0 28520 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_304
timestamp 1649977179
transform 1 0 29072 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_308
timestamp 1649977179
transform 1 0 29440 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_314
timestamp 1649977179
transform 1 0 29992 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_318
timestamp 1649977179
transform 1 0 30360 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_324
timestamp 1649977179
transform 1 0 30912 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_330
timestamp 1649977179
transform 1 0 31464 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_337
timestamp 1649977179
transform 1 0 32108 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_347
timestamp 1649977179
transform 1 0 33028 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_354
timestamp 1649977179
transform 1 0 33672 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_367
timestamp 1649977179
transform 1 0 34868 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_373
timestamp 1649977179
transform 1 0 35420 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_381
timestamp 1649977179
transform 1 0 36156 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_388
timestamp 1649977179
transform 1 0 36800 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_400
timestamp 1649977179
transform 1 0 37904 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_406
timestamp 1649977179
transform 1 0 38456 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_411
timestamp 1649977179
transform 1 0 38916 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_418
timestamp 1649977179
transform 1 0 39560 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_424
timestamp 1649977179
transform 1 0 40112 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_430
timestamp 1649977179
transform 1 0 40664 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_436
timestamp 1649977179
transform 1 0 41216 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_442
timestamp 1649977179
transform 1 0 41768 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_451
timestamp 1649977179
transform 1 0 42596 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_457
timestamp 1649977179
transform 1 0 43148 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_469
timestamp 1649977179
transform 1 0 44252 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_481
timestamp 1649977179
transform 1 0 45356 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_493
timestamp 1649977179
transform 1 0 46460 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_501
timestamp 1649977179
transform 1 0 47196 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_505
timestamp 1649977179
transform 1 0 47564 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_513
timestamp 1649977179
transform 1 0 48300 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_3
timestamp 1649977179
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_11
timestamp 1649977179
transform 1 0 2116 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_23
timestamp 1649977179
transform 1 0 3220 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1649977179
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1649977179
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1649977179
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1649977179
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1649977179
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1649977179
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1649977179
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1649977179
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1649977179
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_109
timestamp 1649977179
transform 1 0 11132 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_115
timestamp 1649977179
transform 1 0 11684 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_118
timestamp 1649977179
transform 1 0 11960 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_124
timestamp 1649977179
transform 1 0 12512 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_130
timestamp 1649977179
transform 1 0 13064 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_136
timestamp 1649977179
transform 1 0 13616 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_141
timestamp 1649977179
transform 1 0 14076 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_147
timestamp 1649977179
transform 1 0 14628 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_155
timestamp 1649977179
transform 1 0 15364 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_162
timestamp 1649977179
transform 1 0 16008 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_168
timestamp 1649977179
transform 1 0 16560 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_174
timestamp 1649977179
transform 1 0 17112 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_180
timestamp 1649977179
transform 1 0 17664 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_192
timestamp 1649977179
transform 1 0 18768 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_204
timestamp 1649977179
transform 1 0 19872 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_213
timestamp 1649977179
transform 1 0 20700 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_220
timestamp 1649977179
transform 1 0 21344 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_231
timestamp 1649977179
transform 1 0 22356 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_239
timestamp 1649977179
transform 1 0 23092 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_243
timestamp 1649977179
transform 1 0 23460 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_248
timestamp 1649977179
transform 1 0 23920 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_253
timestamp 1649977179
transform 1 0 24380 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_262
timestamp 1649977179
transform 1 0 25208 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_271
timestamp 1649977179
transform 1 0 26036 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_279
timestamp 1649977179
transform 1 0 26772 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_304
timestamp 1649977179
transform 1 0 29072 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_326
timestamp 1649977179
transform 1 0 31096 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_330
timestamp 1649977179
transform 1 0 31464 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_334
timestamp 1649977179
transform 1 0 31832 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_343
timestamp 1649977179
transform 1 0 32660 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_352
timestamp 1649977179
transform 1 0 33488 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_360
timestamp 1649977179
transform 1 0 34224 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_370
timestamp 1649977179
transform 1 0 35144 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_378
timestamp 1649977179
transform 1 0 35880 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_385
timestamp 1649977179
transform 1 0 36524 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_394
timestamp 1649977179
transform 1 0 37352 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_403
timestamp 1649977179
transform 1 0 38180 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_409
timestamp 1649977179
transform 1 0 38732 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_415
timestamp 1649977179
transform 1 0 39284 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1649977179
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_423
timestamp 1649977179
transform 1 0 40020 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_429
timestamp 1649977179
transform 1 0 40572 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_435
timestamp 1649977179
transform 1 0 41124 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_441
timestamp 1649977179
transform 1 0 41676 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_447
timestamp 1649977179
transform 1 0 42228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_459
timestamp 1649977179
transform 1 0 43332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_471
timestamp 1649977179
transform 1 0 44436 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1649977179
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1649977179
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1649977179
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_501
timestamp 1649977179
transform 1 0 47196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_504
timestamp 1649977179
transform 1 0 47472 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_512
timestamp 1649977179
transform 1 0 48208 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1649977179
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1649977179
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1649977179
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1649977179
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1649977179
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1649977179
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1649977179
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1649977179
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1649977179
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1649977179
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_105
timestamp 1649977179
transform 1 0 10764 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_108
timestamp 1649977179
transform 1 0 11040 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_113
timestamp 1649977179
transform 1 0 11500 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_119
timestamp 1649977179
transform 1 0 12052 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_125
timestamp 1649977179
transform 1 0 12604 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_131
timestamp 1649977179
transform 1 0 13156 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_137
timestamp 1649977179
transform 1 0 13708 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_144
timestamp 1649977179
transform 1 0 14352 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_153
timestamp 1649977179
transform 1 0 15180 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_164
timestamp 1649977179
transform 1 0 16192 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_176
timestamp 1649977179
transform 1 0 17296 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_183
timestamp 1649977179
transform 1 0 17940 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_187
timestamp 1649977179
transform 1 0 18308 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_192
timestamp 1649977179
transform 1 0 18768 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_204
timestamp 1649977179
transform 1 0 19872 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_211
timestamp 1649977179
transform 1 0 20516 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_217
timestamp 1649977179
transform 1 0 21068 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_220
timestamp 1649977179
transform 1 0 21344 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_230
timestamp 1649977179
transform 1 0 22264 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_237
timestamp 1649977179
transform 1 0 22908 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_243
timestamp 1649977179
transform 1 0 23460 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_249
timestamp 1649977179
transform 1 0 24012 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_257
timestamp 1649977179
transform 1 0 24748 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_263
timestamp 1649977179
transform 1 0 25300 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_268
timestamp 1649977179
transform 1 0 25760 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_274
timestamp 1649977179
transform 1 0 26312 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_71_283
timestamp 1649977179
transform 1 0 27140 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_71_291
timestamp 1649977179
transform 1 0 27876 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_319
timestamp 1649977179
transform 1 0 30452 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_325
timestamp 1649977179
transform 1 0 31004 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_331
timestamp 1649977179
transform 1 0 31556 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1649977179
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_354
timestamp 1649977179
transform 1 0 33672 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_362
timestamp 1649977179
transform 1 0 34408 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_369
timestamp 1649977179
transform 1 0 35052 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_375
timestamp 1649977179
transform 1 0 35604 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_380
timestamp 1649977179
transform 1 0 36064 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_387
timestamp 1649977179
transform 1 0 36708 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1649977179
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_395
timestamp 1649977179
transform 1 0 37444 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_403
timestamp 1649977179
transform 1 0 38180 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_409
timestamp 1649977179
transform 1 0 38732 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_415
timestamp 1649977179
transform 1 0 39284 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_421
timestamp 1649977179
transform 1 0 39836 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_427
timestamp 1649977179
transform 1 0 40388 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_433
timestamp 1649977179
transform 1 0 40940 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_439
timestamp 1649977179
transform 1 0 41492 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1649977179
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1649977179
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1649977179
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1649977179
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1649977179
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1649977179
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1649977179
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_505
timestamp 1649977179
transform 1 0 47564 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_513
timestamp 1649977179
transform 1 0 48300 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1649977179
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1649977179
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1649977179
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1649977179
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1649977179
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1649977179
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1649977179
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1649977179
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1649977179
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1649977179
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1649977179
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_109
timestamp 1649977179
transform 1 0 11132 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_112
timestamp 1649977179
transform 1 0 11408 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_118
timestamp 1649977179
transform 1 0 11960 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_124
timestamp 1649977179
transform 1 0 12512 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_130
timestamp 1649977179
transform 1 0 13064 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_136
timestamp 1649977179
transform 1 0 13616 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_141
timestamp 1649977179
transform 1 0 14076 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_144
timestamp 1649977179
transform 1 0 14352 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_152
timestamp 1649977179
transform 1 0 15088 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_162
timestamp 1649977179
transform 1 0 16008 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_72_178
timestamp 1649977179
transform 1 0 17480 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_186
timestamp 1649977179
transform 1 0 18216 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_190
timestamp 1649977179
transform 1 0 18584 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_197
timestamp 1649977179
transform 1 0 19228 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_204
timestamp 1649977179
transform 1 0 19872 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_212
timestamp 1649977179
transform 1 0 20608 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_215
timestamp 1649977179
transform 1 0 20884 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_221
timestamp 1649977179
transform 1 0 21436 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_229
timestamp 1649977179
transform 1 0 22172 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_233
timestamp 1649977179
transform 1 0 22540 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_236
timestamp 1649977179
transform 1 0 22816 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_242
timestamp 1649977179
transform 1 0 23368 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_248
timestamp 1649977179
transform 1 0 23920 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_256
timestamp 1649977179
transform 1 0 24656 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_264
timestamp 1649977179
transform 1 0 25392 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_267
timestamp 1649977179
transform 1 0 25668 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_291
timestamp 1649977179
transform 1 0 27876 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_297
timestamp 1649977179
transform 1 0 28428 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_303
timestamp 1649977179
transform 1 0 28980 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1649977179
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_328
timestamp 1649977179
transform 1 0 31280 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_334
timestamp 1649977179
transform 1 0 31832 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_72_343
timestamp 1649977179
transform 1 0 32660 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_349
timestamp 1649977179
transform 1 0 33212 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_359
timestamp 1649977179
transform 1 0 34132 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1649977179
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_367
timestamp 1649977179
transform 1 0 34868 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_378
timestamp 1649977179
transform 1 0 35880 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_385
timestamp 1649977179
transform 1 0 36524 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_400
timestamp 1649977179
transform 1 0 37904 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_409
timestamp 1649977179
transform 1 0 38732 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_416
timestamp 1649977179
transform 1 0 39376 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_423
timestamp 1649977179
transform 1 0 40020 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_429
timestamp 1649977179
transform 1 0 40572 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_435
timestamp 1649977179
transform 1 0 41124 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_447
timestamp 1649977179
transform 1 0 42228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_459
timestamp 1649977179
transform 1 0 43332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_471
timestamp 1649977179
transform 1 0 44436 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1649977179
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1649977179
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1649977179
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1649977179
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_513
timestamp 1649977179
transform 1 0 48300 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1649977179
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1649977179
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1649977179
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1649977179
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1649977179
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1649977179
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1649977179
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1649977179
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1649977179
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_93
timestamp 1649977179
transform 1 0 9660 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_99
timestamp 1649977179
transform 1 0 10212 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_102
timestamp 1649977179
transform 1 0 10488 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_108
timestamp 1649977179
transform 1 0 11040 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_113
timestamp 1649977179
transform 1 0 11500 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_117
timestamp 1649977179
transform 1 0 11868 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_123
timestamp 1649977179
transform 1 0 12420 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_132
timestamp 1649977179
transform 1 0 13248 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_142
timestamp 1649977179
transform 1 0 14168 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_148
timestamp 1649977179
transform 1 0 14720 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_154
timestamp 1649977179
transform 1 0 15272 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_164
timestamp 1649977179
transform 1 0 16192 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_172
timestamp 1649977179
transform 1 0 16928 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_178
timestamp 1649977179
transform 1 0 17480 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_184
timestamp 1649977179
transform 1 0 18032 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_195
timestamp 1649977179
transform 1 0 19044 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_201
timestamp 1649977179
transform 1 0 19596 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_207
timestamp 1649977179
transform 1 0 20148 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_213
timestamp 1649977179
transform 1 0 20700 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_220
timestamp 1649977179
transform 1 0 21344 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_233
timestamp 1649977179
transform 1 0 22540 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_240
timestamp 1649977179
transform 1 0 23184 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_250
timestamp 1649977179
transform 1 0 24104 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_259
timestamp 1649977179
transform 1 0 24932 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_266
timestamp 1649977179
transform 1 0 25576 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_270
timestamp 1649977179
transform 1 0 25944 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1649977179
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1649977179
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_281
timestamp 1649977179
transform 1 0 26956 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_299
timestamp 1649977179
transform 1 0 28612 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_322
timestamp 1649977179
transform 1 0 30728 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_328
timestamp 1649977179
transform 1 0 31280 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_354
timestamp 1649977179
transform 1 0 33672 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_360
timestamp 1649977179
transform 1 0 34224 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_368
timestamp 1649977179
transform 1 0 34960 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_375
timestamp 1649977179
transform 1 0 35604 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_384
timestamp 1649977179
transform 1 0 36432 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_400
timestamp 1649977179
transform 1 0 37904 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_408
timestamp 1649977179
transform 1 0 38640 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_415
timestamp 1649977179
transform 1 0 39284 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_421
timestamp 1649977179
transform 1 0 39836 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_427
timestamp 1649977179
transform 1 0 40388 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_433
timestamp 1649977179
transform 1 0 40940 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_445
timestamp 1649977179
transform 1 0 42044 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1649977179
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1649977179
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1649977179
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1649977179
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1649977179
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1649977179
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_505
timestamp 1649977179
transform 1 0 47564 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_513
timestamp 1649977179
transform 1 0 48300 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_7
timestamp 1649977179
transform 1 0 1748 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_13
timestamp 1649977179
transform 1 0 2300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_25
timestamp 1649977179
transform 1 0 3404 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1649977179
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1649977179
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1649977179
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1649977179
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1649977179
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1649977179
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_85
timestamp 1649977179
transform 1 0 8924 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_93
timestamp 1649977179
transform 1 0 9660 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_99
timestamp 1649977179
transform 1 0 10212 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_105
timestamp 1649977179
transform 1 0 10764 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_111
timestamp 1649977179
transform 1 0 11316 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_117
timestamp 1649977179
transform 1 0 11868 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_128
timestamp 1649977179
transform 1 0 12880 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_136
timestamp 1649977179
transform 1 0 13616 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_141
timestamp 1649977179
transform 1 0 14076 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_145
timestamp 1649977179
transform 1 0 14444 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_151
timestamp 1649977179
transform 1 0 14996 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_161
timestamp 1649977179
transform 1 0 15916 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_169
timestamp 1649977179
transform 1 0 16652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_175
timestamp 1649977179
transform 1 0 17204 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_74_186
timestamp 1649977179
transform 1 0 18216 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_192
timestamp 1649977179
transform 1 0 18768 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_203
timestamp 1649977179
transform 1 0 19780 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_215
timestamp 1649977179
transform 1 0 20884 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_229
timestamp 1649977179
transform 1 0 22172 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_238
timestamp 1649977179
transform 1 0 23000 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_242
timestamp 1649977179
transform 1 0 23368 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_248
timestamp 1649977179
transform 1 0 23920 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_259
timestamp 1649977179
transform 1 0 24932 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_268
timestamp 1649977179
transform 1 0 25760 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_274
timestamp 1649977179
transform 1 0 26312 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_280
timestamp 1649977179
transform 1 0 26864 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_284
timestamp 1649977179
transform 1 0 27232 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_304
timestamp 1649977179
transform 1 0 29072 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_328
timestamp 1649977179
transform 1 0 31280 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_351
timestamp 1649977179
transform 1 0 33396 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_360
timestamp 1649977179
transform 1 0 34224 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_374
timestamp 1649977179
transform 1 0 35512 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_386
timestamp 1649977179
transform 1 0 36616 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_397
timestamp 1649977179
transform 1 0 37628 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_405
timestamp 1649977179
transform 1 0 38364 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_411
timestamp 1649977179
transform 1 0 38916 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1649977179
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_423
timestamp 1649977179
transform 1 0 40020 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_429
timestamp 1649977179
transform 1 0 40572 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_441
timestamp 1649977179
transform 1 0 41676 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_453
timestamp 1649977179
transform 1 0 42780 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_465
timestamp 1649977179
transform 1 0 43884 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_473
timestamp 1649977179
transform 1 0 44620 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1649977179
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1649977179
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_501
timestamp 1649977179
transform 1 0 47196 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_505
timestamp 1649977179
transform 1 0 47564 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_512
timestamp 1649977179
transform 1 0 48208 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1649977179
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1649977179
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1649977179
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1649977179
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1649977179
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1649977179
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1649977179
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1649977179
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1649977179
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_93
timestamp 1649977179
transform 1 0 9660 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_96
timestamp 1649977179
transform 1 0 9936 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_102
timestamp 1649977179
transform 1 0 10488 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_108
timestamp 1649977179
transform 1 0 11040 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_113
timestamp 1649977179
transform 1 0 11500 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_116
timestamp 1649977179
transform 1 0 11776 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_122
timestamp 1649977179
transform 1 0 12328 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_129
timestamp 1649977179
transform 1 0 12972 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_140
timestamp 1649977179
transform 1 0 13984 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_144
timestamp 1649977179
transform 1 0 14352 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_152
timestamp 1649977179
transform 1 0 15088 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_156
timestamp 1649977179
transform 1 0 15456 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_164
timestamp 1649977179
transform 1 0 16192 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_172
timestamp 1649977179
transform 1 0 16928 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_176
timestamp 1649977179
transform 1 0 17296 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_183
timestamp 1649977179
transform 1 0 17940 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_195
timestamp 1649977179
transform 1 0 19044 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_199
timestamp 1649977179
transform 1 0 19412 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_207
timestamp 1649977179
transform 1 0 20148 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1649977179
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1649977179
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_233
timestamp 1649977179
transform 1 0 22540 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_245
timestamp 1649977179
transform 1 0 23644 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_256
timestamp 1649977179
transform 1 0 24656 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_276
timestamp 1649977179
transform 1 0 26496 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_283
timestamp 1649977179
transform 1 0 27140 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_289
timestamp 1649977179
transform 1 0 27692 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_295
timestamp 1649977179
transform 1 0 28244 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_319
timestamp 1649977179
transform 1 0 30452 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_325
timestamp 1649977179
transform 1 0 31004 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_331
timestamp 1649977179
transform 1 0 31556 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1649977179
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_354
timestamp 1649977179
transform 1 0 33672 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_375
timestamp 1649977179
transform 1 0 35604 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_386
timestamp 1649977179
transform 1 0 36616 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_393
timestamp 1649977179
transform 1 0 37260 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_397
timestamp 1649977179
transform 1 0 37628 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_401
timestamp 1649977179
transform 1 0 37996 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_408
timestamp 1649977179
transform 1 0 38640 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_414
timestamp 1649977179
transform 1 0 39192 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_420
timestamp 1649977179
transform 1 0 39744 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_426
timestamp 1649977179
transform 1 0 40296 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_438
timestamp 1649977179
transform 1 0 41400 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_446
timestamp 1649977179
transform 1 0 42136 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1649977179
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1649977179
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1649977179
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1649977179
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1649977179
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1649977179
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_505
timestamp 1649977179
transform 1 0 47564 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_513
timestamp 1649977179
transform 1 0 48300 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_5
timestamp 1649977179
transform 1 0 1564 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_17
timestamp 1649977179
transform 1 0 2668 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_25
timestamp 1649977179
transform 1 0 3404 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1649977179
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1649977179
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1649977179
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1649977179
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1649977179
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1649977179
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_85
timestamp 1649977179
transform 1 0 8924 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_95
timestamp 1649977179
transform 1 0 9844 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_101
timestamp 1649977179
transform 1 0 10396 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_107
timestamp 1649977179
transform 1 0 10948 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_113
timestamp 1649977179
transform 1 0 11500 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_119
timestamp 1649977179
transform 1 0 12052 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_125
timestamp 1649977179
transform 1 0 12604 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_136
timestamp 1649977179
transform 1 0 13616 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_76_141
timestamp 1649977179
transform 1 0 14076 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_146
timestamp 1649977179
transform 1 0 14536 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_153
timestamp 1649977179
transform 1 0 15180 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_161
timestamp 1649977179
transform 1 0 15916 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_168
timestamp 1649977179
transform 1 0 16560 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_174
timestamp 1649977179
transform 1 0 17112 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_180
timestamp 1649977179
transform 1 0 17664 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_192
timestamp 1649977179
transform 1 0 18768 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_197
timestamp 1649977179
transform 1 0 19228 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_205
timestamp 1649977179
transform 1 0 19964 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_214
timestamp 1649977179
transform 1 0 20792 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_223
timestamp 1649977179
transform 1 0 21620 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_227
timestamp 1649977179
transform 1 0 21988 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_231
timestamp 1649977179
transform 1 0 22356 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_237
timestamp 1649977179
transform 1 0 22908 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_240
timestamp 1649977179
transform 1 0 23184 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_248
timestamp 1649977179
transform 1 0 23920 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_259
timestamp 1649977179
transform 1 0 24932 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_268
timestamp 1649977179
transform 1 0 25760 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_274
timestamp 1649977179
transform 1 0 26312 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_278
timestamp 1649977179
transform 1 0 26680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_281
timestamp 1649977179
transform 1 0 26956 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_304
timestamp 1649977179
transform 1 0 29072 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_311
timestamp 1649977179
transform 1 0 29716 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_315
timestamp 1649977179
transform 1 0 30084 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_318
timestamp 1649977179
transform 1 0 30360 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_326
timestamp 1649977179
transform 1 0 31096 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_347
timestamp 1649977179
transform 1 0 33028 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_353
timestamp 1649977179
transform 1 0 33580 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_359
timestamp 1649977179
transform 1 0 34132 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1649977179
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_371
timestamp 1649977179
transform 1 0 35236 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_379
timestamp 1649977179
transform 1 0 35972 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_387
timestamp 1649977179
transform 1 0 36708 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_395
timestamp 1649977179
transform 1 0 37444 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_401
timestamp 1649977179
transform 1 0 37996 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_407
timestamp 1649977179
transform 1 0 38548 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1649977179
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1649977179
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1649977179
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1649977179
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1649977179
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1649977179
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1649977179
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1649977179
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1649977179
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1649977179
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_501
timestamp 1649977179
transform 1 0 47196 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_509
timestamp 1649977179
transform 1 0 47932 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_512
timestamp 1649977179
transform 1 0 48208 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_7
timestamp 1649977179
transform 1 0 1748 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_19
timestamp 1649977179
transform 1 0 2852 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_31
timestamp 1649977179
transform 1 0 3956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_43
timestamp 1649977179
transform 1 0 5060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1649977179
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1649977179
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1649977179
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_81
timestamp 1649977179
transform 1 0 8556 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_87
timestamp 1649977179
transform 1 0 9108 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_90
timestamp 1649977179
transform 1 0 9384 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_96
timestamp 1649977179
transform 1 0 9936 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_102
timestamp 1649977179
transform 1 0 10488 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_108
timestamp 1649977179
transform 1 0 11040 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_77_113
timestamp 1649977179
transform 1 0 11500 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_118
timestamp 1649977179
transform 1 0 11960 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_127
timestamp 1649977179
transform 1 0 12788 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_134
timestamp 1649977179
transform 1 0 13432 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_140
timestamp 1649977179
transform 1 0 13984 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_143
timestamp 1649977179
transform 1 0 14260 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_149
timestamp 1649977179
transform 1 0 14812 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_158
timestamp 1649977179
transform 1 0 15640 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_164
timestamp 1649977179
transform 1 0 16192 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_174
timestamp 1649977179
transform 1 0 17112 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_180
timestamp 1649977179
transform 1 0 17664 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_190
timestamp 1649977179
transform 1 0 18584 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_200
timestamp 1649977179
transform 1 0 19504 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_209
timestamp 1649977179
transform 1 0 20332 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_216
timestamp 1649977179
transform 1 0 20976 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_77_231
timestamp 1649977179
transform 1 0 22356 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_239
timestamp 1649977179
transform 1 0 23092 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_242
timestamp 1649977179
transform 1 0 23368 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_249
timestamp 1649977179
transform 1 0 24012 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_258
timestamp 1649977179
transform 1 0 24840 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_77_266
timestamp 1649977179
transform 1 0 25576 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_272
timestamp 1649977179
transform 1 0 26128 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_281
timestamp 1649977179
transform 1 0 26956 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_299
timestamp 1649977179
transform 1 0 28612 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_322
timestamp 1649977179
transform 1 0 30728 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_77_332
timestamp 1649977179
transform 1 0 31648 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_354
timestamp 1649977179
transform 1 0 33672 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_360
timestamp 1649977179
transform 1 0 34224 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_367
timestamp 1649977179
transform 1 0 34868 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_376
timestamp 1649977179
transform 1 0 35696 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_382
timestamp 1649977179
transform 1 0 36248 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_388
timestamp 1649977179
transform 1 0 36800 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_395
timestamp 1649977179
transform 1 0 37444 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_401
timestamp 1649977179
transform 1 0 37996 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_413
timestamp 1649977179
transform 1 0 39100 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_425
timestamp 1649977179
transform 1 0 40204 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_437
timestamp 1649977179
transform 1 0 41308 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_445
timestamp 1649977179
transform 1 0 42044 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1649977179
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1649977179
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1649977179
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1649977179
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1649977179
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1649977179
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_77_505
timestamp 1649977179
transform 1 0 47564 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_512
timestamp 1649977179
transform 1 0 48208 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1649977179
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1649977179
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1649977179
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1649977179
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1649977179
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1649977179
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1649977179
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1649977179
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1649977179
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1649977179
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_99
timestamp 1649977179
transform 1 0 10212 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_105
timestamp 1649977179
transform 1 0 10764 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_111
timestamp 1649977179
transform 1 0 11316 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_117
timestamp 1649977179
transform 1 0 11868 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_123
timestamp 1649977179
transform 1 0 12420 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_130
timestamp 1649977179
transform 1 0 13064 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_136
timestamp 1649977179
transform 1 0 13616 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_149
timestamp 1649977179
transform 1 0 14812 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_153
timestamp 1649977179
transform 1 0 15180 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_157
timestamp 1649977179
transform 1 0 15548 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_163
timestamp 1649977179
transform 1 0 16100 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_174
timestamp 1649977179
transform 1 0 17112 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_180
timestamp 1649977179
transform 1 0 17664 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_186
timestamp 1649977179
transform 1 0 18216 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_192
timestamp 1649977179
transform 1 0 18768 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_200
timestamp 1649977179
transform 1 0 19504 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_204
timestamp 1649977179
transform 1 0 19872 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_207
timestamp 1649977179
transform 1 0 20148 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_218
timestamp 1649977179
transform 1 0 21160 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_229
timestamp 1649977179
transform 1 0 22172 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_236
timestamp 1649977179
transform 1 0 22816 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_242
timestamp 1649977179
transform 1 0 23368 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_248
timestamp 1649977179
transform 1 0 23920 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_253
timestamp 1649977179
transform 1 0 24380 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_262
timestamp 1649977179
transform 1 0 25208 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_268
timestamp 1649977179
transform 1 0 25760 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_274
timestamp 1649977179
transform 1 0 26312 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_78_299
timestamp 1649977179
transform 1 0 28612 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1649977179
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_328
timestamp 1649977179
transform 1 0 31280 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_78_338
timestamp 1649977179
transform 1 0 32200 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_346
timestamp 1649977179
transform 1 0 32936 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_350
timestamp 1649977179
transform 1 0 33304 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_356
timestamp 1649977179
transform 1 0 33856 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_370
timestamp 1649977179
transform 1 0 35144 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_376
timestamp 1649977179
transform 1 0 35696 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_382
timestamp 1649977179
transform 1 0 36248 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_394
timestamp 1649977179
transform 1 0 37352 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_406
timestamp 1649977179
transform 1 0 38456 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_418
timestamp 1649977179
transform 1 0 39560 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1649977179
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1649977179
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1649977179
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1649977179
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1649977179
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1649977179
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1649977179
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1649977179
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_501
timestamp 1649977179
transform 1 0 47196 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_509
timestamp 1649977179
transform 1 0 47932 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_512
timestamp 1649977179
transform 1 0 48208 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_3
timestamp 1649977179
transform 1 0 1380 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_7
timestamp 1649977179
transform 1 0 1748 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_19
timestamp 1649977179
transform 1 0 2852 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_31
timestamp 1649977179
transform 1 0 3956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_43
timestamp 1649977179
transform 1 0 5060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1649977179
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1649977179
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1649977179
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_81
timestamp 1649977179
transform 1 0 8556 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_89
timestamp 1649977179
transform 1 0 9292 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_79_94
timestamp 1649977179
transform 1 0 9752 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_79_102
timestamp 1649977179
transform 1 0 10488 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_108
timestamp 1649977179
transform 1 0 11040 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_113
timestamp 1649977179
transform 1 0 11500 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_119
timestamp 1649977179
transform 1 0 12052 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_125
timestamp 1649977179
transform 1 0 12604 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_133
timestamp 1649977179
transform 1 0 13340 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_144
timestamp 1649977179
transform 1 0 14352 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_150
timestamp 1649977179
transform 1 0 14904 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1649977179
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1649977179
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_173
timestamp 1649977179
transform 1 0 17020 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_180
timestamp 1649977179
transform 1 0 17664 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_79_190
timestamp 1649977179
transform 1 0 18584 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_201
timestamp 1649977179
transform 1 0 19596 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_211
timestamp 1649977179
transform 1 0 20516 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_220
timestamp 1649977179
transform 1 0 21344 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_233
timestamp 1649977179
transform 1 0 22540 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_244
timestamp 1649977179
transform 1 0 23552 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_255
timestamp 1649977179
transform 1 0 24564 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_266
timestamp 1649977179
transform 1 0 25576 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_274
timestamp 1649977179
transform 1 0 26312 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_79_281
timestamp 1649977179
transform 1 0 26956 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_287
timestamp 1649977179
transform 1 0 27508 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_314
timestamp 1649977179
transform 1 0 29992 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_320
timestamp 1649977179
transform 1 0 30544 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_326
timestamp 1649977179
transform 1 0 31096 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_332
timestamp 1649977179
transform 1 0 31648 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_353
timestamp 1649977179
transform 1 0 33580 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_357
timestamp 1649977179
transform 1 0 33948 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_360
timestamp 1649977179
transform 1 0 34224 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_367
timestamp 1649977179
transform 1 0 34868 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1649977179
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1649977179
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1649977179
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1649977179
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1649977179
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1649977179
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1649977179
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1649977179
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1649977179
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1649977179
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1649977179
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1649977179
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1649977179
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1649977179
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1649977179
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_505
timestamp 1649977179
transform 1 0 47564 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_509
timestamp 1649977179
transform 1 0 47932 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_512
timestamp 1649977179
transform 1 0 48208 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_3
timestamp 1649977179
transform 1 0 1380 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_11
timestamp 1649977179
transform 1 0 2116 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_17
timestamp 1649977179
transform 1 0 2668 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_25
timestamp 1649977179
transform 1 0 3404 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1649977179
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1649977179
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1649977179
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1649977179
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1649977179
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1649977179
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_85
timestamp 1649977179
transform 1 0 8924 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_88
timestamp 1649977179
transform 1 0 9200 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_94
timestamp 1649977179
transform 1 0 9752 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_100
timestamp 1649977179
transform 1 0 10304 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_106
timestamp 1649977179
transform 1 0 10856 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_112
timestamp 1649977179
transform 1 0 11408 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_118
timestamp 1649977179
transform 1 0 11960 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_124
timestamp 1649977179
transform 1 0 12512 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_130
timestamp 1649977179
transform 1 0 13064 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_136
timestamp 1649977179
transform 1 0 13616 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_150
timestamp 1649977179
transform 1 0 14904 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_158
timestamp 1649977179
transform 1 0 15640 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_161
timestamp 1649977179
transform 1 0 15916 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_171
timestamp 1649977179
transform 1 0 16836 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_179
timestamp 1649977179
transform 1 0 17572 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_183
timestamp 1649977179
transform 1 0 17940 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_192
timestamp 1649977179
transform 1 0 18768 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_205
timestamp 1649977179
transform 1 0 19964 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_211
timestamp 1649977179
transform 1 0 20516 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_220
timestamp 1649977179
transform 1 0 21344 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_232
timestamp 1649977179
transform 1 0 22448 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_240
timestamp 1649977179
transform 1 0 23184 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_248
timestamp 1649977179
transform 1 0 23920 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_260
timestamp 1649977179
transform 1 0 25024 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_283
timestamp 1649977179
transform 1 0 27140 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_304
timestamp 1649977179
transform 1 0 29072 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_309
timestamp 1649977179
transform 1 0 29532 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_313
timestamp 1649977179
transform 1 0 29900 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_333
timestamp 1649977179
transform 1 0 31740 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_354
timestamp 1649977179
transform 1 0 33672 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_360
timestamp 1649977179
transform 1 0 34224 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_365
timestamp 1649977179
transform 1 0 34684 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_369
timestamp 1649977179
transform 1 0 35052 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_381
timestamp 1649977179
transform 1 0 36156 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_393
timestamp 1649977179
transform 1 0 37260 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_405
timestamp 1649977179
transform 1 0 38364 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_417
timestamp 1649977179
transform 1 0 39468 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1649977179
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1649977179
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1649977179
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1649977179
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1649977179
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1649977179
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1649977179
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_489
timestamp 1649977179
transform 1 0 46092 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_493
timestamp 1649977179
transform 1 0 46460 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_496
timestamp 1649977179
transform 1 0 46736 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_502
timestamp 1649977179
transform 1 0 47288 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_512
timestamp 1649977179
transform 1 0 48208 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_7
timestamp 1649977179
transform 1 0 1748 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_81_17
timestamp 1649977179
transform 1 0 2668 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_23
timestamp 1649977179
transform 1 0 3220 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_35
timestamp 1649977179
transform 1 0 4324 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_47
timestamp 1649977179
transform 1 0 5428 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1649977179
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_57
timestamp 1649977179
transform 1 0 6348 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_63
timestamp 1649977179
transform 1 0 6900 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_75
timestamp 1649977179
transform 1 0 8004 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_81
timestamp 1649977179
transform 1 0 8556 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_84
timestamp 1649977179
transform 1 0 8832 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_90
timestamp 1649977179
transform 1 0 9384 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_96
timestamp 1649977179
transform 1 0 9936 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_102
timestamp 1649977179
transform 1 0 10488 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_108
timestamp 1649977179
transform 1 0 11040 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_113
timestamp 1649977179
transform 1 0 11500 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_118
timestamp 1649977179
transform 1 0 11960 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_124
timestamp 1649977179
transform 1 0 12512 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_131
timestamp 1649977179
transform 1 0 13156 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_142
timestamp 1649977179
transform 1 0 14168 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_149
timestamp 1649977179
transform 1 0 14812 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_160
timestamp 1649977179
transform 1 0 15824 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_81_176
timestamp 1649977179
transform 1 0 17296 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_81_187
timestamp 1649977179
transform 1 0 18308 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_198
timestamp 1649977179
transform 1 0 19320 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_206
timestamp 1649977179
transform 1 0 20056 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_214
timestamp 1649977179
transform 1 0 20792 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_218
timestamp 1649977179
transform 1 0 21160 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_238
timestamp 1649977179
transform 1 0 23000 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_248
timestamp 1649977179
transform 1 0 23920 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_255
timestamp 1649977179
transform 1 0 24564 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_276
timestamp 1649977179
transform 1 0 26496 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_291
timestamp 1649977179
transform 1 0 27876 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_295
timestamp 1649977179
transform 1 0 28244 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_315
timestamp 1649977179
transform 1 0 30084 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_321
timestamp 1649977179
transform 1 0 30636 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_81_332
timestamp 1649977179
transform 1 0 31648 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_354
timestamp 1649977179
transform 1 0 33672 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_362
timestamp 1649977179
transform 1 0 34408 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_368
timestamp 1649977179
transform 1 0 34960 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_373
timestamp 1649977179
transform 1 0 35420 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_379
timestamp 1649977179
transform 1 0 35972 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1649977179
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1649977179
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1649977179
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1649977179
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1649977179
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1649977179
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1649977179
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_451
timestamp 1649977179
transform 1 0 42596 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_463
timestamp 1649977179
transform 1 0 43700 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_475
timestamp 1649977179
transform 1 0 44804 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_481
timestamp 1649977179
transform 1 0 45356 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_489
timestamp 1649977179
transform 1 0 46092 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_492
timestamp 1649977179
transform 1 0 46368 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_500
timestamp 1649977179
transform 1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_505
timestamp 1649977179
transform 1 0 47564 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_512
timestamp 1649977179
transform 1 0 48208 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_13
timestamp 1649977179
transform 1 0 2300 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_21
timestamp 1649977179
transform 1 0 3036 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1649977179
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_29
timestamp 1649977179
transform 1 0 3772 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_34
timestamp 1649977179
transform 1 0 4232 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_40
timestamp 1649977179
transform 1 0 4784 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_52
timestamp 1649977179
transform 1 0 5888 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_61
timestamp 1649977179
transform 1 0 6716 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_69
timestamp 1649977179
transform 1 0 7452 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1649977179
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1649977179
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_82_85
timestamp 1649977179
transform 1 0 8924 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_90
timestamp 1649977179
transform 1 0 9384 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_104
timestamp 1649977179
transform 1 0 10672 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_113
timestamp 1649977179
transform 1 0 11500 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_121
timestamp 1649977179
transform 1 0 12236 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_125
timestamp 1649977179
transform 1 0 12604 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_128
timestamp 1649977179
transform 1 0 12880 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_136
timestamp 1649977179
transform 1 0 13616 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_146
timestamp 1649977179
transform 1 0 14536 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_154
timestamp 1649977179
transform 1 0 15272 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_163
timestamp 1649977179
transform 1 0 16100 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_167
timestamp 1649977179
transform 1 0 16468 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_82_169
timestamp 1649977179
transform 1 0 16652 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_174
timestamp 1649977179
transform 1 0 17112 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_188
timestamp 1649977179
transform 1 0 18400 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_197
timestamp 1649977179
transform 1 0 19228 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_203
timestamp 1649977179
transform 1 0 19780 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_207
timestamp 1649977179
transform 1 0 20148 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_210
timestamp 1649977179
transform 1 0 20424 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_220
timestamp 1649977179
transform 1 0 21344 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_225
timestamp 1649977179
transform 1 0 21804 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_232
timestamp 1649977179
transform 1 0 22448 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_240
timestamp 1649977179
transform 1 0 23184 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1649977179
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1649977179
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_256
timestamp 1649977179
transform 1 0 24656 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_276
timestamp 1649977179
transform 1 0 26496 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_82_281
timestamp 1649977179
transform 1 0 26956 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_304
timestamp 1649977179
transform 1 0 29072 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_328
timestamp 1649977179
transform 1 0 31280 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_354
timestamp 1649977179
transform 1 0 33672 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_360
timestamp 1649977179
transform 1 0 34224 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_382
timestamp 1649977179
transform 1 0 36248 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_388
timestamp 1649977179
transform 1 0 36800 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_397
timestamp 1649977179
transform 1 0 37628 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_405
timestamp 1649977179
transform 1 0 38364 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_412
timestamp 1649977179
transform 1 0 39008 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_421
timestamp 1649977179
transform 1 0 39836 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_426
timestamp 1649977179
transform 1 0 40296 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_434
timestamp 1649977179
transform 1 0 41032 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_446
timestamp 1649977179
transform 1 0 42136 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_449
timestamp 1649977179
transform 1 0 42412 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_455
timestamp 1649977179
transform 1 0 42964 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_467
timestamp 1649977179
transform 1 0 44068 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1649977179
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_477
timestamp 1649977179
transform 1 0 44988 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_485
timestamp 1649977179
transform 1 0 45724 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_82_497
timestamp 1649977179
transform 1 0 46828 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_503
timestamp 1649977179
transform 1 0 47380 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_82_505
timestamp 1649977179
transform 1 0 47564 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_512
timestamp 1649977179
transform 1 0 48208 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1649977179
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1649977179
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1649977179
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1649977179
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1649977179
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1649977179
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1649977179
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1649977179
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1649977179
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1649977179
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1649977179
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1649977179
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1649977179
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1649977179
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1649977179
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1649977179
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1649977179
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1649977179
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1649977179
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1649977179
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1649977179
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1649977179
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1649977179
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1649977179
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1649977179
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1649977179
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1649977179
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1649977179
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1649977179
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1649977179
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1649977179
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1649977179
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1649977179
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1649977179
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1649977179
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1649977179
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1649977179
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1649977179
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1649977179
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1649977179
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1649977179
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1649977179
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1649977179
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1649977179
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1649977179
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1649977179
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1649977179
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1649977179
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1649977179
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1649977179
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1649977179
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1649977179
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1649977179
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1649977179
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1649977179
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1649977179
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1649977179
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1649977179
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1649977179
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1649977179
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1649977179
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1649977179
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1649977179
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1649977179
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1649977179
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1649977179
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1649977179
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1649977179
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1649977179
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1649977179
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1649977179
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1649977179
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1649977179
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1649977179
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1649977179
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1649977179
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1649977179
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1649977179
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1649977179
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1649977179
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1649977179
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1649977179
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1649977179
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1649977179
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1649977179
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1649977179
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1649977179
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1649977179
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1649977179
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1649977179
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1649977179
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1649977179
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1649977179
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1649977179
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1649977179
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1649977179
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1649977179
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1649977179
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1649977179
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1649977179
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1649977179
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1649977179
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1649977179
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1649977179
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1649977179
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1649977179
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1649977179
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1649977179
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1649977179
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1649977179
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1649977179
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1649977179
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1649977179
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1649977179
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1649977179
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1649977179
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1649977179
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1649977179
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1649977179
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1649977179
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1649977179
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1649977179
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1649977179
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1649977179
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1649977179
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1649977179
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1649977179
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1649977179
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1649977179
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1649977179
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1649977179
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1649977179
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1649977179
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1649977179
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1649977179
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1649977179
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1649977179
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1649977179
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1649977179
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1649977179
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1649977179
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1649977179
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1649977179
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1649977179
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1649977179
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1649977179
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1649977179
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1649977179
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1649977179
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1649977179
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1649977179
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1649977179
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1649977179
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1649977179
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1649977179
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1649977179
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1649977179
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1649977179
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1649977179
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1649977179
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1649977179
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1649977179
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1649977179
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1649977179
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1649977179
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1649977179
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1649977179
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1649977179
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1649977179
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1649977179
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1649977179
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1649977179
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1649977179
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1649977179
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1649977179
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1649977179
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1649977179
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1649977179
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1649977179
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1649977179
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1649977179
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1649977179
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1649977179
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1649977179
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1649977179
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1649977179
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1649977179
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1649977179
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1649977179
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1649977179
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1649977179
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1649977179
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1649977179
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1649977179
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1649977179
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1649977179
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1649977179
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1649977179
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1649977179
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1649977179
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1649977179
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1649977179
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1649977179
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1649977179
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1649977179
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1649977179
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1649977179
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1649977179
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1649977179
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1649977179
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1649977179
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1649977179
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1649977179
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1649977179
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1649977179
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1649977179
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1649977179
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1649977179
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1649977179
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1649977179
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1649977179
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1649977179
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1649977179
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1649977179
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1649977179
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1649977179
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1649977179
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1649977179
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1649977179
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1649977179
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1649977179
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1649977179
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1649977179
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1649977179
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1649977179
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1649977179
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1649977179
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1649977179
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1649977179
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1649977179
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1649977179
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1649977179
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1649977179
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1649977179
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1649977179
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1649977179
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1649977179
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1649977179
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1649977179
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1649977179
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _0732_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12696 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0733_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12236 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0734_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12972 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0735_
timestamp 1649977179
transform 1 0 15272 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0736_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14996 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0737_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12788 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0738_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13984 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0739_
timestamp 1649977179
transform 1 0 12328 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0740_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13156 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0741_
timestamp 1649977179
transform -1 0 13064 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0742_
timestamp 1649977179
transform 1 0 13708 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0743_
timestamp 1649977179
transform 1 0 15272 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0744_
timestamp 1649977179
transform 1 0 16468 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0745_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 31648 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0746_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 31464 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _0747_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 34040 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0748_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14720 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0749_
timestamp 1649977179
transform -1 0 14352 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0750_
timestamp 1649977179
transform 1 0 14444 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0751_
timestamp 1649977179
transform -1 0 16560 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0752_
timestamp 1649977179
transform 1 0 14904 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0753_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15364 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0754_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15088 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0755_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 32292 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0756_
timestamp 1649977179
transform -1 0 48024 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0757_
timestamp 1649977179
transform -1 0 30636 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0758_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 29992 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0759_
timestamp 1649977179
transform -1 0 16192 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _0760_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 34408 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _0761_
timestamp 1649977179
transform -1 0 31464 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0762_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 32568 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0763_
timestamp 1649977179
transform 1 0 33396 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0764_
timestamp 1649977179
transform -1 0 17940 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0765_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17480 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0766_
timestamp 1649977179
transform -1 0 17940 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0767_
timestamp 1649977179
transform 1 0 24472 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0768_
timestamp 1649977179
transform -1 0 22724 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0769_
timestamp 1649977179
transform -1 0 14536 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0770_
timestamp 1649977179
transform 1 0 14536 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0771_
timestamp 1649977179
transform -1 0 13156 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0772_
timestamp 1649977179
transform 1 0 12972 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0773_
timestamp 1649977179
transform 1 0 13524 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0774_
timestamp 1649977179
transform 1 0 15180 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0775_
timestamp 1649977179
transform 1 0 17388 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0776_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16652 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0777_
timestamp 1649977179
transform 1 0 16652 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0778_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 31464 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0779_
timestamp 1649977179
transform 1 0 32476 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0780_
timestamp 1649977179
transform 1 0 16744 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0781_
timestamp 1649977179
transform -1 0 16928 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0782_
timestamp 1649977179
transform 1 0 16652 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1649977179
transform 1 0 15732 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0784_
timestamp 1649977179
transform -1 0 16008 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0785_
timestamp 1649977179
transform 1 0 16652 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0786_
timestamp 1649977179
transform 1 0 17112 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1649977179
transform 1 0 34684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0788_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18032 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0789_
timestamp 1649977179
transform -1 0 18584 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0790_
timestamp 1649977179
transform -1 0 24564 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0791_
timestamp 1649977179
transform -1 0 25208 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0792_
timestamp 1649977179
transform -1 0 24656 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0793_
timestamp 1649977179
transform -1 0 14812 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_2  _0794_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 14904 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0795_
timestamp 1649977179
transform -1 0 19596 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0796_
timestamp 1649977179
transform 1 0 18308 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0797_
timestamp 1649977179
transform -1 0 17940 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0798_
timestamp 1649977179
transform 1 0 18032 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0799_
timestamp 1649977179
transform 1 0 15640 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0800_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16284 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0801_
timestamp 1649977179
transform 1 0 18676 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0802_
timestamp 1649977179
transform -1 0 20332 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0803_
timestamp 1649977179
transform 1 0 20700 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0804_
timestamp 1649977179
transform -1 0 19504 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0805_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15640 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0806_
timestamp 1649977179
transform 1 0 18308 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0807_
timestamp 1649977179
transform 1 0 18400 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0808_
timestamp 1649977179
transform -1 0 18768 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0809_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20700 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0810_
timestamp 1649977179
transform -1 0 19412 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0811_
timestamp 1649977179
transform 1 0 19136 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0812_
timestamp 1649977179
transform -1 0 20056 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0813_
timestamp 1649977179
transform 1 0 20884 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0814_
timestamp 1649977179
transform 1 0 20884 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0815_
timestamp 1649977179
transform 1 0 20884 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0816_
timestamp 1649977179
transform 1 0 25944 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0817_
timestamp 1649977179
transform -1 0 25576 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0818_
timestamp 1649977179
transform -1 0 24012 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0819_
timestamp 1649977179
transform 1 0 23460 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0820_
timestamp 1649977179
transform -1 0 24656 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0821_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19228 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0822_
timestamp 1649977179
transform -1 0 23920 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0823_
timestamp 1649977179
transform 1 0 24380 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _0824_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19228 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0825_
timestamp 1649977179
transform -1 0 21344 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0826_
timestamp 1649977179
transform 1 0 21160 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0827_
timestamp 1649977179
transform -1 0 20792 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0828_
timestamp 1649977179
transform 1 0 20516 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0829_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 19964 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0830_
timestamp 1649977179
transform -1 0 47104 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0831_
timestamp 1649977179
transform -1 0 34868 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _0832_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 32016 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _0833_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19228 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0834_
timestamp 1649977179
transform 1 0 20240 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0835_
timestamp 1649977179
transform -1 0 19872 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0836_
timestamp 1649977179
transform -1 0 20148 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0837_
timestamp 1649977179
transform 1 0 30912 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0838_
timestamp 1649977179
transform -1 0 23644 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0839_
timestamp 1649977179
transform 1 0 24380 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _0840_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21804 0 -1 46784
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_1  _0841_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 23920 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0842_
timestamp 1649977179
transform -1 0 22448 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0843_
timestamp 1649977179
transform 1 0 22540 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0844_
timestamp 1649977179
transform 1 0 23920 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0845_
timestamp 1649977179
transform 1 0 25300 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0846_
timestamp 1649977179
transform -1 0 25576 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0847_
timestamp 1649977179
transform -1 0 24840 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0848_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 24472 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0849_
timestamp 1649977179
transform 1 0 23736 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0850_
timestamp 1649977179
transform 1 0 21068 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0851_
timestamp 1649977179
transform 1 0 21804 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0852_
timestamp 1649977179
transform 1 0 22632 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0853_
timestamp 1649977179
transform -1 0 22540 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0854_
timestamp 1649977179
transform -1 0 20884 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0855_
timestamp 1649977179
transform 1 0 21804 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0856_
timestamp 1649977179
transform 1 0 23920 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0857_
timestamp 1649977179
transform 1 0 24472 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _0858_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 25300 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0859_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 24656 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0860_
timestamp 1649977179
transform 1 0 21528 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0861_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 22540 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0862_
timestamp 1649977179
transform 1 0 22908 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0863_
timestamp 1649977179
transform 1 0 34592 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0864_
timestamp 1649977179
transform 1 0 34684 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0865_
timestamp 1649977179
transform -1 0 35696 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0866_
timestamp 1649977179
transform 1 0 34684 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0867_
timestamp 1649977179
transform -1 0 36708 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0868_
timestamp 1649977179
transform -1 0 34224 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0869_
timestamp 1649977179
transform 1 0 18308 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0870_
timestamp 1649977179
transform -1 0 23000 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0871_
timestamp 1649977179
transform 1 0 22080 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0872_
timestamp 1649977179
transform -1 0 23184 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0873_
timestamp 1649977179
transform -1 0 23092 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0874_
timestamp 1649977179
transform 1 0 21712 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0875_
timestamp 1649977179
transform -1 0 26772 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0876_
timestamp 1649977179
transform 1 0 25576 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0877_
timestamp 1649977179
transform -1 0 25944 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0878_
timestamp 1649977179
transform 1 0 25392 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0879_
timestamp 1649977179
transform -1 0 30176 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0880_
timestamp 1649977179
transform 1 0 23276 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0881_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20516 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0882_
timestamp 1649977179
transform 1 0 21804 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _0883_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21712 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _0884_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 25024 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0885_
timestamp 1649977179
transform -1 0 36340 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0886_
timestamp 1649977179
transform 1 0 35236 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0887_
timestamp 1649977179
transform -1 0 36524 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0888_
timestamp 1649977179
transform 1 0 35328 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0889_
timestamp 1649977179
transform 1 0 36248 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0890_
timestamp 1649977179
transform -1 0 35880 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0891_
timestamp 1649977179
transform -1 0 36432 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0892_
timestamp 1649977179
transform -1 0 35972 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0893_
timestamp 1649977179
transform 1 0 35972 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0894_
timestamp 1649977179
transform -1 0 38640 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0895_
timestamp 1649977179
transform 1 0 37536 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0896_
timestamp 1649977179
transform 1 0 37720 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0897_
timestamp 1649977179
transform -1 0 22172 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _0898_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21804 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__o41a_2  _0899_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 22172 0 1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_1  _0900_
timestamp 1649977179
transform -1 0 37628 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0901_
timestamp 1649977179
transform -1 0 33488 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0902_
timestamp 1649977179
transform 1 0 33396 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0903_
timestamp 1649977179
transform -1 0 32660 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0904_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 35512 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0905_
timestamp 1649977179
transform 1 0 34316 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0906_
timestamp 1649977179
transform -1 0 38548 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0907_
timestamp 1649977179
transform 1 0 38088 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0908_
timestamp 1649977179
transform 1 0 37444 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0909_
timestamp 1649977179
transform 1 0 36340 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0910_
timestamp 1649977179
transform 1 0 35972 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0911_
timestamp 1649977179
transform -1 0 37260 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0912_
timestamp 1649977179
transform 1 0 37260 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0913_
timestamp 1649977179
transform -1 0 35696 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _0914_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 35052 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _0915_
timestamp 1649977179
transform -1 0 36616 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0916_
timestamp 1649977179
transform 1 0 36524 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0917_
timestamp 1649977179
transform -1 0 35328 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0918_
timestamp 1649977179
transform 1 0 34776 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0919_
timestamp 1649977179
transform 1 0 34684 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0920_
timestamp 1649977179
transform 1 0 38272 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0921_
timestamp 1649977179
transform 1 0 39008 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0922_
timestamp 1649977179
transform -1 0 39376 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0923_
timestamp 1649977179
transform 1 0 37996 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0924_
timestamp 1649977179
transform -1 0 37904 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0925_
timestamp 1649977179
transform -1 0 35420 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0926_
timestamp 1649977179
transform 1 0 34684 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0927_
timestamp 1649977179
transform -1 0 34224 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0928_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 31556 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0929_
timestamp 1649977179
transform -1 0 36708 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0930_
timestamp 1649977179
transform -1 0 36800 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0931_
timestamp 1649977179
transform 1 0 36892 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0932_
timestamp 1649977179
transform -1 0 38732 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0933_
timestamp 1649977179
transform 1 0 38272 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0934_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 37260 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0935_
timestamp 1649977179
transform -1 0 36524 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0936_
timestamp 1649977179
transform -1 0 38180 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0937_
timestamp 1649977179
transform -1 0 36708 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0938_
timestamp 1649977179
transform 1 0 32200 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0939_
timestamp 1649977179
transform -1 0 34224 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0940_
timestamp 1649977179
transform 1 0 34040 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0941_
timestamp 1649977179
transform -1 0 36340 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0942_
timestamp 1649977179
transform -1 0 37904 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0943_
timestamp 1649977179
transform -1 0 37812 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0944_
timestamp 1649977179
transform -1 0 40480 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0945_
timestamp 1649977179
transform -1 0 38180 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0946_
timestamp 1649977179
transform 1 0 39100 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0947_
timestamp 1649977179
transform 1 0 38272 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1649977179
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0949_
timestamp 1649977179
transform 1 0 38180 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0950_
timestamp 1649977179
transform -1 0 39284 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0951_
timestamp 1649977179
transform 1 0 38088 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0952_
timestamp 1649977179
transform 1 0 38916 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0953_
timestamp 1649977179
transform -1 0 36064 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0954_
timestamp 1649977179
transform 1 0 36064 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0955_
timestamp 1649977179
transform -1 0 35696 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _0956_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 33304 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _0957_
timestamp 1649977179
transform 1 0 32476 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _0958_
timestamp 1649977179
transform -1 0 41584 0 1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__a22oi_2  _0959_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 39100 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_2  _0960_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 40296 0 -1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0961_
timestamp 1649977179
transform -1 0 41952 0 -1 36992
box -38 -48 1234 592
use sky130_fd_sc_hd__o21bai_1  _0962_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 38548 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _0963_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 37904 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0964_
timestamp 1649977179
transform -1 0 38824 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0965_
timestamp 1649977179
transform 1 0 32752 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0966_
timestamp 1649977179
transform -1 0 40296 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0967_
timestamp 1649977179
transform 1 0 39284 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0968_
timestamp 1649977179
transform 1 0 39836 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0969_
timestamp 1649977179
transform 1 0 35696 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0970_
timestamp 1649977179
transform 1 0 35512 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0971_
timestamp 1649977179
transform -1 0 35880 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0972_
timestamp 1649977179
transform -1 0 34868 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0973_
timestamp 1649977179
transform -1 0 34316 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0974_
timestamp 1649977179
transform 1 0 35144 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0975_
timestamp 1649977179
transform -1 0 36984 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0976_
timestamp 1649977179
transform 1 0 37168 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0977_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 38180 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0978_
timestamp 1649977179
transform 1 0 40388 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0979_
timestamp 1649977179
transform 1 0 39836 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0980_
timestamp 1649977179
transform 1 0 37260 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0981_
timestamp 1649977179
transform 1 0 36156 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0982_
timestamp 1649977179
transform -1 0 39376 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0983_
timestamp 1649977179
transform 1 0 39836 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0984_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 40388 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _0985_
timestamp 1649977179
transform 1 0 39744 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0986_
timestamp 1649977179
transform 1 0 40480 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0987_
timestamp 1649977179
transform -1 0 40756 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0988_
timestamp 1649977179
transform -1 0 37536 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0989_
timestamp 1649977179
transform -1 0 36892 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0990_
timestamp 1649977179
transform -1 0 36432 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0991_
timestamp 1649977179
transform -1 0 39192 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0992_
timestamp 1649977179
transform -1 0 38916 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0993_
timestamp 1649977179
transform 1 0 37260 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0994_
timestamp 1649977179
transform -1 0 37352 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0995_
timestamp 1649977179
transform -1 0 33856 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0996_
timestamp 1649977179
transform 1 0 32660 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0997_
timestamp 1649977179
transform 1 0 33580 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0998_
timestamp 1649977179
transform -1 0 34224 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0999_
timestamp 1649977179
transform 1 0 34316 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1000_
timestamp 1649977179
transform -1 0 32292 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1001_
timestamp 1649977179
transform 1 0 32108 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1002_
timestamp 1649977179
transform 1 0 24748 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1003_
timestamp 1649977179
transform 1 0 32476 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1004_
timestamp 1649977179
transform 1 0 32844 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1005_
timestamp 1649977179
transform 1 0 33396 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1006_
timestamp 1649977179
transform -1 0 35880 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1007_
timestamp 1649977179
transform 1 0 34684 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1008_
timestamp 1649977179
transform -1 0 35972 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1009_
timestamp 1649977179
transform -1 0 35236 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1010_
timestamp 1649977179
transform 1 0 36340 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1011_
timestamp 1649977179
transform -1 0 39376 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1012_
timestamp 1649977179
transform -1 0 36156 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _1013_
timestamp 1649977179
transform -1 0 41492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1014_
timestamp 1649977179
transform 1 0 39836 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _1015_
timestamp 1649977179
transform 1 0 33488 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1016_
timestamp 1649977179
transform -1 0 35144 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1017_
timestamp 1649977179
transform -1 0 34500 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1018_
timestamp 1649977179
transform 1 0 33212 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1019_
timestamp 1649977179
transform -1 0 35052 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1020_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 33212 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1021_
timestamp 1649977179
transform -1 0 39468 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1022_
timestamp 1649977179
transform 1 0 38088 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1023_
timestamp 1649977179
transform 1 0 38732 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1024_
timestamp 1649977179
transform 1 0 35972 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1025_
timestamp 1649977179
transform -1 0 36340 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1026_
timestamp 1649977179
transform 1 0 32476 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1027_
timestamp 1649977179
transform -1 0 29440 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1028_
timestamp 1649977179
transform 1 0 33028 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1649977179
transform 1 0 35696 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1030_
timestamp 1649977179
transform 1 0 33120 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1031_
timestamp 1649977179
transform -1 0 34776 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1032_
timestamp 1649977179
transform 1 0 34684 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1033_
timestamp 1649977179
transform 1 0 34960 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1034_
timestamp 1649977179
transform -1 0 34684 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1035_
timestamp 1649977179
transform -1 0 35880 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1036_
timestamp 1649977179
transform -1 0 31188 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1037_
timestamp 1649977179
transform -1 0 30544 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1038_
timestamp 1649977179
transform 1 0 30084 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1039_
timestamp 1649977179
transform -1 0 38640 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1040_
timestamp 1649977179
transform -1 0 37812 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1041_
timestamp 1649977179
transform 1 0 37720 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1042_
timestamp 1649977179
transform 1 0 31004 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1043_
timestamp 1649977179
transform -1 0 34040 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1044_
timestamp 1649977179
transform 1 0 33672 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1045_
timestamp 1649977179
transform -1 0 33304 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1046_
timestamp 1649977179
transform 1 0 32476 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _1047_
timestamp 1649977179
transform -1 0 33764 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1048_
timestamp 1649977179
transform 1 0 26220 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1049_
timestamp 1649977179
transform 1 0 28704 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1050_
timestamp 1649977179
transform -1 0 29992 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1051_
timestamp 1649977179
transform -1 0 27968 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1052_
timestamp 1649977179
transform -1 0 28704 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1053_
timestamp 1649977179
transform 1 0 30912 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1054_
timestamp 1649977179
transform 1 0 31004 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1055_
timestamp 1649977179
transform 1 0 32108 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1056_
timestamp 1649977179
transform -1 0 32568 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1057_
timestamp 1649977179
transform 1 0 32844 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1058_
timestamp 1649977179
transform -1 0 33396 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _1059_
timestamp 1649977179
transform -1 0 33120 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__nor3_1  _1060_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 34224 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1061_
timestamp 1649977179
transform 1 0 34776 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1062_
timestamp 1649977179
transform 1 0 34592 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1063_
timestamp 1649977179
transform 1 0 33580 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1064_
timestamp 1649977179
transform -1 0 31832 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1065_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 28244 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1066_
timestamp 1649977179
transform 1 0 28336 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1067_
timestamp 1649977179
transform 1 0 28612 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1068_
timestamp 1649977179
transform 1 0 33764 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_1  _1069_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 35236 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1070_
timestamp 1649977179
transform -1 0 37720 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_4  _1071_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 37720 0 1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_1  _1072_
timestamp 1649977179
transform -1 0 31096 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1073_
timestamp 1649977179
transform -1 0 33120 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1074_
timestamp 1649977179
transform 1 0 31464 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1075_
timestamp 1649977179
transform 1 0 12328 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1076_
timestamp 1649977179
transform 1 0 12328 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1077_
timestamp 1649977179
transform -1 0 13248 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1078_
timestamp 1649977179
transform 1 0 15180 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1079_
timestamp 1649977179
transform 1 0 14812 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1080_
timestamp 1649977179
transform 1 0 15548 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1081_
timestamp 1649977179
transform 1 0 31188 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1082_
timestamp 1649977179
transform 1 0 31280 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1083_
timestamp 1649977179
transform 1 0 33488 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1084_
timestamp 1649977179
transform -1 0 33212 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1085_
timestamp 1649977179
transform -1 0 32660 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1086_
timestamp 1649977179
transform -1 0 32384 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1087_
timestamp 1649977179
transform 1 0 27232 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1088_
timestamp 1649977179
transform 1 0 28336 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1089_
timestamp 1649977179
transform 1 0 15732 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1090_
timestamp 1649977179
transform 1 0 15088 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1091_
timestamp 1649977179
transform -1 0 16468 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1092_
timestamp 1649977179
transform 1 0 29900 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1093_
timestamp 1649977179
transform -1 0 29900 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1094_
timestamp 1649977179
transform -1 0 30176 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1095_
timestamp 1649977179
transform -1 0 17848 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1096_
timestamp 1649977179
transform 1 0 18216 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1097_
timestamp 1649977179
transform 1 0 19228 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1098_
timestamp 1649977179
transform 1 0 27232 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1099_
timestamp 1649977179
transform 1 0 14812 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1100_
timestamp 1649977179
transform -1 0 14444 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1101_
timestamp 1649977179
transform 1 0 15640 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1102_
timestamp 1649977179
transform 1 0 16652 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1103_
timestamp 1649977179
transform -1 0 17020 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1104_
timestamp 1649977179
transform -1 0 17112 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1105_
timestamp 1649977179
transform -1 0 13984 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1106_
timestamp 1649977179
transform 1 0 14352 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1107_
timestamp 1649977179
transform 1 0 13156 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _1108_
timestamp 1649977179
transform -1 0 14444 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1109_
timestamp 1649977179
transform -1 0 13984 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1110_
timestamp 1649977179
transform -1 0 15272 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1111_
timestamp 1649977179
transform -1 0 16008 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1112_
timestamp 1649977179
transform -1 0 15732 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1113_
timestamp 1649977179
transform -1 0 33764 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1114_
timestamp 1649977179
transform -1 0 33212 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1115_
timestamp 1649977179
transform -1 0 32752 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1116_
timestamp 1649977179
transform 1 0 33396 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1117_
timestamp 1649977179
transform 1 0 32292 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _1118_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 32200 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1119_
timestamp 1649977179
transform 1 0 17572 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1120_
timestamp 1649977179
transform -1 0 16284 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1121_
timestamp 1649977179
transform 1 0 17848 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1122_
timestamp 1649977179
transform -1 0 28612 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1123_
timestamp 1649977179
transform -1 0 27508 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1124_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 27600 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1125_
timestamp 1649977179
transform -1 0 26496 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1126_
timestamp 1649977179
transform 1 0 25484 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1127_
timestamp 1649977179
transform -1 0 26772 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1128_
timestamp 1649977179
transform -1 0 13616 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1129_
timestamp 1649977179
transform -1 0 14536 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1130_
timestamp 1649977179
transform -1 0 13616 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1131_
timestamp 1649977179
transform -1 0 15456 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1132_
timestamp 1649977179
transform 1 0 14720 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1133_
timestamp 1649977179
transform 1 0 14996 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1134_
timestamp 1649977179
transform 1 0 11500 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1135_
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1136_
timestamp 1649977179
transform 1 0 10856 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1137_
timestamp 1649977179
transform -1 0 12696 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1138_
timestamp 1649977179
transform -1 0 13892 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1139_
timestamp 1649977179
transform 1 0 12972 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1140_
timestamp 1649977179
transform 1 0 14260 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1141_
timestamp 1649977179
transform -1 0 14536 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1142_
timestamp 1649977179
transform 1 0 14536 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1143_
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1144_
timestamp 1649977179
transform 1 0 16652 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1145_
timestamp 1649977179
transform -1 0 18400 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1146_
timestamp 1649977179
transform -1 0 27324 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1147_
timestamp 1649977179
transform 1 0 12512 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1148_
timestamp 1649977179
transform 1 0 13156 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1149_
timestamp 1649977179
transform 1 0 14076 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1150_
timestamp 1649977179
transform -1 0 14628 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1151_
timestamp 1649977179
transform 1 0 14260 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1152_
timestamp 1649977179
transform 1 0 23460 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1153_
timestamp 1649977179
transform -1 0 24932 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1154_
timestamp 1649977179
transform 1 0 25300 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1155_
timestamp 1649977179
transform 1 0 12604 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1156_
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1157_
timestamp 1649977179
transform 1 0 10764 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1158_
timestamp 1649977179
transform -1 0 12052 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1159_
timestamp 1649977179
transform 1 0 12512 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1160_
timestamp 1649977179
transform -1 0 12972 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1161_
timestamp 1649977179
transform -1 0 14628 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1162_
timestamp 1649977179
transform 1 0 13248 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1163_
timestamp 1649977179
transform -1 0 16468 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1164_
timestamp 1649977179
transform -1 0 14168 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1165_
timestamp 1649977179
transform -1 0 15456 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1166_
timestamp 1649977179
transform 1 0 15180 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1167_
timestamp 1649977179
transform -1 0 24932 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1168_
timestamp 1649977179
transform -1 0 24748 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1169_
timestamp 1649977179
transform 1 0 12696 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1170_
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1171_
timestamp 1649977179
transform -1 0 15824 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1172_
timestamp 1649977179
transform 1 0 11500 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1173_
timestamp 1649977179
transform -1 0 13156 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1174_
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1175_
timestamp 1649977179
transform 1 0 15916 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1176_
timestamp 1649977179
transform 1 0 16836 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1177_
timestamp 1649977179
transform -1 0 16468 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1178_
timestamp 1649977179
transform -1 0 17204 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1179_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _1180_
timestamp 1649977179
transform -1 0 16192 0 -1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__a21boi_1  _1181_
timestamp 1649977179
transform 1 0 15088 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1182_
timestamp 1649977179
transform 1 0 15456 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1183_
timestamp 1649977179
transform -1 0 24564 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1184_
timestamp 1649977179
transform 1 0 23184 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1185_
timestamp 1649977179
transform 1 0 23644 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1186_
timestamp 1649977179
transform -1 0 25024 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1187_
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1188_
timestamp 1649977179
transform 1 0 16468 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1189_
timestamp 1649977179
transform 1 0 17296 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1190_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15640 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1191_
timestamp 1649977179
transform -1 0 13708 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1192_
timestamp 1649977179
transform -1 0 15548 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1193_
timestamp 1649977179
transform -1 0 14628 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1194_
timestamp 1649977179
transform -1 0 19044 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1195_
timestamp 1649977179
transform 1 0 17664 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1196_
timestamp 1649977179
transform 1 0 24380 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1197_
timestamp 1649977179
transform -1 0 23920 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1198_
timestamp 1649977179
transform -1 0 23552 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1199_
timestamp 1649977179
transform 1 0 17388 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1200_
timestamp 1649977179
transform 1 0 19688 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1201_
timestamp 1649977179
transform 1 0 17204 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1202_
timestamp 1649977179
transform -1 0 18216 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1203_
timestamp 1649977179
transform -1 0 18768 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1204_
timestamp 1649977179
transform 1 0 17940 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1205_
timestamp 1649977179
transform -1 0 19320 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1206_
timestamp 1649977179
transform 1 0 17940 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1207_
timestamp 1649977179
transform -1 0 17756 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1208_
timestamp 1649977179
transform -1 0 17940 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1209_
timestamp 1649977179
transform 1 0 18032 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1210_
timestamp 1649977179
transform 1 0 17112 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1211_
timestamp 1649977179
transform 1 0 19228 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1212_
timestamp 1649977179
transform 1 0 15364 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1213_
timestamp 1649977179
transform 1 0 16652 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1214_
timestamp 1649977179
transform -1 0 15088 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1215_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16836 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1216_
timestamp 1649977179
transform -1 0 17112 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a311oi_2  _1217_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15364 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__a21bo_1  _1218_
timestamp 1649977179
transform 1 0 18584 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1219_
timestamp 1649977179
transform -1 0 19872 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1220_
timestamp 1649977179
transform -1 0 19320 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1221_
timestamp 1649977179
transform -1 0 23920 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1222_
timestamp 1649977179
transform -1 0 19964 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1223_
timestamp 1649977179
transform 1 0 19780 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1224_
timestamp 1649977179
transform 1 0 20332 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1225_
timestamp 1649977179
transform -1 0 19504 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1226_
timestamp 1649977179
transform -1 0 17940 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1227_
timestamp 1649977179
transform 1 0 20884 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1228_
timestamp 1649977179
transform 1 0 20056 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1229_
timestamp 1649977179
transform 1 0 22724 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1230_
timestamp 1649977179
transform 1 0 22908 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1231_
timestamp 1649977179
transform 1 0 17572 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1232_
timestamp 1649977179
transform -1 0 18124 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1233_
timestamp 1649977179
transform 1 0 17848 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1234_
timestamp 1649977179
transform 1 0 18860 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1235_
timestamp 1649977179
transform -1 0 20700 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1236_
timestamp 1649977179
transform -1 0 19596 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1237_
timestamp 1649977179
transform -1 0 19320 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1238_
timestamp 1649977179
transform -1 0 18584 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1239_
timestamp 1649977179
transform 1 0 18308 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1240_
timestamp 1649977179
transform -1 0 20056 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1241_
timestamp 1649977179
transform -1 0 19964 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1242_
timestamp 1649977179
transform -1 0 19780 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1243_
timestamp 1649977179
transform 1 0 19780 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1244_
timestamp 1649977179
transform -1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _1245_
timestamp 1649977179
transform -1 0 22448 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _1246_
timestamp 1649977179
transform 1 0 21804 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1247_
timestamp 1649977179
transform 1 0 27692 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1248_
timestamp 1649977179
transform -1 0 20700 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1249_
timestamp 1649977179
transform 1 0 20332 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1250_
timestamp 1649977179
transform -1 0 20700 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1251_
timestamp 1649977179
transform -1 0 20608 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1252_
timestamp 1649977179
transform -1 0 20976 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1253_
timestamp 1649977179
transform -1 0 21252 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1254_
timestamp 1649977179
transform -1 0 23276 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1255_
timestamp 1649977179
transform 1 0 23368 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1256_
timestamp 1649977179
transform -1 0 20608 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1257_
timestamp 1649977179
transform -1 0 20332 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1258_
timestamp 1649977179
transform 1 0 19688 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1259_
timestamp 1649977179
transform -1 0 19872 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1260_
timestamp 1649977179
transform 1 0 19504 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1261_
timestamp 1649977179
transform 1 0 20424 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1262_
timestamp 1649977179
transform -1 0 20056 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1263_
timestamp 1649977179
transform 1 0 20700 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1264_
timestamp 1649977179
transform 1 0 19780 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _1265_
timestamp 1649977179
transform -1 0 19320 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1266_
timestamp 1649977179
transform 1 0 19688 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1267_
timestamp 1649977179
transform 1 0 20516 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1268_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 23000 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1269_
timestamp 1649977179
transform -1 0 22356 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1270_
timestamp 1649977179
transform 1 0 20792 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1271_
timestamp 1649977179
transform -1 0 20700 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1272_
timestamp 1649977179
transform 1 0 19044 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _1273_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18400 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1274_
timestamp 1649977179
transform 1 0 22448 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1275_
timestamp 1649977179
transform -1 0 22080 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1276_
timestamp 1649977179
transform -1 0 22080 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _1277_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20516 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1278_
timestamp 1649977179
transform 1 0 20608 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1279_
timestamp 1649977179
transform 1 0 21160 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1280_
timestamp 1649977179
transform -1 0 21896 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1281_
timestamp 1649977179
transform 1 0 21436 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1282_
timestamp 1649977179
transform 1 0 21528 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1283_
timestamp 1649977179
transform 1 0 22448 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1284_
timestamp 1649977179
transform 1 0 22356 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1285_
timestamp 1649977179
transform 1 0 23276 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1286_
timestamp 1649977179
transform 1 0 18216 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1287_
timestamp 1649977179
transform 1 0 19412 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1288_
timestamp 1649977179
transform 1 0 18308 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1289_
timestamp 1649977179
transform -1 0 20976 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _1290_
timestamp 1649977179
transform 1 0 21804 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1291_
timestamp 1649977179
transform -1 0 21988 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1292_
timestamp 1649977179
transform 1 0 22080 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1293_
timestamp 1649977179
transform 1 0 22540 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1294_
timestamp 1649977179
transform -1 0 23828 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_2  _1295_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22356 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _1296_
timestamp 1649977179
transform -1 0 25392 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1297_
timestamp 1649977179
transform 1 0 25116 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1298_
timestamp 1649977179
transform -1 0 26036 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1299_
timestamp 1649977179
transform 1 0 20516 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  _1300_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20792 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1301_
timestamp 1649977179
transform -1 0 20148 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1302_
timestamp 1649977179
transform -1 0 21344 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1303_
timestamp 1649977179
transform 1 0 20608 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1304_
timestamp 1649977179
transform -1 0 22632 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1305_
timestamp 1649977179
transform 1 0 20608 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1306_
timestamp 1649977179
transform 1 0 20424 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1307_
timestamp 1649977179
transform -1 0 24656 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1308_
timestamp 1649977179
transform 1 0 21988 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1309_
timestamp 1649977179
transform -1 0 21344 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1310_
timestamp 1649977179
transform -1 0 22356 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1311_
timestamp 1649977179
transform 1 0 23000 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1312_
timestamp 1649977179
transform 1 0 22172 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1313_
timestamp 1649977179
transform 1 0 22632 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1314_
timestamp 1649977179
transform -1 0 23828 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1315_
timestamp 1649977179
transform 1 0 23736 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1316_
timestamp 1649977179
transform 1 0 23828 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1317_
timestamp 1649977179
transform 1 0 25576 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1318_
timestamp 1649977179
transform -1 0 22908 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1319_
timestamp 1649977179
transform 1 0 21620 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1320_
timestamp 1649977179
transform 1 0 21712 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1321_
timestamp 1649977179
transform 1 0 23276 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1322_
timestamp 1649977179
transform 1 0 22632 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1323_
timestamp 1649977179
transform 1 0 24196 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1324_
timestamp 1649977179
transform -1 0 25208 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1325_
timestamp 1649977179
transform -1 0 23092 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1326_
timestamp 1649977179
transform -1 0 25024 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1327_
timestamp 1649977179
transform 1 0 24656 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1328_
timestamp 1649977179
transform -1 0 26036 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1329_
timestamp 1649977179
transform -1 0 25208 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1330_
timestamp 1649977179
transform -1 0 24472 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _1331_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 24748 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1332_
timestamp 1649977179
transform 1 0 23460 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1333_
timestamp 1649977179
transform -1 0 23092 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1334_
timestamp 1649977179
transform 1 0 23552 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1335_
timestamp 1649977179
transform 1 0 21528 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1336_
timestamp 1649977179
transform 1 0 22816 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1337_
timestamp 1649977179
transform 1 0 22816 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1338_
timestamp 1649977179
transform 1 0 24472 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1339_
timestamp 1649977179
transform -1 0 25392 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1340_
timestamp 1649977179
transform 1 0 24932 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1341_
timestamp 1649977179
transform 1 0 25944 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1342_
timestamp 1649977179
transform 1 0 25208 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1343_
timestamp 1649977179
transform -1 0 26404 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1344_
timestamp 1649977179
transform 1 0 25024 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1345_
timestamp 1649977179
transform -1 0 25760 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1346_
timestamp 1649977179
transform 1 0 26128 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1347_
timestamp 1649977179
transform -1 0 25576 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1348_
timestamp 1649977179
transform -1 0 26220 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1349_
timestamp 1649977179
transform 1 0 25576 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1350_
timestamp 1649977179
transform 1 0 25392 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1351_
timestamp 1649977179
transform 1 0 26772 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1352_
timestamp 1649977179
transform -1 0 23184 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1353_
timestamp 1649977179
transform 1 0 25852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1354_
timestamp 1649977179
transform -1 0 25392 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1355_
timestamp 1649977179
transform -1 0 24288 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1356_
timestamp 1649977179
transform 1 0 24840 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1357_
timestamp 1649977179
transform 1 0 25668 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1358_
timestamp 1649977179
transform 1 0 26036 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1359_
timestamp 1649977179
transform -1 0 26312 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1360_
timestamp 1649977179
transform 1 0 26772 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1361_
timestamp 1649977179
transform 1 0 25760 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1362_
timestamp 1649977179
transform 1 0 26772 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1363_
timestamp 1649977179
transform -1 0 25024 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1364_
timestamp 1649977179
transform -1 0 25760 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _1365_
timestamp 1649977179
transform -1 0 27508 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1366_
timestamp 1649977179
transform -1 0 28612 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1367_
timestamp 1649977179
transform 1 0 27508 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1368_
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1369_
timestamp 1649977179
transform -1 0 27508 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _1370_
timestamp 1649977179
transform 1 0 27324 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1371_
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1372_
timestamp 1649977179
transform 1 0 23736 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1373_
timestamp 1649977179
transform -1 0 24840 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1374_
timestamp 1649977179
transform -1 0 25484 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1375_
timestamp 1649977179
transform 1 0 24656 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1376_
timestamp 1649977179
transform 1 0 24656 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1377_
timestamp 1649977179
transform -1 0 27692 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1378_
timestamp 1649977179
transform 1 0 27692 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1379_
timestamp 1649977179
transform -1 0 27968 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1380_
timestamp 1649977179
transform 1 0 27508 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1381_
timestamp 1649977179
transform -1 0 24932 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1382_
timestamp 1649977179
transform 1 0 23184 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1383_
timestamp 1649977179
transform 1 0 22448 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1384_
timestamp 1649977179
transform 1 0 23276 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _1385_
timestamp 1649977179
transform -1 0 25208 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1386_
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1387_
timestamp 1649977179
transform 1 0 26772 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1388_
timestamp 1649977179
transform 1 0 28244 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1389_
timestamp 1649977179
transform -1 0 26956 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1390_
timestamp 1649977179
transform 1 0 27324 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1391_
timestamp 1649977179
transform 1 0 27876 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1392_
timestamp 1649977179
transform -1 0 27600 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1393_
timestamp 1649977179
transform -1 0 28060 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1394_
timestamp 1649977179
transform 1 0 27600 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1395_
timestamp 1649977179
transform -1 0 27968 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1396_
timestamp 1649977179
transform 1 0 27968 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1397_
timestamp 1649977179
transform 1 0 30360 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1398_
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1399_
timestamp 1649977179
transform -1 0 29992 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1400_
timestamp 1649977179
transform 1 0 28336 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1401_
timestamp 1649977179
transform -1 0 29072 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _1402_
timestamp 1649977179
transform -1 0 29164 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1403_
timestamp 1649977179
transform -1 0 28244 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1404_
timestamp 1649977179
transform 1 0 27140 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1405_
timestamp 1649977179
transform -1 0 28336 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1406_
timestamp 1649977179
transform 1 0 24564 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1407_
timestamp 1649977179
transform 1 0 27048 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1408_
timestamp 1649977179
transform 1 0 27416 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1409_
timestamp 1649977179
transform -1 0 27600 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1410_
timestamp 1649977179
transform -1 0 28336 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1411_
timestamp 1649977179
transform -1 0 26404 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1412_
timestamp 1649977179
transform -1 0 27324 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _1413_
timestamp 1649977179
transform 1 0 27876 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1414_
timestamp 1649977179
transform -1 0 28428 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1415_
timestamp 1649977179
transform -1 0 29072 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1416_
timestamp 1649977179
transform -1 0 29992 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1417_
timestamp 1649977179
transform 1 0 28704 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _1418_
timestamp 1649977179
transform 1 0 28428 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1419_
timestamp 1649977179
transform -1 0 28796 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1420_
timestamp 1649977179
transform 1 0 28428 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1421_
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1422_
timestamp 1649977179
transform -1 0 31280 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1423_
timestamp 1649977179
transform -1 0 31556 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1424_
timestamp 1649977179
transform 1 0 30268 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1425_
timestamp 1649977179
transform 1 0 26680 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1426_
timestamp 1649977179
transform 1 0 27324 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1427_
timestamp 1649977179
transform 1 0 29716 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1428_
timestamp 1649977179
transform -1 0 30728 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1429_
timestamp 1649977179
transform 1 0 30176 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1430_
timestamp 1649977179
transform 1 0 30268 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1431_
timestamp 1649977179
transform -1 0 29900 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1432_
timestamp 1649977179
transform 1 0 29532 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1433_
timestamp 1649977179
transform -1 0 31372 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1434_
timestamp 1649977179
transform 1 0 31188 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1435_
timestamp 1649977179
transform -1 0 31280 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1436_
timestamp 1649977179
transform -1 0 31188 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1437_
timestamp 1649977179
transform -1 0 30820 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _1438_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 29532 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1439_
timestamp 1649977179
transform -1 0 30176 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1440_
timestamp 1649977179
transform -1 0 31004 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1441_
timestamp 1649977179
transform 1 0 29808 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1442_
timestamp 1649977179
transform 1 0 29164 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1443_
timestamp 1649977179
transform -1 0 32016 0 1 39168
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1444_
timestamp 1649977179
transform -1 0 30728 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1445_
timestamp 1649977179
transform 1 0 30176 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1446_
timestamp 1649977179
transform -1 0 31004 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1447_
timestamp 1649977179
transform -1 0 31096 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1448_
timestamp 1649977179
transform -1 0 29716 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1449_
timestamp 1649977179
transform -1 0 30544 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1450_
timestamp 1649977179
transform 1 0 28244 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1451_
timestamp 1649977179
transform 1 0 29256 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1452_
timestamp 1649977179
transform 1 0 30084 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1453_
timestamp 1649977179
transform -1 0 31280 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1454_
timestamp 1649977179
transform 1 0 30268 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1455_
timestamp 1649977179
transform 1 0 30360 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1456_
timestamp 1649977179
transform 1 0 15180 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1457_
timestamp 1649977179
transform 1 0 16652 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1458_
timestamp 1649977179
transform 1 0 15548 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1459_
timestamp 1649977179
transform 1 0 17940 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1460_
timestamp 1649977179
transform -1 0 19044 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1461_
timestamp 1649977179
transform -1 0 19504 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1462_
timestamp 1649977179
transform -1 0 18584 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1463_
timestamp 1649977179
transform -1 0 18768 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1464_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 33672 0 -1 43520
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1465_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 29532 0 1 46784
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1466_
timestamp 1649977179
transform -1 0 29992 0 -1 45696
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1467_
timestamp 1649977179
transform -1 0 33672 0 -1 44608
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1468_
timestamp 1649977179
transform 1 0 27324 0 1 42432
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1469_
timestamp 1649977179
transform 1 0 32108 0 1 46784
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1470_
timestamp 1649977179
transform 1 0 32108 0 -1 46784
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1471_
timestamp 1649977179
transform 1 0 29532 0 1 40256
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1472_
timestamp 1649977179
transform 1 0 27508 0 1 40256
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1473_
timestamp 1649977179
transform -1 0 28612 0 -1 42432
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1474_
timestamp 1649977179
transform 1 0 27508 0 1 45696
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1475_
timestamp 1649977179
transform 1 0 27324 0 1 43520
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1476_
timestamp 1649977179
transform 1 0 27048 0 1 44608
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1477_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 25024 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1478_
timestamp 1649977179
transform 1 0 28336 0 -1 46784
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1479_
timestamp 1649977179
transform 1 0 29532 0 1 41344
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1480_
timestamp 1649977179
transform -1 0 26496 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1481_
timestamp 1649977179
transform 1 0 32108 0 1 45696
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1482_
timestamp 1649977179
transform -1 0 31280 0 1 44608
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1483_
timestamp 1649977179
transform 1 0 28980 0 -1 44608
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1484_
timestamp 1649977179
transform 1 0 34040 0 -1 43520
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1485_
timestamp 1649977179
transform -1 0 33396 0 1 42432
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1486_
timestamp 1649977179
transform 1 0 24932 0 -1 46784
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1487_
timestamp 1649977179
transform -1 0 28612 0 -1 44608
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1488_
timestamp 1649977179
transform 1 0 29992 0 1 45696
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1489_
timestamp 1649977179
transform 1 0 34684 0 1 46784
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1490_
timestamp 1649977179
transform 1 0 29532 0 1 42432
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1491_
timestamp 1649977179
transform 1 0 28980 0 -1 42432
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1492_
timestamp 1649977179
transform 1 0 32108 0 -1 41344
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1493_
timestamp 1649977179
transform 1 0 32108 0 -1 42432
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1494_
timestamp 1649977179
transform 1 0 25576 0 1 45696
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1495_
timestamp 1649977179
transform -1 0 33580 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 30452 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1649977179
transform -1 0 27876 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1649977179
transform -1 0 29072 0 1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1649977179
transform -1 0 30452 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1649977179
transform 1 0 31188 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  input1 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 48208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform 1 0 47932 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1649977179
transform -1 0 48208 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 1649977179
transform 1 0 1748 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input5
timestamp 1649977179
transform 1 0 43884 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 1649977179
transform 1 0 1380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1649977179
transform -1 0 48208 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input8
timestamp 1649977179
transform 1 0 36156 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input9
timestamp 1649977179
transform 1 0 1748 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1649977179
transform 1 0 1748 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1649977179
transform 1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1649977179
transform 1 0 1748 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input13
timestamp 1649977179
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1649977179
transform 1 0 1748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1649977179
transform 1 0 1748 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1649977179
transform -1 0 48208 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1649977179
transform -1 0 23644 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1649977179
transform 1 0 42412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1649977179
transform 1 0 1748 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1649977179
transform 1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1649977179
transform 1 0 1748 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1649977179
transform -1 0 28796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1649977179
transform 1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input24
timestamp 1649977179
transform -1 0 48208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 48208 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform -1 0 31648 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1649977179
transform 1 0 17480 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1649977179
transform -1 0 48208 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input30
timestamp 1649977179
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input31
timestamp 1649977179
transform 1 0 1748 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1649977179
transform -1 0 48208 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input33
timestamp 1649977179
transform 1 0 19412 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1649977179
transform -1 0 48208 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1649977179
transform -1 0 48208 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input36
timestamp 1649977179
transform 1 0 20792 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input37
timestamp 1649977179
transform 1 0 40020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input38
timestamp 1649977179
transform -1 0 48208 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1649977179
transform 1 0 7820 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1649977179
transform 1 0 1748 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1649977179
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1649977179
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp 1649977179
transform 1 0 30360 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1649977179
transform 1 0 9752 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1649977179
transform 1 0 26956 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1649977179
transform 1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp 1649977179
transform -1 0 2300 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1649977179
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1649977179
transform -1 0 45724 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1649977179
transform -1 0 35420 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1649977179
transform 1 0 22632 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1649977179
transform -1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1649977179
transform -1 0 48208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1649977179
transform 1 0 2668 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1649977179
transform -1 0 48208 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1649977179
transform 1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1649977179
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1649977179
transform 1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input60
timestamp 1649977179
transform -1 0 48208 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input62
timestamp 1649977179
transform -1 0 41032 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1649977179
transform 1 0 38732 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1649977179
transform -1 0 4232 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1649977179
transform 1 0 11868 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input66
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input67
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input68
timestamp 1649977179
transform 1 0 1380 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input69
timestamp 1649977179
transform -1 0 48208 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform 1 0 13248 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform -1 0 32660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform -1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform 1 0 47840 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform 1 0 47748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform 1 0 47840 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform 1 0 37260 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform 1 0 14904 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform 1 0 46736 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform 1 0 47840 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform 1 0 46460 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform 1 0 27140 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform -1 0 1748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform 1 0 47840 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform -1 0 1748 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform -1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform 1 0 34040 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform -1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform 1 0 42596 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform -1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform -1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform -1 0 15272 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform 1 0 45816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform 1 0 47840 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform 1 0 47840 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform -1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform -1 0 1748 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform 1 0 47840 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform -1 0 6716 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform 1 0 47840 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform 1 0 47840 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  repeater102
timestamp 1649977179
transform -1 0 27508 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  repeater103
timestamp 1649977179
transform 1 0 29348 0 -1 38080
box -38 -48 406 592
<< labels >>
flabel metal3 s 49200 7488 50000 7608 0 FreeSans 480 0 0 0 alu_branch
port 0 nsew signal input
flabel metal3 s 49200 42168 50000 42288 0 FreeSans 480 0 0 0 branch
port 1 nsew signal input
flabel metal2 s 28998 49200 29054 50000 0 FreeSans 224 90 0 0 clk
port 2 nsew signal input
flabel metal3 s 49200 48288 50000 48408 0 FreeSans 480 0 0 0 immediate[0]
port 3 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 immediate[10]
port 4 nsew signal input
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 immediate[11]
port 5 nsew signal input
flabel metal3 s 0 46248 800 46368 0 FreeSans 480 0 0 0 immediate[12]
port 6 nsew signal input
flabel metal2 s 48318 49200 48374 50000 0 FreeSans 224 90 0 0 immediate[13]
port 7 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 immediate[14]
port 8 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 immediate[15]
port 9 nsew signal input
flabel metal3 s 0 38088 800 38208 0 FreeSans 480 0 0 0 immediate[16]
port 10 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 immediate[17]
port 11 nsew signal input
flabel metal3 s 0 48288 800 48408 0 FreeSans 480 0 0 0 immediate[18]
port 12 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 immediate[19]
port 13 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 immediate[1]
port 14 nsew signal input
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 immediate[20]
port 15 nsew signal input
flabel metal3 s 49200 36048 50000 36168 0 FreeSans 480 0 0 0 immediate[21]
port 16 nsew signal input
flabel metal2 s 23202 49200 23258 50000 0 FreeSans 224 90 0 0 immediate[22]
port 17 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 immediate[23]
port 18 nsew signal input
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 immediate[24]
port 19 nsew signal input
flabel metal3 s 0 40128 800 40248 0 FreeSans 480 0 0 0 immediate[25]
port 20 nsew signal input
flabel metal3 s 0 34008 800 34128 0 FreeSans 480 0 0 0 immediate[26]
port 21 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 immediate[27]
port 22 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 immediate[28]
port 23 nsew signal input
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 immediate[29]
port 24 nsew signal input
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 immediate[2]
port 25 nsew signal input
flabel metal3 s 49200 25848 50000 25968 0 FreeSans 480 0 0 0 immediate[30]
port 26 nsew signal input
flabel metal2 s 30930 49200 30986 50000 0 FreeSans 224 90 0 0 immediate[31]
port 27 nsew signal input
flabel metal2 s 17406 49200 17462 50000 0 FreeSans 224 90 0 0 immediate[3]
port 28 nsew signal input
flabel metal3 s 49200 46248 50000 46368 0 FreeSans 480 0 0 0 immediate[4]
port 29 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 immediate[5]
port 30 nsew signal input
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 immediate[6]
port 31 nsew signal input
flabel metal3 s 49200 44208 50000 44328 0 FreeSans 480 0 0 0 immediate[7]
port 32 nsew signal input
flabel metal2 s 19338 49200 19394 50000 0 FreeSans 224 90 0 0 immediate[8]
port 33 nsew signal input
flabel metal3 s 49200 11568 50000 11688 0 FreeSans 480 0 0 0 immediate[9]
port 34 nsew signal input
flabel metal3 s 49200 15648 50000 15768 0 FreeSans 480 0 0 0 jump_jal
port 35 nsew signal input
flabel metal2 s 21270 49200 21326 50000 0 FreeSans 224 90 0 0 jump_jalr
port 36 nsew signal input
flabel metal2 s 13542 49200 13598 50000 0 FreeSans 224 90 0 0 pc_out[0]
port 37 nsew signal tristate
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 pc_out[10]
port 38 nsew signal tristate
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 pc_out[11]
port 39 nsew signal tristate
flabel metal3 s 49200 38088 50000 38208 0 FreeSans 480 0 0 0 pc_out[12]
port 40 nsew signal tristate
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 pc_out[13]
port 41 nsew signal tristate
flabel metal3 s 49200 19728 50000 19848 0 FreeSans 480 0 0 0 pc_out[14]
port 42 nsew signal tristate
flabel metal2 s 36726 49200 36782 50000 0 FreeSans 224 90 0 0 pc_out[15]
port 43 nsew signal tristate
flabel metal2 s 15474 49200 15530 50000 0 FreeSans 224 90 0 0 pc_out[16]
port 44 nsew signal tristate
flabel metal3 s 49200 1368 50000 1488 0 FreeSans 480 0 0 0 pc_out[17]
port 45 nsew signal tristate
flabel metal3 s 49200 40128 50000 40248 0 FreeSans 480 0 0 0 pc_out[18]
port 46 nsew signal tristate
flabel metal2 s 46386 49200 46442 50000 0 FreeSans 224 90 0 0 pc_out[19]
port 47 nsew signal tristate
flabel metal2 s 27066 49200 27122 50000 0 FreeSans 224 90 0 0 pc_out[1]
port 48 nsew signal tristate
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 pc_out[20]
port 49 nsew signal tristate
flabel metal3 s 49200 9528 50000 9648 0 FreeSans 480 0 0 0 pc_out[21]
port 50 nsew signal tristate
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 pc_out[22]
port 51 nsew signal tristate
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 pc_out[23]
port 52 nsew signal tristate
flabel metal2 s 32862 49200 32918 50000 0 FreeSans 224 90 0 0 pc_out[24]
port 53 nsew signal tristate
flabel metal3 s 0 36048 800 36168 0 FreeSans 480 0 0 0 pc_out[25]
port 54 nsew signal tristate
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 pc_out[26]
port 55 nsew signal tristate
flabel metal2 s 42522 49200 42578 50000 0 FreeSans 224 90 0 0 pc_out[27]
port 56 nsew signal tristate
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 pc_out[28]
port 57 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 pc_out[29]
port 58 nsew signal tristate
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 pc_out[2]
port 59 nsew signal tristate
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 pc_out[30]
port 60 nsew signal tristate
flabel metal3 s 49200 21768 50000 21888 0 FreeSans 480 0 0 0 pc_out[31]
port 61 nsew signal tristate
flabel metal3 s 49200 13608 50000 13728 0 FreeSans 480 0 0 0 pc_out[3]
port 62 nsew signal tristate
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 pc_out[4]
port 63 nsew signal tristate
flabel metal3 s 0 42168 800 42288 0 FreeSans 480 0 0 0 pc_out[5]
port 64 nsew signal tristate
flabel metal3 s 49200 3408 50000 3528 0 FreeSans 480 0 0 0 pc_out[6]
port 65 nsew signal tristate
flabel metal2 s 5814 49200 5870 50000 0 FreeSans 224 90 0 0 pc_out[7]
port 66 nsew signal tristate
flabel metal3 s 49200 17688 50000 17808 0 FreeSans 480 0 0 0 pc_out[8]
port 67 nsew signal tristate
flabel metal3 s 49200 31968 50000 32088 0 FreeSans 480 0 0 0 pc_out[9]
port 68 nsew signal tristate
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 rs1_data[0]
port 69 nsew signal input
flabel metal3 s 49200 34008 50000 34128 0 FreeSans 480 0 0 0 rs1_data[10]
port 70 nsew signal input
flabel metal2 s 7746 49200 7802 50000 0 FreeSans 224 90 0 0 rs1_data[11]
port 71 nsew signal input
flabel metal3 s 0 29928 800 30048 0 FreeSans 480 0 0 0 rs1_data[12]
port 72 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 rs1_data[13]
port 73 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 rs1_data[14]
port 74 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 rs1_data[15]
port 75 nsew signal input
flabel metal2 s 9678 49200 9734 50000 0 FreeSans 224 90 0 0 rs1_data[16]
port 76 nsew signal input
flabel metal2 s 25134 49200 25190 50000 0 FreeSans 224 90 0 0 rs1_data[17]
port 77 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 rs1_data[18]
port 78 nsew signal input
flabel metal2 s 18 49200 74 50000 0 FreeSans 224 90 0 0 rs1_data[19]
port 79 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 rs1_data[1]
port 80 nsew signal input
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 rs1_data[20]
port 81 nsew signal input
flabel metal2 s 44454 49200 44510 50000 0 FreeSans 224 90 0 0 rs1_data[21]
port 82 nsew signal input
flabel metal2 s 34794 49200 34850 50000 0 FreeSans 224 90 0 0 rs1_data[22]
port 83 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 rs1_data[23]
port 84 nsew signal input
flabel metal2 s 49606 49200 49662 50000 0 FreeSans 224 90 0 0 rs1_data[24]
port 85 nsew signal input
flabel metal3 s 49200 5448 50000 5568 0 FreeSans 480 0 0 0 rs1_data[25]
port 86 nsew signal input
flabel metal2 s 1950 49200 2006 50000 0 FreeSans 224 90 0 0 rs1_data[26]
port 87 nsew signal input
flabel metal3 s 49200 27888 50000 28008 0 FreeSans 480 0 0 0 rs1_data[27]
port 88 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 rs1_data[28]
port 89 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 rs1_data[29]
port 90 nsew signal input
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 rs1_data[2]
port 91 nsew signal input
flabel metal3 s 49200 29928 50000 30048 0 FreeSans 480 0 0 0 rs1_data[30]
port 92 nsew signal input
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 rs1_data[31]
port 93 nsew signal input
flabel metal2 s 40590 49200 40646 50000 0 FreeSans 224 90 0 0 rs1_data[3]
port 94 nsew signal input
flabel metal2 s 38658 49200 38714 50000 0 FreeSans 224 90 0 0 rs1_data[4]
port 95 nsew signal input
flabel metal2 s 3882 49200 3938 50000 0 FreeSans 224 90 0 0 rs1_data[5]
port 96 nsew signal input
flabel metal2 s 11610 49200 11666 50000 0 FreeSans 224 90 0 0 rs1_data[6]
port 97 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 rs1_data[7]
port 98 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 rs1_data[8]
port 99 nsew signal input
flabel metal3 s 0 44208 800 44328 0 FreeSans 480 0 0 0 rs1_data[9]
port 100 nsew signal input
flabel metal3 s 49200 23808 50000 23928 0 FreeSans 480 0 0 0 rst_n
port 101 nsew signal input
flabel metal4 s 4208 2128 4528 47376 0 FreeSans 1920 90 0 0 vccd1
port 102 nsew power bidirectional
flabel metal4 s 34928 2128 35248 47376 0 FreeSans 1920 90 0 0 vccd1
port 102 nsew power bidirectional
flabel metal4 s 19568 2128 19888 47376 0 FreeSans 1920 90 0 0 vssd1
port 103 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
