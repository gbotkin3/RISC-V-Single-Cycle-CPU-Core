magic
tech sky130B
magscale 1 2
timestamp 1663796782
<< obsli1 >>
rect 1104 2159 562856 681649
<< obsm1 >>
rect 14 2128 562856 681680
<< metal2 >>
rect 18 683200 74 684000
rect 6458 683200 6514 684000
rect 12898 683200 12954 684000
rect 19338 683200 19394 684000
rect 25778 683200 25834 684000
rect 31574 683200 31630 684000
rect 38014 683200 38070 684000
rect 44454 683200 44510 684000
rect 50894 683200 50950 684000
rect 56690 683200 56746 684000
rect 63130 683200 63186 684000
rect 69570 683200 69626 684000
rect 76010 683200 76066 684000
rect 82450 683200 82506 684000
rect 88246 683200 88302 684000
rect 94686 683200 94742 684000
rect 101126 683200 101182 684000
rect 107566 683200 107622 684000
rect 113362 683200 113418 684000
rect 119802 683200 119858 684000
rect 126242 683200 126298 684000
rect 132682 683200 132738 684000
rect 139122 683200 139178 684000
rect 144918 683200 144974 684000
rect 151358 683200 151414 684000
rect 157798 683200 157854 684000
rect 164238 683200 164294 684000
rect 170034 683200 170090 684000
rect 176474 683200 176530 684000
rect 182914 683200 182970 684000
rect 189354 683200 189410 684000
rect 195794 683200 195850 684000
rect 201590 683200 201646 684000
rect 208030 683200 208086 684000
rect 214470 683200 214526 684000
rect 220910 683200 220966 684000
rect 226706 683200 226762 684000
rect 233146 683200 233202 684000
rect 239586 683200 239642 684000
rect 246026 683200 246082 684000
rect 252466 683200 252522 684000
rect 258262 683200 258318 684000
rect 264702 683200 264758 684000
rect 271142 683200 271198 684000
rect 277582 683200 277638 684000
rect 283378 683200 283434 684000
rect 289818 683200 289874 684000
rect 296258 683200 296314 684000
rect 302698 683200 302754 684000
rect 309138 683200 309194 684000
rect 314934 683200 314990 684000
rect 321374 683200 321430 684000
rect 327814 683200 327870 684000
rect 334254 683200 334310 684000
rect 340050 683200 340106 684000
rect 346490 683200 346546 684000
rect 352930 683200 352986 684000
rect 359370 683200 359426 684000
rect 365810 683200 365866 684000
rect 371606 683200 371662 684000
rect 378046 683200 378102 684000
rect 384486 683200 384542 684000
rect 390926 683200 390982 684000
rect 396722 683200 396778 684000
rect 403162 683200 403218 684000
rect 409602 683200 409658 684000
rect 416042 683200 416098 684000
rect 422482 683200 422538 684000
rect 428278 683200 428334 684000
rect 434718 683200 434774 684000
rect 441158 683200 441214 684000
rect 447598 683200 447654 684000
rect 453394 683200 453450 684000
rect 459834 683200 459890 684000
rect 466274 683200 466330 684000
rect 472714 683200 472770 684000
rect 479154 683200 479210 684000
rect 484950 683200 485006 684000
rect 491390 683200 491446 684000
rect 497830 683200 497886 684000
rect 504270 683200 504326 684000
rect 510066 683200 510122 684000
rect 516506 683200 516562 684000
rect 522946 683200 523002 684000
rect 529386 683200 529442 684000
rect 535826 683200 535882 684000
rect 541622 683200 541678 684000
rect 548062 683200 548118 684000
rect 554502 683200 554558 684000
rect 560942 683200 560998 684000
rect 18 0 74 800
rect 5814 0 5870 800
rect 12254 0 12310 800
rect 18694 0 18750 800
rect 25134 0 25190 800
rect 30930 0 30986 800
rect 37370 0 37426 800
rect 43810 0 43866 800
rect 50250 0 50306 800
rect 56046 0 56102 800
rect 62486 0 62542 800
rect 68926 0 68982 800
rect 75366 0 75422 800
rect 81806 0 81862 800
rect 87602 0 87658 800
rect 94042 0 94098 800
rect 100482 0 100538 800
rect 106922 0 106978 800
rect 112718 0 112774 800
rect 119158 0 119214 800
rect 125598 0 125654 800
rect 132038 0 132094 800
rect 138478 0 138534 800
rect 144274 0 144330 800
rect 150714 0 150770 800
rect 157154 0 157210 800
rect 163594 0 163650 800
rect 169390 0 169446 800
rect 175830 0 175886 800
rect 182270 0 182326 800
rect 188710 0 188766 800
rect 195150 0 195206 800
rect 200946 0 201002 800
rect 207386 0 207442 800
rect 213826 0 213882 800
rect 220266 0 220322 800
rect 226062 0 226118 800
rect 232502 0 232558 800
rect 238942 0 238998 800
rect 245382 0 245438 800
rect 251822 0 251878 800
rect 257618 0 257674 800
rect 264058 0 264114 800
rect 270498 0 270554 800
rect 276938 0 276994 800
rect 282734 0 282790 800
rect 289174 0 289230 800
rect 295614 0 295670 800
rect 302054 0 302110 800
rect 308494 0 308550 800
rect 314290 0 314346 800
rect 320730 0 320786 800
rect 327170 0 327226 800
rect 333610 0 333666 800
rect 339406 0 339462 800
rect 345846 0 345902 800
rect 352286 0 352342 800
rect 358726 0 358782 800
rect 365166 0 365222 800
rect 370962 0 371018 800
rect 377402 0 377458 800
rect 383842 0 383898 800
rect 390282 0 390338 800
rect 396078 0 396134 800
rect 402518 0 402574 800
rect 408958 0 409014 800
rect 415398 0 415454 800
rect 421838 0 421894 800
rect 427634 0 427690 800
rect 434074 0 434130 800
rect 440514 0 440570 800
rect 446954 0 447010 800
rect 452750 0 452806 800
rect 459190 0 459246 800
rect 465630 0 465686 800
rect 472070 0 472126 800
rect 478510 0 478566 800
rect 484306 0 484362 800
rect 490746 0 490802 800
rect 497186 0 497242 800
rect 503626 0 503682 800
rect 509422 0 509478 800
rect 515862 0 515918 800
rect 522302 0 522358 800
rect 528742 0 528798 800
rect 535182 0 535238 800
rect 540978 0 541034 800
rect 547418 0 547474 800
rect 553858 0 553914 800
rect 560298 0 560354 800
<< obsm2 >>
rect 130 683144 6402 683346
rect 6570 683144 12842 683346
rect 13010 683144 19282 683346
rect 19450 683144 25722 683346
rect 25890 683144 31518 683346
rect 31686 683144 37958 683346
rect 38126 683144 44398 683346
rect 44566 683144 50838 683346
rect 51006 683144 56634 683346
rect 56802 683144 63074 683346
rect 63242 683144 69514 683346
rect 69682 683144 75954 683346
rect 76122 683144 82394 683346
rect 82562 683144 88190 683346
rect 88358 683144 94630 683346
rect 94798 683144 101070 683346
rect 101238 683144 107510 683346
rect 107678 683144 113306 683346
rect 113474 683144 119746 683346
rect 119914 683144 126186 683346
rect 126354 683144 132626 683346
rect 132794 683144 139066 683346
rect 139234 683144 144862 683346
rect 145030 683144 151302 683346
rect 151470 683144 157742 683346
rect 157910 683144 164182 683346
rect 164350 683144 169978 683346
rect 170146 683144 176418 683346
rect 176586 683144 182858 683346
rect 183026 683144 189298 683346
rect 189466 683144 195738 683346
rect 195906 683144 201534 683346
rect 201702 683144 207974 683346
rect 208142 683144 214414 683346
rect 214582 683144 220854 683346
rect 221022 683144 226650 683346
rect 226818 683144 233090 683346
rect 233258 683144 239530 683346
rect 239698 683144 245970 683346
rect 246138 683144 252410 683346
rect 252578 683144 258206 683346
rect 258374 683144 264646 683346
rect 264814 683144 271086 683346
rect 271254 683144 277526 683346
rect 277694 683144 283322 683346
rect 283490 683144 289762 683346
rect 289930 683144 296202 683346
rect 296370 683144 302642 683346
rect 302810 683144 309082 683346
rect 309250 683144 314878 683346
rect 315046 683144 321318 683346
rect 321486 683144 327758 683346
rect 327926 683144 334198 683346
rect 334366 683144 339994 683346
rect 340162 683144 346434 683346
rect 346602 683144 352874 683346
rect 353042 683144 359314 683346
rect 359482 683144 365754 683346
rect 365922 683144 371550 683346
rect 371718 683144 377990 683346
rect 378158 683144 384430 683346
rect 384598 683144 390870 683346
rect 391038 683144 396666 683346
rect 396834 683144 403106 683346
rect 403274 683144 409546 683346
rect 409714 683144 415986 683346
rect 416154 683144 422426 683346
rect 422594 683144 428222 683346
rect 428390 683144 434662 683346
rect 434830 683144 441102 683346
rect 441270 683144 447542 683346
rect 447710 683144 453338 683346
rect 453506 683144 459778 683346
rect 459946 683144 466218 683346
rect 466386 683144 472658 683346
rect 472826 683144 479098 683346
rect 479266 683144 484894 683346
rect 485062 683144 491334 683346
rect 491502 683144 497774 683346
rect 497942 683144 504214 683346
rect 504382 683144 510010 683346
rect 510178 683144 516450 683346
rect 516618 683144 522890 683346
rect 523058 683144 529330 683346
rect 529498 683144 535770 683346
rect 535938 683144 541566 683346
rect 541734 683144 548006 683346
rect 548174 683144 554446 683346
rect 554614 683144 560886 683346
rect 561054 683144 562194 683346
rect 20 856 562194 683144
rect 130 800 5758 856
rect 5926 800 12198 856
rect 12366 800 18638 856
rect 18806 800 25078 856
rect 25246 800 30874 856
rect 31042 800 37314 856
rect 37482 800 43754 856
rect 43922 800 50194 856
rect 50362 800 55990 856
rect 56158 800 62430 856
rect 62598 800 68870 856
rect 69038 800 75310 856
rect 75478 800 81750 856
rect 81918 800 87546 856
rect 87714 800 93986 856
rect 94154 800 100426 856
rect 100594 800 106866 856
rect 107034 800 112662 856
rect 112830 800 119102 856
rect 119270 800 125542 856
rect 125710 800 131982 856
rect 132150 800 138422 856
rect 138590 800 144218 856
rect 144386 800 150658 856
rect 150826 800 157098 856
rect 157266 800 163538 856
rect 163706 800 169334 856
rect 169502 800 175774 856
rect 175942 800 182214 856
rect 182382 800 188654 856
rect 188822 800 195094 856
rect 195262 800 200890 856
rect 201058 800 207330 856
rect 207498 800 213770 856
rect 213938 800 220210 856
rect 220378 800 226006 856
rect 226174 800 232446 856
rect 232614 800 238886 856
rect 239054 800 245326 856
rect 245494 800 251766 856
rect 251934 800 257562 856
rect 257730 800 264002 856
rect 264170 800 270442 856
rect 270610 800 276882 856
rect 277050 800 282678 856
rect 282846 800 289118 856
rect 289286 800 295558 856
rect 295726 800 301998 856
rect 302166 800 308438 856
rect 308606 800 314234 856
rect 314402 800 320674 856
rect 320842 800 327114 856
rect 327282 800 333554 856
rect 333722 800 339350 856
rect 339518 800 345790 856
rect 345958 800 352230 856
rect 352398 800 358670 856
rect 358838 800 365110 856
rect 365278 800 370906 856
rect 371074 800 377346 856
rect 377514 800 383786 856
rect 383954 800 390226 856
rect 390394 800 396022 856
rect 396190 800 402462 856
rect 402630 800 408902 856
rect 409070 800 415342 856
rect 415510 800 421782 856
rect 421950 800 427578 856
rect 427746 800 434018 856
rect 434186 800 440458 856
rect 440626 800 446898 856
rect 447066 800 452694 856
rect 452862 800 459134 856
rect 459302 800 465574 856
rect 465742 800 472014 856
rect 472182 800 478454 856
rect 478622 800 484250 856
rect 484418 800 490690 856
rect 490858 800 497130 856
rect 497298 800 503570 856
rect 503738 800 509366 856
rect 509534 800 515806 856
rect 515974 800 522246 856
rect 522414 800 528686 856
rect 528854 800 535126 856
rect 535294 800 540922 856
rect 541090 800 547362 856
rect 547530 800 553802 856
rect 553970 800 560242 856
rect 560410 800 562194 856
<< metal3 >>
rect 563200 680688 564000 680808
rect 0 677968 800 678088
rect 563200 673888 564000 674008
rect 0 671168 800 671288
rect 563200 667088 564000 667208
rect 0 664368 800 664488
rect 563200 660288 564000 660408
rect 0 657568 800 657688
rect 563200 654168 564000 654288
rect 0 651448 800 651568
rect 563200 647368 564000 647488
rect 0 644648 800 644768
rect 563200 640568 564000 640688
rect 0 637848 800 637968
rect 563200 633768 564000 633888
rect 0 631048 800 631168
rect 563200 626968 564000 627088
rect 0 624928 800 625048
rect 563200 620848 564000 620968
rect 0 618128 800 618248
rect 563200 614048 564000 614168
rect 0 611328 800 611448
rect 563200 607248 564000 607368
rect 0 604528 800 604648
rect 563200 600448 564000 600568
rect 0 597728 800 597848
rect 563200 594328 564000 594448
rect 0 591608 800 591728
rect 563200 587528 564000 587648
rect 0 584808 800 584928
rect 563200 580728 564000 580848
rect 0 578008 800 578128
rect 563200 573928 564000 574048
rect 0 571208 800 571328
rect 563200 567128 564000 567248
rect 0 565088 800 565208
rect 563200 561008 564000 561128
rect 0 558288 800 558408
rect 563200 554208 564000 554328
rect 0 551488 800 551608
rect 563200 547408 564000 547528
rect 0 544688 800 544808
rect 563200 540608 564000 540728
rect 0 537888 800 538008
rect 563200 534488 564000 534608
rect 0 531768 800 531888
rect 563200 527688 564000 527808
rect 0 524968 800 525088
rect 563200 520888 564000 521008
rect 0 518168 800 518288
rect 563200 514088 564000 514208
rect 0 511368 800 511488
rect 563200 507288 564000 507408
rect 0 505248 800 505368
rect 563200 501168 564000 501288
rect 0 498448 800 498568
rect 563200 494368 564000 494488
rect 0 491648 800 491768
rect 563200 487568 564000 487688
rect 0 484848 800 484968
rect 563200 480768 564000 480888
rect 0 478048 800 478168
rect 563200 474648 564000 474768
rect 0 471928 800 472048
rect 563200 467848 564000 467968
rect 0 465128 800 465248
rect 563200 461048 564000 461168
rect 0 458328 800 458448
rect 563200 454248 564000 454368
rect 0 451528 800 451648
rect 563200 447448 564000 447568
rect 0 445408 800 445528
rect 563200 441328 564000 441448
rect 0 438608 800 438728
rect 563200 434528 564000 434648
rect 0 431808 800 431928
rect 563200 427728 564000 427848
rect 0 425008 800 425128
rect 563200 420928 564000 421048
rect 0 418208 800 418328
rect 563200 414808 564000 414928
rect 0 412088 800 412208
rect 563200 408008 564000 408128
rect 0 405288 800 405408
rect 563200 401208 564000 401328
rect 0 398488 800 398608
rect 563200 394408 564000 394528
rect 0 391688 800 391808
rect 563200 387608 564000 387728
rect 0 385568 800 385688
rect 563200 381488 564000 381608
rect 0 378768 800 378888
rect 563200 374688 564000 374808
rect 0 371968 800 372088
rect 563200 367888 564000 368008
rect 0 365168 800 365288
rect 563200 361088 564000 361208
rect 0 358368 800 358488
rect 563200 354968 564000 355088
rect 0 352248 800 352368
rect 563200 348168 564000 348288
rect 0 345448 800 345568
rect 563200 341368 564000 341488
rect 0 338648 800 338768
rect 563200 334568 564000 334688
rect 0 331848 800 331968
rect 563200 327768 564000 327888
rect 0 325728 800 325848
rect 563200 321648 564000 321768
rect 0 318928 800 319048
rect 563200 314848 564000 314968
rect 0 312128 800 312248
rect 563200 308048 564000 308168
rect 0 305328 800 305448
rect 563200 301248 564000 301368
rect 0 298528 800 298648
rect 563200 295128 564000 295248
rect 0 292408 800 292528
rect 563200 288328 564000 288448
rect 0 285608 800 285728
rect 563200 281528 564000 281648
rect 0 278808 800 278928
rect 563200 274728 564000 274848
rect 0 272008 800 272128
rect 563200 267928 564000 268048
rect 0 265888 800 266008
rect 563200 261808 564000 261928
rect 0 259088 800 259208
rect 563200 255008 564000 255128
rect 0 252288 800 252408
rect 563200 248208 564000 248328
rect 0 245488 800 245608
rect 563200 241408 564000 241528
rect 0 238688 800 238808
rect 563200 235288 564000 235408
rect 0 232568 800 232688
rect 563200 228488 564000 228608
rect 0 225768 800 225888
rect 563200 221688 564000 221808
rect 0 218968 800 219088
rect 563200 214888 564000 215008
rect 0 212168 800 212288
rect 563200 208088 564000 208208
rect 0 206048 800 206168
rect 563200 201968 564000 202088
rect 0 199248 800 199368
rect 563200 195168 564000 195288
rect 0 192448 800 192568
rect 563200 188368 564000 188488
rect 0 185648 800 185768
rect 563200 181568 564000 181688
rect 0 178848 800 178968
rect 563200 175448 564000 175568
rect 0 172728 800 172848
rect 563200 168648 564000 168768
rect 0 165928 800 166048
rect 563200 161848 564000 161968
rect 0 159128 800 159248
rect 563200 155048 564000 155168
rect 0 152328 800 152448
rect 563200 148248 564000 148368
rect 0 146208 800 146328
rect 563200 142128 564000 142248
rect 0 139408 800 139528
rect 563200 135328 564000 135448
rect 0 132608 800 132728
rect 563200 128528 564000 128648
rect 0 125808 800 125928
rect 563200 121728 564000 121848
rect 0 119008 800 119128
rect 563200 115608 564000 115728
rect 0 112888 800 113008
rect 563200 108808 564000 108928
rect 0 106088 800 106208
rect 563200 102008 564000 102128
rect 0 99288 800 99408
rect 563200 95208 564000 95328
rect 0 92488 800 92608
rect 563200 88408 564000 88528
rect 0 86368 800 86488
rect 563200 82288 564000 82408
rect 0 79568 800 79688
rect 563200 75488 564000 75608
rect 0 72768 800 72888
rect 563200 68688 564000 68808
rect 0 65968 800 66088
rect 563200 61888 564000 62008
rect 0 59168 800 59288
rect 563200 55768 564000 55888
rect 0 53048 800 53168
rect 563200 48968 564000 49088
rect 0 46248 800 46368
rect 563200 42168 564000 42288
rect 0 39448 800 39568
rect 563200 35368 564000 35488
rect 0 32648 800 32768
rect 563200 29248 564000 29368
rect 0 26528 800 26648
rect 563200 22448 564000 22568
rect 0 19728 800 19848
rect 563200 15648 564000 15768
rect 0 12928 800 13048
rect 563200 8848 564000 8968
rect 0 6128 800 6248
rect 563200 2048 564000 2168
<< obsm3 >>
rect 800 680888 563200 681665
rect 800 680608 563120 680888
rect 800 678168 563200 680608
rect 880 677888 563200 678168
rect 800 674088 563200 677888
rect 800 673808 563120 674088
rect 800 671368 563200 673808
rect 880 671088 563200 671368
rect 800 667288 563200 671088
rect 800 667008 563120 667288
rect 800 664568 563200 667008
rect 880 664288 563200 664568
rect 800 660488 563200 664288
rect 800 660208 563120 660488
rect 800 657768 563200 660208
rect 880 657488 563200 657768
rect 800 654368 563200 657488
rect 800 654088 563120 654368
rect 800 651648 563200 654088
rect 880 651368 563200 651648
rect 800 647568 563200 651368
rect 800 647288 563120 647568
rect 800 644848 563200 647288
rect 880 644568 563200 644848
rect 800 640768 563200 644568
rect 800 640488 563120 640768
rect 800 638048 563200 640488
rect 880 637768 563200 638048
rect 800 633968 563200 637768
rect 800 633688 563120 633968
rect 800 631248 563200 633688
rect 880 630968 563200 631248
rect 800 627168 563200 630968
rect 800 626888 563120 627168
rect 800 625128 563200 626888
rect 880 624848 563200 625128
rect 800 621048 563200 624848
rect 800 620768 563120 621048
rect 800 618328 563200 620768
rect 880 618048 563200 618328
rect 800 614248 563200 618048
rect 800 613968 563120 614248
rect 800 611528 563200 613968
rect 880 611248 563200 611528
rect 800 607448 563200 611248
rect 800 607168 563120 607448
rect 800 604728 563200 607168
rect 880 604448 563200 604728
rect 800 600648 563200 604448
rect 800 600368 563120 600648
rect 800 597928 563200 600368
rect 880 597648 563200 597928
rect 800 594528 563200 597648
rect 800 594248 563120 594528
rect 800 591808 563200 594248
rect 880 591528 563200 591808
rect 800 587728 563200 591528
rect 800 587448 563120 587728
rect 800 585008 563200 587448
rect 880 584728 563200 585008
rect 800 580928 563200 584728
rect 800 580648 563120 580928
rect 800 578208 563200 580648
rect 880 577928 563200 578208
rect 800 574128 563200 577928
rect 800 573848 563120 574128
rect 800 571408 563200 573848
rect 880 571128 563200 571408
rect 800 567328 563200 571128
rect 800 567048 563120 567328
rect 800 565288 563200 567048
rect 880 565008 563200 565288
rect 800 561208 563200 565008
rect 800 560928 563120 561208
rect 800 558488 563200 560928
rect 880 558208 563200 558488
rect 800 554408 563200 558208
rect 800 554128 563120 554408
rect 800 551688 563200 554128
rect 880 551408 563200 551688
rect 800 547608 563200 551408
rect 800 547328 563120 547608
rect 800 544888 563200 547328
rect 880 544608 563200 544888
rect 800 540808 563200 544608
rect 800 540528 563120 540808
rect 800 538088 563200 540528
rect 880 537808 563200 538088
rect 800 534688 563200 537808
rect 800 534408 563120 534688
rect 800 531968 563200 534408
rect 880 531688 563200 531968
rect 800 527888 563200 531688
rect 800 527608 563120 527888
rect 800 525168 563200 527608
rect 880 524888 563200 525168
rect 800 521088 563200 524888
rect 800 520808 563120 521088
rect 800 518368 563200 520808
rect 880 518088 563200 518368
rect 800 514288 563200 518088
rect 800 514008 563120 514288
rect 800 511568 563200 514008
rect 880 511288 563200 511568
rect 800 507488 563200 511288
rect 800 507208 563120 507488
rect 800 505448 563200 507208
rect 880 505168 563200 505448
rect 800 501368 563200 505168
rect 800 501088 563120 501368
rect 800 498648 563200 501088
rect 880 498368 563200 498648
rect 800 494568 563200 498368
rect 800 494288 563120 494568
rect 800 491848 563200 494288
rect 880 491568 563200 491848
rect 800 487768 563200 491568
rect 800 487488 563120 487768
rect 800 485048 563200 487488
rect 880 484768 563200 485048
rect 800 480968 563200 484768
rect 800 480688 563120 480968
rect 800 478248 563200 480688
rect 880 477968 563200 478248
rect 800 474848 563200 477968
rect 800 474568 563120 474848
rect 800 472128 563200 474568
rect 880 471848 563200 472128
rect 800 468048 563200 471848
rect 800 467768 563120 468048
rect 800 465328 563200 467768
rect 880 465048 563200 465328
rect 800 461248 563200 465048
rect 800 460968 563120 461248
rect 800 458528 563200 460968
rect 880 458248 563200 458528
rect 800 454448 563200 458248
rect 800 454168 563120 454448
rect 800 451728 563200 454168
rect 880 451448 563200 451728
rect 800 447648 563200 451448
rect 800 447368 563120 447648
rect 800 445608 563200 447368
rect 880 445328 563200 445608
rect 800 441528 563200 445328
rect 800 441248 563120 441528
rect 800 438808 563200 441248
rect 880 438528 563200 438808
rect 800 434728 563200 438528
rect 800 434448 563120 434728
rect 800 432008 563200 434448
rect 880 431728 563200 432008
rect 800 427928 563200 431728
rect 800 427648 563120 427928
rect 800 425208 563200 427648
rect 880 424928 563200 425208
rect 800 421128 563200 424928
rect 800 420848 563120 421128
rect 800 418408 563200 420848
rect 880 418128 563200 418408
rect 800 415008 563200 418128
rect 800 414728 563120 415008
rect 800 412288 563200 414728
rect 880 412008 563200 412288
rect 800 408208 563200 412008
rect 800 407928 563120 408208
rect 800 405488 563200 407928
rect 880 405208 563200 405488
rect 800 401408 563200 405208
rect 800 401128 563120 401408
rect 800 398688 563200 401128
rect 880 398408 563200 398688
rect 800 394608 563200 398408
rect 800 394328 563120 394608
rect 800 391888 563200 394328
rect 880 391608 563200 391888
rect 800 387808 563200 391608
rect 800 387528 563120 387808
rect 800 385768 563200 387528
rect 880 385488 563200 385768
rect 800 381688 563200 385488
rect 800 381408 563120 381688
rect 800 378968 563200 381408
rect 880 378688 563200 378968
rect 800 374888 563200 378688
rect 800 374608 563120 374888
rect 800 372168 563200 374608
rect 880 371888 563200 372168
rect 800 368088 563200 371888
rect 800 367808 563120 368088
rect 800 365368 563200 367808
rect 880 365088 563200 365368
rect 800 361288 563200 365088
rect 800 361008 563120 361288
rect 800 358568 563200 361008
rect 880 358288 563200 358568
rect 800 355168 563200 358288
rect 800 354888 563120 355168
rect 800 352448 563200 354888
rect 880 352168 563200 352448
rect 800 348368 563200 352168
rect 800 348088 563120 348368
rect 800 345648 563200 348088
rect 880 345368 563200 345648
rect 800 341568 563200 345368
rect 800 341288 563120 341568
rect 800 338848 563200 341288
rect 880 338568 563200 338848
rect 800 334768 563200 338568
rect 800 334488 563120 334768
rect 800 332048 563200 334488
rect 880 331768 563200 332048
rect 800 327968 563200 331768
rect 800 327688 563120 327968
rect 800 325928 563200 327688
rect 880 325648 563200 325928
rect 800 321848 563200 325648
rect 800 321568 563120 321848
rect 800 319128 563200 321568
rect 880 318848 563200 319128
rect 800 315048 563200 318848
rect 800 314768 563120 315048
rect 800 312328 563200 314768
rect 880 312048 563200 312328
rect 800 308248 563200 312048
rect 800 307968 563120 308248
rect 800 305528 563200 307968
rect 880 305248 563200 305528
rect 800 301448 563200 305248
rect 800 301168 563120 301448
rect 800 298728 563200 301168
rect 880 298448 563200 298728
rect 800 295328 563200 298448
rect 800 295048 563120 295328
rect 800 292608 563200 295048
rect 880 292328 563200 292608
rect 800 288528 563200 292328
rect 800 288248 563120 288528
rect 800 285808 563200 288248
rect 880 285528 563200 285808
rect 800 281728 563200 285528
rect 800 281448 563120 281728
rect 800 279008 563200 281448
rect 880 278728 563200 279008
rect 800 274928 563200 278728
rect 800 274648 563120 274928
rect 800 272208 563200 274648
rect 880 271928 563200 272208
rect 800 268128 563200 271928
rect 800 267848 563120 268128
rect 800 266088 563200 267848
rect 880 265808 563200 266088
rect 800 262008 563200 265808
rect 800 261728 563120 262008
rect 800 259288 563200 261728
rect 880 259008 563200 259288
rect 800 255208 563200 259008
rect 800 254928 563120 255208
rect 800 252488 563200 254928
rect 880 252208 563200 252488
rect 800 248408 563200 252208
rect 800 248128 563120 248408
rect 800 245688 563200 248128
rect 880 245408 563200 245688
rect 800 241608 563200 245408
rect 800 241328 563120 241608
rect 800 238888 563200 241328
rect 880 238608 563200 238888
rect 800 235488 563200 238608
rect 800 235208 563120 235488
rect 800 232768 563200 235208
rect 880 232488 563200 232768
rect 800 228688 563200 232488
rect 800 228408 563120 228688
rect 800 225968 563200 228408
rect 880 225688 563200 225968
rect 800 221888 563200 225688
rect 800 221608 563120 221888
rect 800 219168 563200 221608
rect 880 218888 563200 219168
rect 800 215088 563200 218888
rect 800 214808 563120 215088
rect 800 212368 563200 214808
rect 880 212088 563200 212368
rect 800 208288 563200 212088
rect 800 208008 563120 208288
rect 800 206248 563200 208008
rect 880 205968 563200 206248
rect 800 202168 563200 205968
rect 800 201888 563120 202168
rect 800 199448 563200 201888
rect 880 199168 563200 199448
rect 800 195368 563200 199168
rect 800 195088 563120 195368
rect 800 192648 563200 195088
rect 880 192368 563200 192648
rect 800 188568 563200 192368
rect 800 188288 563120 188568
rect 800 185848 563200 188288
rect 880 185568 563200 185848
rect 800 181768 563200 185568
rect 800 181488 563120 181768
rect 800 179048 563200 181488
rect 880 178768 563200 179048
rect 800 175648 563200 178768
rect 800 175368 563120 175648
rect 800 172928 563200 175368
rect 880 172648 563200 172928
rect 800 168848 563200 172648
rect 800 168568 563120 168848
rect 800 166128 563200 168568
rect 880 165848 563200 166128
rect 800 162048 563200 165848
rect 800 161768 563120 162048
rect 800 159328 563200 161768
rect 880 159048 563200 159328
rect 800 155248 563200 159048
rect 800 154968 563120 155248
rect 800 152528 563200 154968
rect 880 152248 563200 152528
rect 800 148448 563200 152248
rect 800 148168 563120 148448
rect 800 146408 563200 148168
rect 880 146128 563200 146408
rect 800 142328 563200 146128
rect 800 142048 563120 142328
rect 800 139608 563200 142048
rect 880 139328 563200 139608
rect 800 135528 563200 139328
rect 800 135248 563120 135528
rect 800 132808 563200 135248
rect 880 132528 563200 132808
rect 800 128728 563200 132528
rect 800 128448 563120 128728
rect 800 126008 563200 128448
rect 880 125728 563200 126008
rect 800 121928 563200 125728
rect 800 121648 563120 121928
rect 800 119208 563200 121648
rect 880 118928 563200 119208
rect 800 115808 563200 118928
rect 800 115528 563120 115808
rect 800 113088 563200 115528
rect 880 112808 563200 113088
rect 800 109008 563200 112808
rect 800 108728 563120 109008
rect 800 106288 563200 108728
rect 880 106008 563200 106288
rect 800 102208 563200 106008
rect 800 101928 563120 102208
rect 800 99488 563200 101928
rect 880 99208 563200 99488
rect 800 95408 563200 99208
rect 800 95128 563120 95408
rect 800 92688 563200 95128
rect 880 92408 563200 92688
rect 800 88608 563200 92408
rect 800 88328 563120 88608
rect 800 86568 563200 88328
rect 880 86288 563200 86568
rect 800 82488 563200 86288
rect 800 82208 563120 82488
rect 800 79768 563200 82208
rect 880 79488 563200 79768
rect 800 75688 563200 79488
rect 800 75408 563120 75688
rect 800 72968 563200 75408
rect 880 72688 563200 72968
rect 800 68888 563200 72688
rect 800 68608 563120 68888
rect 800 66168 563200 68608
rect 880 65888 563200 66168
rect 800 62088 563200 65888
rect 800 61808 563120 62088
rect 800 59368 563200 61808
rect 880 59088 563200 59368
rect 800 55968 563200 59088
rect 800 55688 563120 55968
rect 800 53248 563200 55688
rect 880 52968 563200 53248
rect 800 49168 563200 52968
rect 800 48888 563120 49168
rect 800 46448 563200 48888
rect 880 46168 563200 46448
rect 800 42368 563200 46168
rect 800 42088 563120 42368
rect 800 39648 563200 42088
rect 880 39368 563200 39648
rect 800 35568 563200 39368
rect 800 35288 563120 35568
rect 800 32848 563200 35288
rect 880 32568 563200 32848
rect 800 29448 563200 32568
rect 800 29168 563120 29448
rect 800 26728 563200 29168
rect 880 26448 563200 26728
rect 800 22648 563200 26448
rect 800 22368 563120 22648
rect 800 19928 563200 22368
rect 880 19648 563200 19928
rect 800 15848 563200 19648
rect 800 15568 563120 15848
rect 800 13128 563200 15568
rect 880 12848 563200 13128
rect 800 9048 563200 12848
rect 800 8768 563120 9048
rect 800 6328 563200 8768
rect 880 6048 563200 6328
rect 800 2248 563200 6048
rect 800 2075 563120 2248
<< metal4 >>
rect 4208 2128 4528 681680
rect 19568 2128 19888 681680
rect 34928 2128 35248 681680
rect 50288 2128 50608 681680
rect 65648 2128 65968 681680
rect 81008 2128 81328 681680
rect 96368 2128 96688 681680
rect 111728 2128 112048 681680
rect 127088 2128 127408 681680
rect 142448 2128 142768 681680
rect 157808 2128 158128 681680
rect 173168 2128 173488 681680
rect 188528 2128 188848 681680
rect 203888 2128 204208 681680
rect 219248 2128 219568 681680
rect 234608 2128 234928 681680
rect 249968 2128 250288 681680
rect 265328 2128 265648 681680
rect 280688 2128 281008 681680
rect 296048 2128 296368 681680
rect 311408 2128 311728 681680
rect 326768 2128 327088 681680
rect 342128 2128 342448 681680
rect 357488 2128 357808 681680
rect 372848 2128 373168 681680
rect 388208 2128 388528 681680
rect 403568 2128 403888 681680
rect 418928 2128 419248 681680
rect 434288 2128 434608 681680
rect 449648 2128 449968 681680
rect 465008 2128 465328 681680
rect 480368 2128 480688 681680
rect 495728 2128 496048 681680
rect 511088 2128 511408 681680
rect 526448 2128 526768 681680
rect 541808 2128 542128 681680
rect 557168 2128 557488 681680
<< obsm4 >>
rect 174491 2347 188448 681325
rect 188928 2347 203808 681325
rect 204288 2347 219168 681325
rect 219648 2347 234528 681325
rect 235008 2347 249888 681325
rect 250368 2347 265248 681325
rect 265728 2347 280608 681325
rect 281088 2347 295968 681325
rect 296448 2347 311328 681325
rect 311808 2347 326688 681325
rect 327168 2347 342048 681325
rect 342528 2347 357408 681325
rect 357888 2347 372768 681325
rect 373248 2347 378429 681325
<< labels >>
rlabel metal3 s 0 265888 800 266008 6 clk
port 1 nsew signal input
rlabel metal2 s 522946 683200 523002 684000 6 la_data_in[0]
port 2 nsew signal input
rlabel metal3 s 0 152328 800 152448 6 la_data_in[100]
port 3 nsew signal input
rlabel metal2 s 453394 683200 453450 684000 6 la_data_in[101]
port 4 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 la_data_in[102]
port 5 nsew signal input
rlabel metal3 s 0 385568 800 385688 6 la_data_in[103]
port 6 nsew signal input
rlabel metal3 s 0 352248 800 352368 6 la_data_in[104]
port 7 nsew signal input
rlabel metal3 s 563200 161848 564000 161968 6 la_data_in[105]
port 8 nsew signal input
rlabel metal3 s 0 558288 800 558408 6 la_data_in[106]
port 9 nsew signal input
rlabel metal2 s 201590 683200 201646 684000 6 la_data_in[107]
port 10 nsew signal input
rlabel metal2 s 164238 683200 164294 684000 6 la_data_in[108]
port 11 nsew signal input
rlabel metal2 s 371606 683200 371662 684000 6 la_data_in[109]
port 12 nsew signal input
rlabel metal3 s 563200 188368 564000 188488 6 la_data_in[10]
port 13 nsew signal input
rlabel metal2 s 497830 683200 497886 684000 6 la_data_in[110]
port 14 nsew signal input
rlabel metal3 s 0 412088 800 412208 6 la_data_in[111]
port 15 nsew signal input
rlabel metal2 s 320730 0 320786 800 6 la_data_in[112]
port 16 nsew signal input
rlabel metal3 s 563200 248208 564000 248328 6 la_data_in[113]
port 17 nsew signal input
rlabel metal2 s 541622 683200 541678 684000 6 la_data_in[114]
port 18 nsew signal input
rlabel metal3 s 0 511368 800 511488 6 la_data_in[115]
port 19 nsew signal input
rlabel metal3 s 0 165928 800 166048 6 la_data_in[116]
port 20 nsew signal input
rlabel metal3 s 563200 647368 564000 647488 6 la_data_in[117]
port 21 nsew signal input
rlabel metal3 s 563200 427728 564000 427848 6 la_data_in[118]
port 22 nsew signal input
rlabel metal2 s 547418 0 547474 800 6 la_data_in[119]
port 23 nsew signal input
rlabel metal2 s 428278 683200 428334 684000 6 la_data_in[11]
port 24 nsew signal input
rlabel metal2 s 383842 0 383898 800 6 la_data_in[120]
port 25 nsew signal input
rlabel metal3 s 0 624928 800 625048 6 la_data_in[121]
port 26 nsew signal input
rlabel metal2 s 189354 683200 189410 684000 6 la_data_in[122]
port 27 nsew signal input
rlabel metal3 s 563200 587528 564000 587648 6 la_data_in[123]
port 28 nsew signal input
rlabel metal3 s 563200 274728 564000 274848 6 la_data_in[124]
port 29 nsew signal input
rlabel metal3 s 0 611328 800 611448 6 la_data_in[125]
port 30 nsew signal input
rlabel metal2 s 409602 683200 409658 684000 6 la_data_in[126]
port 31 nsew signal input
rlabel metal3 s 563200 507288 564000 507408 6 la_data_in[127]
port 32 nsew signal input
rlabel metal2 s 138478 0 138534 800 6 la_data_in[12]
port 33 nsew signal input
rlabel metal3 s 563200 381488 564000 381608 6 la_data_in[13]
port 34 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 la_data_in[14]
port 35 nsew signal input
rlabel metal3 s 563200 29248 564000 29368 6 la_data_in[15]
port 36 nsew signal input
rlabel metal2 s 370962 0 371018 800 6 la_data_in[16]
port 37 nsew signal input
rlabel metal3 s 0 199248 800 199368 6 la_data_in[17]
port 38 nsew signal input
rlabel metal3 s 0 206048 800 206168 6 la_data_in[18]
port 39 nsew signal input
rlabel metal3 s 563200 195168 564000 195288 6 la_data_in[19]
port 40 nsew signal input
rlabel metal3 s 563200 640568 564000 640688 6 la_data_in[1]
port 41 nsew signal input
rlabel metal2 s 535182 0 535238 800 6 la_data_in[20]
port 42 nsew signal input
rlabel metal3 s 563200 474648 564000 474768 6 la_data_in[21]
port 43 nsew signal input
rlabel metal3 s 563200 680688 564000 680808 6 la_data_in[22]
port 44 nsew signal input
rlabel metal2 s 396078 0 396134 800 6 la_data_in[23]
port 45 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 la_data_in[24]
port 46 nsew signal input
rlabel metal2 s 107566 683200 107622 684000 6 la_data_in[25]
port 47 nsew signal input
rlabel metal2 s 94686 683200 94742 684000 6 la_data_in[26]
port 48 nsew signal input
rlabel metal2 s 264702 683200 264758 684000 6 la_data_in[27]
port 49 nsew signal input
rlabel metal3 s 0 478048 800 478168 6 la_data_in[28]
port 50 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_data_in[29]
port 51 nsew signal input
rlabel metal3 s 563200 554208 564000 554328 6 la_data_in[2]
port 52 nsew signal input
rlabel metal3 s 563200 354968 564000 355088 6 la_data_in[30]
port 53 nsew signal input
rlabel metal3 s 0 664368 800 664488 6 la_data_in[31]
port 54 nsew signal input
rlabel metal3 s 563200 2048 564000 2168 6 la_data_in[32]
port 55 nsew signal input
rlabel metal3 s 563200 128528 564000 128648 6 la_data_in[33]
port 56 nsew signal input
rlabel metal3 s 563200 441328 564000 441448 6 la_data_in[34]
port 57 nsew signal input
rlabel metal3 s 0 99288 800 99408 6 la_data_in[35]
port 58 nsew signal input
rlabel metal3 s 563200 673888 564000 674008 6 la_data_in[36]
port 59 nsew signal input
rlabel metal3 s 563200 327768 564000 327888 6 la_data_in[37]
port 60 nsew signal input
rlabel metal3 s 563200 614048 564000 614168 6 la_data_in[38]
port 61 nsew signal input
rlabel metal3 s 0 465128 800 465248 6 la_data_in[39]
port 62 nsew signal input
rlabel metal2 s 346490 683200 346546 684000 6 la_data_in[3]
port 63 nsew signal input
rlabel metal3 s 0 498448 800 498568 6 la_data_in[40]
port 64 nsew signal input
rlabel metal2 s 144274 0 144330 800 6 la_data_in[41]
port 65 nsew signal input
rlabel metal2 s 522302 0 522358 800 6 la_data_in[42]
port 66 nsew signal input
rlabel metal2 s 252466 683200 252522 684000 6 la_data_in[43]
port 67 nsew signal input
rlabel metal2 s 427634 0 427690 800 6 la_data_in[44]
port 68 nsew signal input
rlabel metal2 s 441158 683200 441214 684000 6 la_data_in[45]
port 69 nsew signal input
rlabel metal3 s 563200 22448 564000 22568 6 la_data_in[46]
port 70 nsew signal input
rlabel metal2 s 339406 0 339462 800 6 la_data_in[47]
port 71 nsew signal input
rlabel metal2 s 309138 683200 309194 684000 6 la_data_in[48]
port 72 nsew signal input
rlabel metal2 s 308494 0 308550 800 6 la_data_in[49]
port 73 nsew signal input
rlabel metal3 s 563200 561008 564000 561128 6 la_data_in[4]
port 74 nsew signal input
rlabel metal2 s 214470 683200 214526 684000 6 la_data_in[50]
port 75 nsew signal input
rlabel metal3 s 563200 374688 564000 374808 6 la_data_in[51]
port 76 nsew signal input
rlabel metal2 s 472070 0 472126 800 6 la_data_in[52]
port 77 nsew signal input
rlabel metal3 s 563200 527688 564000 527808 6 la_data_in[53]
port 78 nsew signal input
rlabel metal3 s 563200 520888 564000 521008 6 la_data_in[54]
port 79 nsew signal input
rlabel metal2 s 264058 0 264114 800 6 la_data_in[55]
port 80 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 la_data_in[56]
port 81 nsew signal input
rlabel metal3 s 0 418208 800 418328 6 la_data_in[57]
port 82 nsew signal input
rlabel metal3 s 563200 168648 564000 168768 6 la_data_in[58]
port 83 nsew signal input
rlabel metal2 s 76010 683200 76066 684000 6 la_data_in[59]
port 84 nsew signal input
rlabel metal2 s 484306 0 484362 800 6 la_data_in[5]
port 85 nsew signal input
rlabel metal3 s 563200 55768 564000 55888 6 la_data_in[60]
port 86 nsew signal input
rlabel metal3 s 0 651448 800 651568 6 la_data_in[61]
port 87 nsew signal input
rlabel metal3 s 0 238688 800 238808 6 la_data_in[62]
port 88 nsew signal input
rlabel metal3 s 563200 654168 564000 654288 6 la_data_in[63]
port 89 nsew signal input
rlabel metal2 s 226062 0 226118 800 6 la_data_in[64]
port 90 nsew signal input
rlabel metal2 s 282734 0 282790 800 6 la_data_in[65]
port 91 nsew signal input
rlabel metal2 s 56690 683200 56746 684000 6 la_data_in[66]
port 92 nsew signal input
rlabel metal3 s 563200 600448 564000 600568 6 la_data_in[67]
port 93 nsew signal input
rlabel metal2 s 113362 683200 113418 684000 6 la_data_in[68]
port 94 nsew signal input
rlabel metal3 s 0 677968 800 678088 6 la_data_in[69]
port 95 nsew signal input
rlabel metal3 s 0 484848 800 484968 6 la_data_in[6]
port 96 nsew signal input
rlabel metal2 s 44454 683200 44510 684000 6 la_data_in[70]
port 97 nsew signal input
rlabel metal3 s 563200 201968 564000 202088 6 la_data_in[71]
port 98 nsew signal input
rlabel metal2 s 182270 0 182326 800 6 la_data_in[72]
port 99 nsew signal input
rlabel metal2 s 233146 683200 233202 684000 6 la_data_in[73]
port 100 nsew signal input
rlabel metal3 s 0 159128 800 159248 6 la_data_in[74]
port 101 nsew signal input
rlabel metal2 s 258262 683200 258318 684000 6 la_data_in[75]
port 102 nsew signal input
rlabel metal3 s 563200 108808 564000 108928 6 la_data_in[76]
port 103 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 la_data_in[77]
port 104 nsew signal input
rlabel metal2 s 314934 683200 314990 684000 6 la_data_in[78]
port 105 nsew signal input
rlabel metal3 s 563200 480768 564000 480888 6 la_data_in[79]
port 106 nsew signal input
rlabel metal3 s 563200 88408 564000 88528 6 la_data_in[7]
port 107 nsew signal input
rlabel metal2 s 560942 683200 560998 684000 6 la_data_in[80]
port 108 nsew signal input
rlabel metal3 s 0 365168 800 365288 6 la_data_in[81]
port 109 nsew signal input
rlabel metal2 s 321374 683200 321430 684000 6 la_data_in[82]
port 110 nsew signal input
rlabel metal2 s 484950 683200 485006 684000 6 la_data_in[83]
port 111 nsew signal input
rlabel metal3 s 563200 573928 564000 574048 6 la_data_in[84]
port 112 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 la_data_in[85]
port 113 nsew signal input
rlabel metal3 s 563200 567128 564000 567248 6 la_data_in[86]
port 114 nsew signal input
rlabel metal3 s 0 278808 800 278928 6 la_data_in[87]
port 115 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 la_data_in[88]
port 116 nsew signal input
rlabel metal2 s 19338 683200 19394 684000 6 la_data_in[89]
port 117 nsew signal input
rlabel metal3 s 0 445408 800 445528 6 la_data_in[8]
port 118 nsew signal input
rlabel metal2 s 251822 0 251878 800 6 la_data_in[90]
port 119 nsew signal input
rlabel metal2 s 200946 0 201002 800 6 la_data_in[91]
port 120 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 la_data_in[92]
port 121 nsew signal input
rlabel metal2 s 528742 0 528798 800 6 la_data_in[93]
port 122 nsew signal input
rlabel metal2 s 169390 0 169446 800 6 la_data_in[94]
port 123 nsew signal input
rlabel metal3 s 0 637848 800 637968 6 la_data_in[95]
port 124 nsew signal input
rlabel metal3 s 0 451528 800 451648 6 la_data_in[96]
port 125 nsew signal input
rlabel metal2 s 139122 683200 139178 684000 6 la_data_in[97]
port 126 nsew signal input
rlabel metal3 s 0 192448 800 192568 6 la_data_in[98]
port 127 nsew signal input
rlabel metal2 s 239586 683200 239642 684000 6 la_data_in[99]
port 128 nsew signal input
rlabel metal3 s 563200 288328 564000 288448 6 la_data_in[9]
port 129 nsew signal input
rlabel metal2 s 245382 0 245438 800 6 la_data_out[0]
port 130 nsew signal output
rlabel metal3 s 563200 148248 564000 148368 6 la_data_out[100]
port 131 nsew signal output
rlabel metal3 s 0 644648 800 644768 6 la_data_out[101]
port 132 nsew signal output
rlabel metal3 s 563200 121728 564000 121848 6 la_data_out[102]
port 133 nsew signal output
rlabel metal3 s 0 185648 800 185768 6 la_data_out[103]
port 134 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 la_data_out[104]
port 135 nsew signal output
rlabel metal2 s 553858 0 553914 800 6 la_data_out[105]
port 136 nsew signal output
rlabel metal2 s 195150 0 195206 800 6 la_data_out[106]
port 137 nsew signal output
rlabel metal2 s 466274 683200 466330 684000 6 la_data_out[107]
port 138 nsew signal output
rlabel metal3 s 0 391688 800 391808 6 la_data_out[108]
port 139 nsew signal output
rlabel metal2 s 6458 683200 6514 684000 6 la_data_out[109]
port 140 nsew signal output
rlabel metal2 s 276938 0 276994 800 6 la_data_out[10]
port 141 nsew signal output
rlabel metal3 s 0 604528 800 604648 6 la_data_out[110]
port 142 nsew signal output
rlabel metal2 s 296258 683200 296314 684000 6 la_data_out[111]
port 143 nsew signal output
rlabel metal2 s 327814 683200 327870 684000 6 la_data_out[112]
port 144 nsew signal output
rlabel metal3 s 563200 181568 564000 181688 6 la_data_out[113]
port 145 nsew signal output
rlabel metal3 s 563200 620848 564000 620968 6 la_data_out[114]
port 146 nsew signal output
rlabel metal2 s 497186 0 497242 800 6 la_data_out[115]
port 147 nsew signal output
rlabel metal3 s 563200 267928 564000 268048 6 la_data_out[116]
port 148 nsew signal output
rlabel metal3 s 563200 281528 564000 281648 6 la_data_out[117]
port 149 nsew signal output
rlabel metal2 s 390282 0 390338 800 6 la_data_out[118]
port 150 nsew signal output
rlabel metal2 s 175830 0 175886 800 6 la_data_out[119]
port 151 nsew signal output
rlabel metal2 s 207386 0 207442 800 6 la_data_out[11]
port 152 nsew signal output
rlabel metal3 s 563200 214888 564000 215008 6 la_data_out[120]
port 153 nsew signal output
rlabel metal3 s 563200 547408 564000 547528 6 la_data_out[121]
port 154 nsew signal output
rlabel metal3 s 0 458328 800 458448 6 la_data_out[122]
port 155 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 la_data_out[123]
port 156 nsew signal output
rlabel metal3 s 563200 461048 564000 461168 6 la_data_out[124]
port 157 nsew signal output
rlabel metal3 s 0 398488 800 398608 6 la_data_out[125]
port 158 nsew signal output
rlabel metal3 s 563200 255008 564000 255128 6 la_data_out[126]
port 159 nsew signal output
rlabel metal3 s 0 671168 800 671288 6 la_data_out[127]
port 160 nsew signal output
rlabel metal3 s 563200 394408 564000 394528 6 la_data_out[12]
port 161 nsew signal output
rlabel metal2 s 334254 683200 334310 684000 6 la_data_out[13]
port 162 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 la_data_out[14]
port 163 nsew signal output
rlabel metal3 s 563200 155048 564000 155168 6 la_data_out[15]
port 164 nsew signal output
rlabel metal2 s 283378 683200 283434 684000 6 la_data_out[16]
port 165 nsew signal output
rlabel metal3 s 0 112888 800 113008 6 la_data_out[17]
port 166 nsew signal output
rlabel metal2 s 88246 683200 88302 684000 6 la_data_out[18]
port 167 nsew signal output
rlabel metal3 s 563200 454248 564000 454368 6 la_data_out[19]
port 168 nsew signal output
rlabel metal2 s 238942 0 238998 800 6 la_data_out[1]
port 169 nsew signal output
rlabel metal2 s 213826 0 213882 800 6 la_data_out[20]
port 170 nsew signal output
rlabel metal3 s 563200 261808 564000 261928 6 la_data_out[21]
port 171 nsew signal output
rlabel metal2 s 151358 683200 151414 684000 6 la_data_out[22]
port 172 nsew signal output
rlabel metal2 s 50894 683200 50950 684000 6 la_data_out[23]
port 173 nsew signal output
rlabel metal3 s 563200 102008 564000 102128 6 la_data_out[24]
port 174 nsew signal output
rlabel metal2 s 270498 0 270554 800 6 la_data_out[25]
port 175 nsew signal output
rlabel metal2 s 491390 683200 491446 684000 6 la_data_out[26]
port 176 nsew signal output
rlabel metal3 s 563200 467848 564000 467968 6 la_data_out[27]
port 177 nsew signal output
rlabel metal3 s 0 106088 800 106208 6 la_data_out[28]
port 178 nsew signal output
rlabel metal3 s 0 618128 800 618248 6 la_data_out[29]
port 179 nsew signal output
rlabel metal3 s 0 259088 800 259208 6 la_data_out[2]
port 180 nsew signal output
rlabel metal2 s 352286 0 352342 800 6 la_data_out[30]
port 181 nsew signal output
rlabel metal2 s 101126 683200 101182 684000 6 la_data_out[31]
port 182 nsew signal output
rlabel metal2 s 472714 683200 472770 684000 6 la_data_out[32]
port 183 nsew signal output
rlabel metal3 s 563200 494368 564000 494488 6 la_data_out[33]
port 184 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 la_data_out[34]
port 185 nsew signal output
rlabel metal3 s 0 537888 800 538008 6 la_data_out[35]
port 186 nsew signal output
rlabel metal2 s 18 683200 74 684000 6 la_data_out[36]
port 187 nsew signal output
rlabel metal2 s 340050 683200 340106 684000 6 la_data_out[37]
port 188 nsew signal output
rlabel metal3 s 0 491648 800 491768 6 la_data_out[38]
port 189 nsew signal output
rlabel metal3 s 0 86368 800 86488 6 la_data_out[39]
port 190 nsew signal output
rlabel metal2 s 509422 0 509478 800 6 la_data_out[3]
port 191 nsew signal output
rlabel metal3 s 563200 308048 564000 308168 6 la_data_out[40]
port 192 nsew signal output
rlabel metal3 s 563200 68688 564000 68808 6 la_data_out[41]
port 193 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 la_data_out[42]
port 194 nsew signal output
rlabel metal2 s 226706 683200 226762 684000 6 la_data_out[43]
port 195 nsew signal output
rlabel metal2 s 314290 0 314346 800 6 la_data_out[44]
port 196 nsew signal output
rlabel metal3 s 0 631048 800 631168 6 la_data_out[45]
port 197 nsew signal output
rlabel metal2 s 289174 0 289230 800 6 la_data_out[46]
port 198 nsew signal output
rlabel metal3 s 563200 142128 564000 142248 6 la_data_out[47]
port 199 nsew signal output
rlabel metal2 s 504270 683200 504326 684000 6 la_data_out[48]
port 200 nsew signal output
rlabel metal3 s 0 125808 800 125928 6 la_data_out[49]
port 201 nsew signal output
rlabel metal2 s 302698 683200 302754 684000 6 la_data_out[4]
port 202 nsew signal output
rlabel metal3 s 0 225768 800 225888 6 la_data_out[50]
port 203 nsew signal output
rlabel metal2 s 529386 683200 529442 684000 6 la_data_out[51]
port 204 nsew signal output
rlabel metal2 s 63130 683200 63186 684000 6 la_data_out[52]
port 205 nsew signal output
rlabel metal3 s 0 172728 800 172848 6 la_data_out[53]
port 206 nsew signal output
rlabel metal3 s 563200 48968 564000 49088 6 la_data_out[54]
port 207 nsew signal output
rlabel metal3 s 0 584808 800 584928 6 la_data_out[55]
port 208 nsew signal output
rlabel metal3 s 0 544688 800 544808 6 la_data_out[56]
port 209 nsew signal output
rlabel metal2 s 358726 0 358782 800 6 la_data_out[57]
port 210 nsew signal output
rlabel metal3 s 563200 295128 564000 295248 6 la_data_out[58]
port 211 nsew signal output
rlabel metal3 s 563200 235288 564000 235408 6 la_data_out[59]
port 212 nsew signal output
rlabel metal2 s 170034 683200 170090 684000 6 la_data_out[5]
port 213 nsew signal output
rlabel metal3 s 563200 348168 564000 348288 6 la_data_out[60]
port 214 nsew signal output
rlabel metal2 s 434074 0 434130 800 6 la_data_out[61]
port 215 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 la_data_out[62]
port 216 nsew signal output
rlabel metal2 s 421838 0 421894 800 6 la_data_out[63]
port 217 nsew signal output
rlabel metal2 s 503626 0 503682 800 6 la_data_out[64]
port 218 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 la_data_out[65]
port 219 nsew signal output
rlabel metal3 s 0 431808 800 431928 6 la_data_out[66]
port 220 nsew signal output
rlabel metal2 s 459190 0 459246 800 6 la_data_out[67]
port 221 nsew signal output
rlabel metal3 s 0 298528 800 298648 6 la_data_out[68]
port 222 nsew signal output
rlabel metal3 s 0 471928 800 472048 6 la_data_out[69]
port 223 nsew signal output
rlabel metal3 s 563200 667088 564000 667208 6 la_data_out[6]
port 224 nsew signal output
rlabel metal3 s 0 132608 800 132728 6 la_data_out[70]
port 225 nsew signal output
rlabel metal3 s 0 345448 800 345568 6 la_data_out[71]
port 226 nsew signal output
rlabel metal2 s 163594 0 163650 800 6 la_data_out[72]
port 227 nsew signal output
rlabel metal3 s 563200 387608 564000 387728 6 la_data_out[73]
port 228 nsew signal output
rlabel metal2 s 515862 0 515918 800 6 la_data_out[74]
port 229 nsew signal output
rlabel metal2 s 434718 683200 434774 684000 6 la_data_out[75]
port 230 nsew signal output
rlabel metal2 s 106922 0 106978 800 6 la_data_out[76]
port 231 nsew signal output
rlabel metal2 s 82450 683200 82506 684000 6 la_data_out[77]
port 232 nsew signal output
rlabel metal3 s 563200 594328 564000 594448 6 la_data_out[78]
port 233 nsew signal output
rlabel metal3 s 0 232568 800 232688 6 la_data_out[79]
port 234 nsew signal output
rlabel metal3 s 563200 540608 564000 540728 6 la_data_out[7]
port 235 nsew signal output
rlabel metal2 s 289818 683200 289874 684000 6 la_data_out[80]
port 236 nsew signal output
rlabel metal3 s 0 65968 800 66088 6 la_data_out[81]
port 237 nsew signal output
rlabel metal3 s 0 285608 800 285728 6 la_data_out[82]
port 238 nsew signal output
rlabel metal3 s 0 378768 800 378888 6 la_data_out[83]
port 239 nsew signal output
rlabel metal2 s 220910 683200 220966 684000 6 la_data_out[84]
port 240 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 la_data_out[85]
port 241 nsew signal output
rlabel metal2 s 126242 683200 126298 684000 6 la_data_out[86]
port 242 nsew signal output
rlabel metal2 s 302054 0 302110 800 6 la_data_out[87]
port 243 nsew signal output
rlabel metal3 s 563200 42168 564000 42288 6 la_data_out[88]
port 244 nsew signal output
rlabel metal3 s 563200 660288 564000 660408 6 la_data_out[89]
port 245 nsew signal output
rlabel metal3 s 563200 95208 564000 95328 6 la_data_out[8]
port 246 nsew signal output
rlabel metal2 s 246026 683200 246082 684000 6 la_data_out[90]
port 247 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 la_data_out[91]
port 248 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 la_data_out[92]
port 249 nsew signal output
rlabel metal2 s 257618 0 257674 800 6 la_data_out[93]
port 250 nsew signal output
rlabel metal2 s 510066 683200 510122 684000 6 la_data_out[94]
port 251 nsew signal output
rlabel metal3 s 0 518168 800 518288 6 la_data_out[95]
port 252 nsew signal output
rlabel metal2 s 220266 0 220322 800 6 la_data_out[96]
port 253 nsew signal output
rlabel metal3 s 0 26528 800 26648 6 la_data_out[97]
port 254 nsew signal output
rlabel metal3 s 563200 321648 564000 321768 6 la_data_out[98]
port 255 nsew signal output
rlabel metal3 s 0 578008 800 578128 6 la_data_out[99]
port 256 nsew signal output
rlabel metal2 s 452750 0 452806 800 6 la_data_out[9]
port 257 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 la_oenb[0]
port 258 nsew signal input
rlabel metal3 s 563200 15648 564000 15768 6 la_oenb[100]
port 259 nsew signal input
rlabel metal3 s 563200 414808 564000 414928 6 la_oenb[101]
port 260 nsew signal input
rlabel metal2 s 416042 683200 416098 684000 6 la_oenb[102]
port 261 nsew signal input
rlabel metal3 s 563200 341368 564000 341488 6 la_oenb[103]
port 262 nsew signal input
rlabel metal3 s 0 505248 800 505368 6 la_oenb[104]
port 263 nsew signal input
rlabel metal3 s 0 371968 800 372088 6 la_oenb[105]
port 264 nsew signal input
rlabel metal3 s 563200 82288 564000 82408 6 la_oenb[106]
port 265 nsew signal input
rlabel metal2 s 365810 683200 365866 684000 6 la_oenb[107]
port 266 nsew signal input
rlabel metal2 s 540978 0 541034 800 6 la_oenb[108]
port 267 nsew signal input
rlabel metal2 s 31574 683200 31630 684000 6 la_oenb[109]
port 268 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_oenb[10]
port 269 nsew signal input
rlabel metal3 s 563200 334568 564000 334688 6 la_oenb[110]
port 270 nsew signal input
rlabel metal3 s 0 657568 800 657688 6 la_oenb[111]
port 271 nsew signal input
rlabel metal3 s 563200 434528 564000 434648 6 la_oenb[112]
port 272 nsew signal input
rlabel metal2 s 150714 0 150770 800 6 la_oenb[113]
port 273 nsew signal input
rlabel metal2 s 560298 0 560354 800 6 la_oenb[114]
port 274 nsew signal input
rlabel metal2 s 182914 683200 182970 684000 6 la_oenb[115]
port 275 nsew signal input
rlabel metal2 s 516506 683200 516562 684000 6 la_oenb[116]
port 276 nsew signal input
rlabel metal3 s 563200 501168 564000 501288 6 la_oenb[117]
port 277 nsew signal input
rlabel metal2 s 157798 683200 157854 684000 6 la_oenb[118]
port 278 nsew signal input
rlabel metal2 s 208030 683200 208086 684000 6 la_oenb[119]
port 279 nsew signal input
rlabel metal3 s 563200 135328 564000 135448 6 la_oenb[11]
port 280 nsew signal input
rlabel metal3 s 0 338648 800 338768 6 la_oenb[120]
port 281 nsew signal input
rlabel metal3 s 0 305328 800 305448 6 la_oenb[121]
port 282 nsew signal input
rlabel metal2 s 396722 683200 396778 684000 6 la_oenb[122]
port 283 nsew signal input
rlabel metal2 s 271142 683200 271198 684000 6 la_oenb[123]
port 284 nsew signal input
rlabel metal2 s 38014 683200 38070 684000 6 la_oenb[124]
port 285 nsew signal input
rlabel metal3 s 0 252288 800 252408 6 la_oenb[125]
port 286 nsew signal input
rlabel metal3 s 0 597728 800 597848 6 la_oenb[126]
port 287 nsew signal input
rlabel metal3 s 563200 487568 564000 487688 6 la_oenb[127]
port 288 nsew signal input
rlabel metal3 s 563200 447448 564000 447568 6 la_oenb[12]
port 289 nsew signal input
rlabel metal2 s 377402 0 377458 800 6 la_oenb[13]
port 290 nsew signal input
rlabel metal3 s 563200 408008 564000 408128 6 la_oenb[14]
port 291 nsew signal input
rlabel metal3 s 0 312128 800 312248 6 la_oenb[15]
port 292 nsew signal input
rlabel metal3 s 563200 8848 564000 8968 6 la_oenb[16]
port 293 nsew signal input
rlabel metal2 s 378046 683200 378102 684000 6 la_oenb[17]
port 294 nsew signal input
rlabel metal2 s 548062 683200 548118 684000 6 la_oenb[18]
port 295 nsew signal input
rlabel metal2 s 333610 0 333666 800 6 la_oenb[19]
port 296 nsew signal input
rlabel metal3 s 0 178848 800 178968 6 la_oenb[1]
port 297 nsew signal input
rlabel metal3 s 563200 175448 564000 175568 6 la_oenb[20]
port 298 nsew signal input
rlabel metal2 s 69570 683200 69626 684000 6 la_oenb[21]
port 299 nsew signal input
rlabel metal3 s 0 119008 800 119128 6 la_oenb[22]
port 300 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_oenb[23]
port 301 nsew signal input
rlabel metal2 s 195794 683200 195850 684000 6 la_oenb[24]
port 302 nsew signal input
rlabel metal3 s 0 245488 800 245608 6 la_oenb[25]
port 303 nsew signal input
rlabel metal3 s 563200 633768 564000 633888 6 la_oenb[26]
port 304 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 la_oenb[27]
port 305 nsew signal input
rlabel metal2 s 459834 683200 459890 684000 6 la_oenb[28]
port 306 nsew signal input
rlabel metal3 s 563200 301248 564000 301368 6 la_oenb[29]
port 307 nsew signal input
rlabel metal2 s 465630 0 465686 800 6 la_oenb[2]
port 308 nsew signal input
rlabel metal3 s 0 272008 800 272128 6 la_oenb[30]
port 309 nsew signal input
rlabel metal2 s 446954 0 447010 800 6 la_oenb[31]
port 310 nsew signal input
rlabel metal3 s 0 331848 800 331968 6 la_oenb[32]
port 311 nsew signal input
rlabel metal3 s 0 438608 800 438728 6 la_oenb[33]
port 312 nsew signal input
rlabel metal3 s 563200 35368 564000 35488 6 la_oenb[34]
port 313 nsew signal input
rlabel metal3 s 563200 208088 564000 208208 6 la_oenb[35]
port 314 nsew signal input
rlabel metal2 s 176474 683200 176530 684000 6 la_oenb[36]
port 315 nsew signal input
rlabel metal3 s 563200 580728 564000 580848 6 la_oenb[37]
port 316 nsew signal input
rlabel metal3 s 0 524968 800 525088 6 la_oenb[38]
port 317 nsew signal input
rlabel metal3 s 0 571208 800 571328 6 la_oenb[39]
port 318 nsew signal input
rlabel metal3 s 0 551488 800 551608 6 la_oenb[3]
port 319 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 la_oenb[40]
port 320 nsew signal input
rlabel metal3 s 0 146208 800 146328 6 la_oenb[41]
port 321 nsew signal input
rlabel metal3 s 563200 367888 564000 368008 6 la_oenb[42]
port 322 nsew signal input
rlabel metal2 s 345846 0 345902 800 6 la_oenb[43]
port 323 nsew signal input
rlabel metal2 s 390926 683200 390982 684000 6 la_oenb[44]
port 324 nsew signal input
rlabel metal2 s 535826 683200 535882 684000 6 la_oenb[45]
port 325 nsew signal input
rlabel metal2 s 12898 683200 12954 684000 6 la_oenb[46]
port 326 nsew signal input
rlabel metal3 s 0 292408 800 292528 6 la_oenb[47]
port 327 nsew signal input
rlabel metal3 s 0 325728 800 325848 6 la_oenb[48]
port 328 nsew signal input
rlabel metal2 s 554502 683200 554558 684000 6 la_oenb[49]
port 329 nsew signal input
rlabel metal3 s 0 405288 800 405408 6 la_oenb[4]
port 330 nsew signal input
rlabel metal3 s 0 92488 800 92608 6 la_oenb[50]
port 331 nsew signal input
rlabel metal3 s 563200 241408 564000 241528 6 la_oenb[51]
port 332 nsew signal input
rlabel metal2 s 415398 0 415454 800 6 la_oenb[52]
port 333 nsew signal input
rlabel metal2 s 479154 683200 479210 684000 6 la_oenb[53]
port 334 nsew signal input
rlabel metal2 s 119802 683200 119858 684000 6 la_oenb[54]
port 335 nsew signal input
rlabel metal2 s 188710 0 188766 800 6 la_oenb[55]
port 336 nsew signal input
rlabel metal3 s 563200 420928 564000 421048 6 la_oenb[56]
port 337 nsew signal input
rlabel metal2 s 490746 0 490802 800 6 la_oenb[57]
port 338 nsew signal input
rlabel metal3 s 563200 228488 564000 228608 6 la_oenb[58]
port 339 nsew signal input
rlabel metal3 s 0 358368 800 358488 6 la_oenb[59]
port 340 nsew signal input
rlabel metal3 s 563200 61888 564000 62008 6 la_oenb[5]
port 341 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_oenb[60]
port 342 nsew signal input
rlabel metal2 s 295614 0 295670 800 6 la_oenb[61]
port 343 nsew signal input
rlabel metal3 s 563200 314848 564000 314968 6 la_oenb[62]
port 344 nsew signal input
rlabel metal2 s 447598 683200 447654 684000 6 la_oenb[63]
port 345 nsew signal input
rlabel metal3 s 563200 607248 564000 607368 6 la_oenb[64]
port 346 nsew signal input
rlabel metal3 s 563200 75488 564000 75608 6 la_oenb[65]
port 347 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_oenb[66]
port 348 nsew signal input
rlabel metal3 s 563200 401208 564000 401328 6 la_oenb[67]
port 349 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 la_oenb[68]
port 350 nsew signal input
rlabel metal3 s 563200 626968 564000 627088 6 la_oenb[69]
port 351 nsew signal input
rlabel metal2 s 422482 683200 422538 684000 6 la_oenb[6]
port 352 nsew signal input
rlabel metal3 s 563200 115608 564000 115728 6 la_oenb[70]
port 353 nsew signal input
rlabel metal2 s 403162 683200 403218 684000 6 la_oenb[71]
port 354 nsew signal input
rlabel metal2 s 408958 0 409014 800 6 la_oenb[72]
port 355 nsew signal input
rlabel metal3 s 0 212168 800 212288 6 la_oenb[73]
port 356 nsew signal input
rlabel metal2 s 402518 0 402574 800 6 la_oenb[74]
port 357 nsew signal input
rlabel metal2 s 18 0 74 800 6 la_oenb[75]
port 358 nsew signal input
rlabel metal2 s 478510 0 478566 800 6 la_oenb[76]
port 359 nsew signal input
rlabel metal3 s 0 318928 800 319048 6 la_oenb[77]
port 360 nsew signal input
rlabel metal3 s 0 565088 800 565208 6 la_oenb[78]
port 361 nsew signal input
rlabel metal2 s 132682 683200 132738 684000 6 la_oenb[79]
port 362 nsew signal input
rlabel metal3 s 0 218968 800 219088 6 la_oenb[7]
port 363 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 la_oenb[80]
port 364 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 la_oenb[81]
port 365 nsew signal input
rlabel metal2 s 277582 683200 277638 684000 6 la_oenb[82]
port 366 nsew signal input
rlabel metal2 s 144918 683200 144974 684000 6 la_oenb[83]
port 367 nsew signal input
rlabel metal2 s 327170 0 327226 800 6 la_oenb[84]
port 368 nsew signal input
rlabel metal2 s 384486 683200 384542 684000 6 la_oenb[85]
port 369 nsew signal input
rlabel metal3 s 563200 221688 564000 221808 6 la_oenb[86]
port 370 nsew signal input
rlabel metal3 s 0 425008 800 425128 6 la_oenb[87]
port 371 nsew signal input
rlabel metal3 s 563200 534488 564000 534608 6 la_oenb[88]
port 372 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 la_oenb[89]
port 373 nsew signal input
rlabel metal2 s 232502 0 232558 800 6 la_oenb[8]
port 374 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 la_oenb[90]
port 375 nsew signal input
rlabel metal3 s 563200 514088 564000 514208 6 la_oenb[91]
port 376 nsew signal input
rlabel metal2 s 365166 0 365222 800 6 la_oenb[92]
port 377 nsew signal input
rlabel metal2 s 359370 683200 359426 684000 6 la_oenb[93]
port 378 nsew signal input
rlabel metal2 s 352930 683200 352986 684000 6 la_oenb[94]
port 379 nsew signal input
rlabel metal3 s 0 591608 800 591728 6 la_oenb[95]
port 380 nsew signal input
rlabel metal2 s 25778 683200 25834 684000 6 la_oenb[96]
port 381 nsew signal input
rlabel metal2 s 440514 0 440570 800 6 la_oenb[97]
port 382 nsew signal input
rlabel metal3 s 0 139408 800 139528 6 la_oenb[98]
port 383 nsew signal input
rlabel metal3 s 0 531768 800 531888 6 la_oenb[99]
port 384 nsew signal input
rlabel metal3 s 563200 361088 564000 361208 6 la_oenb[9]
port 385 nsew signal input
rlabel metal4 s 4208 2128 4528 681680 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 681680 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 681680 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 681680 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 681680 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 681680 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 681680 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 681680 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 681680 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 681680 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 681680 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 681680 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 681680 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 681680 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 681680 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 681680 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 681680 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 681680 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 557168 2128 557488 681680 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 681680 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 681680 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 681680 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 681680 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 681680 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 681680 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 681680 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 681680 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 681680 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 681680 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 681680 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 681680 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 681680 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 681680 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 681680 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 681680 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 681680 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 541808 2128 542128 681680 6 vssd1
port 387 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 564000 684000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 170997486
string GDS_FILE /home/drewarosa/RISC-V-Single-Cycle-CPU-Core/openlane/RISC_V/runs/22_09_21_14_02/results/signoff/RISC_V.magic.gds
string GDS_START 1198964
<< end >>

