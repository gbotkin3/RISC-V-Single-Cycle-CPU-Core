magic
tech sky130B
magscale 1 2
timestamp 1663362282
<< obsli1 >>
rect 1104 2159 160448 161041
<< obsm1 >>
rect 14 2128 161078 161220
<< metal2 >>
rect 1306 162936 1362 163736
rect 3238 162936 3294 163736
rect 5814 162936 5870 163736
rect 8390 162936 8446 163736
rect 10322 162936 10378 163736
rect 12898 162936 12954 163736
rect 15474 162936 15530 163736
rect 17406 162936 17462 163736
rect 19982 162936 20038 163736
rect 21914 162936 21970 163736
rect 24490 162936 24546 163736
rect 27066 162936 27122 163736
rect 28998 162936 29054 163736
rect 31574 162936 31630 163736
rect 34150 162936 34206 163736
rect 36082 162936 36138 163736
rect 38658 162936 38714 163736
rect 41234 162936 41290 163736
rect 43166 162936 43222 163736
rect 45742 162936 45798 163736
rect 47674 162936 47730 163736
rect 50250 162936 50306 163736
rect 52826 162936 52882 163736
rect 54758 162936 54814 163736
rect 57334 162936 57390 163736
rect 59910 162936 59966 163736
rect 61842 162936 61898 163736
rect 64418 162936 64474 163736
rect 66350 162936 66406 163736
rect 68926 162936 68982 163736
rect 71502 162936 71558 163736
rect 73434 162936 73490 163736
rect 76010 162936 76066 163736
rect 78586 162936 78642 163736
rect 80518 162936 80574 163736
rect 83094 162936 83150 163736
rect 85026 162936 85082 163736
rect 87602 162936 87658 163736
rect 90178 162936 90234 163736
rect 92110 162936 92166 163736
rect 94686 162936 94742 163736
rect 97262 162936 97318 163736
rect 99194 162936 99250 163736
rect 101770 162936 101826 163736
rect 104346 162936 104402 163736
rect 106278 162936 106334 163736
rect 108854 162936 108910 163736
rect 110786 162936 110842 163736
rect 113362 162936 113418 163736
rect 115938 162936 115994 163736
rect 117870 162936 117926 163736
rect 120446 162936 120502 163736
rect 123022 162936 123078 163736
rect 124954 162936 125010 163736
rect 127530 162936 127586 163736
rect 129462 162936 129518 163736
rect 132038 162936 132094 163736
rect 134614 162936 134670 163736
rect 136546 162936 136602 163736
rect 139122 162936 139178 163736
rect 141698 162936 141754 163736
rect 143630 162936 143686 163736
rect 146206 162936 146262 163736
rect 148782 162936 148838 163736
rect 150714 162936 150770 163736
rect 153290 162936 153346 163736
rect 155222 162936 155278 163736
rect 157798 162936 157854 163736
rect 160374 162936 160430 163736
rect 18 0 74 800
rect 1950 0 2006 800
rect 4526 0 4582 800
rect 6458 0 6514 800
rect 9034 0 9090 800
rect 11610 0 11666 800
rect 13542 0 13598 800
rect 16118 0 16174 800
rect 18694 0 18750 800
rect 20626 0 20682 800
rect 23202 0 23258 800
rect 25134 0 25190 800
rect 27710 0 27766 800
rect 30286 0 30342 800
rect 32218 0 32274 800
rect 34794 0 34850 800
rect 37370 0 37426 800
rect 39302 0 39358 800
rect 41878 0 41934 800
rect 43810 0 43866 800
rect 46386 0 46442 800
rect 48962 0 49018 800
rect 50894 0 50950 800
rect 53470 0 53526 800
rect 56046 0 56102 800
rect 57978 0 58034 800
rect 60554 0 60610 800
rect 63130 0 63186 800
rect 65062 0 65118 800
rect 67638 0 67694 800
rect 69570 0 69626 800
rect 72146 0 72202 800
rect 74722 0 74778 800
rect 76654 0 76710 800
rect 79230 0 79286 800
rect 81806 0 81862 800
rect 83738 0 83794 800
rect 86314 0 86370 800
rect 88246 0 88302 800
rect 90822 0 90878 800
rect 93398 0 93454 800
rect 95330 0 95386 800
rect 97906 0 97962 800
rect 100482 0 100538 800
rect 102414 0 102470 800
rect 104990 0 105046 800
rect 107566 0 107622 800
rect 109498 0 109554 800
rect 112074 0 112130 800
rect 114006 0 114062 800
rect 116582 0 116638 800
rect 119158 0 119214 800
rect 121090 0 121146 800
rect 123666 0 123722 800
rect 126242 0 126298 800
rect 128174 0 128230 800
rect 130750 0 130806 800
rect 132682 0 132738 800
rect 135258 0 135314 800
rect 137834 0 137890 800
rect 139766 0 139822 800
rect 142342 0 142398 800
rect 144918 0 144974 800
rect 146850 0 146906 800
rect 149426 0 149482 800
rect 152002 0 152058 800
rect 153934 0 153990 800
rect 156510 0 156566 800
rect 158442 0 158498 800
rect 161018 0 161074 800
<< obsm2 >>
rect 20 162880 1250 163010
rect 1418 162880 3182 163010
rect 3350 162880 5758 163010
rect 5926 162880 8334 163010
rect 8502 162880 10266 163010
rect 10434 162880 12842 163010
rect 13010 162880 15418 163010
rect 15586 162880 17350 163010
rect 17518 162880 19926 163010
rect 20094 162880 21858 163010
rect 22026 162880 24434 163010
rect 24602 162880 27010 163010
rect 27178 162880 28942 163010
rect 29110 162880 31518 163010
rect 31686 162880 34094 163010
rect 34262 162880 36026 163010
rect 36194 162880 38602 163010
rect 38770 162880 41178 163010
rect 41346 162880 43110 163010
rect 43278 162880 45686 163010
rect 45854 162880 47618 163010
rect 47786 162880 50194 163010
rect 50362 162880 52770 163010
rect 52938 162880 54702 163010
rect 54870 162880 57278 163010
rect 57446 162880 59854 163010
rect 60022 162880 61786 163010
rect 61954 162880 64362 163010
rect 64530 162880 66294 163010
rect 66462 162880 68870 163010
rect 69038 162880 71446 163010
rect 71614 162880 73378 163010
rect 73546 162880 75954 163010
rect 76122 162880 78530 163010
rect 78698 162880 80462 163010
rect 80630 162880 83038 163010
rect 83206 162880 84970 163010
rect 85138 162880 87546 163010
rect 87714 162880 90122 163010
rect 90290 162880 92054 163010
rect 92222 162880 94630 163010
rect 94798 162880 97206 163010
rect 97374 162880 99138 163010
rect 99306 162880 101714 163010
rect 101882 162880 104290 163010
rect 104458 162880 106222 163010
rect 106390 162880 108798 163010
rect 108966 162880 110730 163010
rect 110898 162880 113306 163010
rect 113474 162880 115882 163010
rect 116050 162880 117814 163010
rect 117982 162880 120390 163010
rect 120558 162880 122966 163010
rect 123134 162880 124898 163010
rect 125066 162880 127474 163010
rect 127642 162880 129406 163010
rect 129574 162880 131982 163010
rect 132150 162880 134558 163010
rect 134726 162880 136490 163010
rect 136658 162880 139066 163010
rect 139234 162880 141642 163010
rect 141810 162880 143574 163010
rect 143742 162880 146150 163010
rect 146318 162880 148726 163010
rect 148894 162880 150658 163010
rect 150826 162880 153234 163010
rect 153402 162880 155166 163010
rect 155334 162880 157742 163010
rect 157910 162880 160318 163010
rect 160486 162880 161072 163010
rect 20 856 161072 162880
rect 130 800 1894 856
rect 2062 800 4470 856
rect 4638 800 6402 856
rect 6570 800 8978 856
rect 9146 800 11554 856
rect 11722 800 13486 856
rect 13654 800 16062 856
rect 16230 800 18638 856
rect 18806 800 20570 856
rect 20738 800 23146 856
rect 23314 800 25078 856
rect 25246 800 27654 856
rect 27822 800 30230 856
rect 30398 800 32162 856
rect 32330 800 34738 856
rect 34906 800 37314 856
rect 37482 800 39246 856
rect 39414 800 41822 856
rect 41990 800 43754 856
rect 43922 800 46330 856
rect 46498 800 48906 856
rect 49074 800 50838 856
rect 51006 800 53414 856
rect 53582 800 55990 856
rect 56158 800 57922 856
rect 58090 800 60498 856
rect 60666 800 63074 856
rect 63242 800 65006 856
rect 65174 800 67582 856
rect 67750 800 69514 856
rect 69682 800 72090 856
rect 72258 800 74666 856
rect 74834 800 76598 856
rect 76766 800 79174 856
rect 79342 800 81750 856
rect 81918 800 83682 856
rect 83850 800 86258 856
rect 86426 800 88190 856
rect 88358 800 90766 856
rect 90934 800 93342 856
rect 93510 800 95274 856
rect 95442 800 97850 856
rect 98018 800 100426 856
rect 100594 800 102358 856
rect 102526 800 104934 856
rect 105102 800 107510 856
rect 107678 800 109442 856
rect 109610 800 112018 856
rect 112186 800 113950 856
rect 114118 800 116526 856
rect 116694 800 119102 856
rect 119270 800 121034 856
rect 121202 800 123610 856
rect 123778 800 126186 856
rect 126354 800 128118 856
rect 128286 800 130694 856
rect 130862 800 132626 856
rect 132794 800 135202 856
rect 135370 800 137778 856
rect 137946 800 139710 856
rect 139878 800 142286 856
rect 142454 800 144862 856
rect 145030 800 146794 856
rect 146962 800 149370 856
rect 149538 800 151946 856
rect 152114 800 153878 856
rect 154046 800 156454 856
rect 156622 800 158386 856
rect 158554 800 160962 856
<< metal3 >>
rect 0 162528 800 162648
rect 160792 162528 161592 162648
rect 0 160488 800 160608
rect 160792 159808 161592 159928
rect 0 157768 800 157888
rect 160792 157088 161592 157208
rect 0 155048 800 155168
rect 160792 155048 161592 155168
rect 0 153008 800 153128
rect 160792 152328 161592 152448
rect 0 150288 800 150408
rect 160792 150288 161592 150408
rect 0 147568 800 147688
rect 160792 147568 161592 147688
rect 0 145528 800 145648
rect 160792 144848 161592 144968
rect 0 142808 800 142928
rect 160792 142808 161592 142928
rect 0 140088 800 140208
rect 160792 140088 161592 140208
rect 0 138048 800 138168
rect 160792 137368 161592 137488
rect 0 135328 800 135448
rect 160792 135328 161592 135448
rect 0 133288 800 133408
rect 160792 132608 161592 132728
rect 0 130568 800 130688
rect 160792 129888 161592 130008
rect 0 127848 800 127968
rect 160792 127848 161592 127968
rect 0 125808 800 125928
rect 160792 125128 161592 125248
rect 0 123088 800 123208
rect 160792 123088 161592 123208
rect 0 120368 800 120488
rect 160792 120368 161592 120488
rect 0 118328 800 118448
rect 160792 117648 161592 117768
rect 0 115608 800 115728
rect 160792 115608 161592 115728
rect 0 113568 800 113688
rect 160792 112888 161592 113008
rect 0 110848 800 110968
rect 160792 110168 161592 110288
rect 0 108128 800 108248
rect 160792 108128 161592 108248
rect 0 106088 800 106208
rect 160792 105408 161592 105528
rect 0 103368 800 103488
rect 160792 103368 161592 103488
rect 0 100648 800 100768
rect 160792 100648 161592 100768
rect 0 98608 800 98728
rect 160792 97928 161592 98048
rect 0 95888 800 96008
rect 160792 95888 161592 96008
rect 0 93168 800 93288
rect 160792 93168 161592 93288
rect 0 91128 800 91248
rect 160792 90448 161592 90568
rect 0 88408 800 88528
rect 160792 88408 161592 88528
rect 0 86368 800 86488
rect 160792 85688 161592 85808
rect 0 83648 800 83768
rect 160792 82968 161592 83088
rect 0 80928 800 81048
rect 160792 80928 161592 81048
rect 0 78888 800 79008
rect 160792 78208 161592 78328
rect 0 76168 800 76288
rect 160792 76168 161592 76288
rect 0 73448 800 73568
rect 160792 73448 161592 73568
rect 0 71408 800 71528
rect 160792 70728 161592 70848
rect 0 68688 800 68808
rect 160792 68688 161592 68808
rect 0 66648 800 66768
rect 160792 65968 161592 66088
rect 0 63928 800 64048
rect 160792 63248 161592 63368
rect 0 61208 800 61328
rect 160792 61208 161592 61328
rect 0 59168 800 59288
rect 160792 58488 161592 58608
rect 0 56448 800 56568
rect 160792 56448 161592 56568
rect 0 53728 800 53848
rect 160792 53728 161592 53848
rect 0 51688 800 51808
rect 160792 51008 161592 51128
rect 0 48968 800 49088
rect 160792 48968 161592 49088
rect 0 46248 800 46368
rect 160792 46248 161592 46368
rect 0 44208 800 44328
rect 160792 43528 161592 43648
rect 0 41488 800 41608
rect 160792 41488 161592 41608
rect 0 39448 800 39568
rect 160792 38768 161592 38888
rect 0 36728 800 36848
rect 160792 36728 161592 36848
rect 0 34008 800 34128
rect 160792 34008 161592 34128
rect 0 31968 800 32088
rect 160792 31288 161592 31408
rect 0 29248 800 29368
rect 160792 29248 161592 29368
rect 0 26528 800 26648
rect 160792 26528 161592 26648
rect 0 24488 800 24608
rect 160792 23808 161592 23928
rect 0 21768 800 21888
rect 160792 21768 161592 21888
rect 0 19728 800 19848
rect 160792 19048 161592 19168
rect 0 17008 800 17128
rect 160792 16328 161592 16448
rect 0 14288 800 14408
rect 160792 14288 161592 14408
rect 0 12248 800 12368
rect 160792 11568 161592 11688
rect 0 9528 800 9648
rect 160792 9528 161592 9648
rect 0 6808 800 6928
rect 160792 6808 161592 6928
rect 0 4768 800 4888
rect 160792 4088 161592 4208
rect 0 2048 800 2168
rect 160792 2048 161592 2168
<< obsm3 >>
rect 880 162448 160712 162621
rect 800 160688 160792 162448
rect 880 160408 160792 160688
rect 800 160008 160792 160408
rect 800 159728 160712 160008
rect 800 157968 160792 159728
rect 880 157688 160792 157968
rect 800 157288 160792 157688
rect 800 157008 160712 157288
rect 800 155248 160792 157008
rect 880 154968 160712 155248
rect 800 153208 160792 154968
rect 880 152928 160792 153208
rect 800 152528 160792 152928
rect 800 152248 160712 152528
rect 800 150488 160792 152248
rect 880 150208 160712 150488
rect 800 147768 160792 150208
rect 880 147488 160712 147768
rect 800 145728 160792 147488
rect 880 145448 160792 145728
rect 800 145048 160792 145448
rect 800 144768 160712 145048
rect 800 143008 160792 144768
rect 880 142728 160712 143008
rect 800 140288 160792 142728
rect 880 140008 160712 140288
rect 800 138248 160792 140008
rect 880 137968 160792 138248
rect 800 137568 160792 137968
rect 800 137288 160712 137568
rect 800 135528 160792 137288
rect 880 135248 160712 135528
rect 800 133488 160792 135248
rect 880 133208 160792 133488
rect 800 132808 160792 133208
rect 800 132528 160712 132808
rect 800 130768 160792 132528
rect 880 130488 160792 130768
rect 800 130088 160792 130488
rect 800 129808 160712 130088
rect 800 128048 160792 129808
rect 880 127768 160712 128048
rect 800 126008 160792 127768
rect 880 125728 160792 126008
rect 800 125328 160792 125728
rect 800 125048 160712 125328
rect 800 123288 160792 125048
rect 880 123008 160712 123288
rect 800 120568 160792 123008
rect 880 120288 160712 120568
rect 800 118528 160792 120288
rect 880 118248 160792 118528
rect 800 117848 160792 118248
rect 800 117568 160712 117848
rect 800 115808 160792 117568
rect 880 115528 160712 115808
rect 800 113768 160792 115528
rect 880 113488 160792 113768
rect 800 113088 160792 113488
rect 800 112808 160712 113088
rect 800 111048 160792 112808
rect 880 110768 160792 111048
rect 800 110368 160792 110768
rect 800 110088 160712 110368
rect 800 108328 160792 110088
rect 880 108048 160712 108328
rect 800 106288 160792 108048
rect 880 106008 160792 106288
rect 800 105608 160792 106008
rect 800 105328 160712 105608
rect 800 103568 160792 105328
rect 880 103288 160712 103568
rect 800 100848 160792 103288
rect 880 100568 160712 100848
rect 800 98808 160792 100568
rect 880 98528 160792 98808
rect 800 98128 160792 98528
rect 800 97848 160712 98128
rect 800 96088 160792 97848
rect 880 95808 160712 96088
rect 800 93368 160792 95808
rect 880 93088 160712 93368
rect 800 91328 160792 93088
rect 880 91048 160792 91328
rect 800 90648 160792 91048
rect 800 90368 160712 90648
rect 800 88608 160792 90368
rect 880 88328 160712 88608
rect 800 86568 160792 88328
rect 880 86288 160792 86568
rect 800 85888 160792 86288
rect 800 85608 160712 85888
rect 800 83848 160792 85608
rect 880 83568 160792 83848
rect 800 83168 160792 83568
rect 800 82888 160712 83168
rect 800 81128 160792 82888
rect 880 80848 160712 81128
rect 800 79088 160792 80848
rect 880 78808 160792 79088
rect 800 78408 160792 78808
rect 800 78128 160712 78408
rect 800 76368 160792 78128
rect 880 76088 160712 76368
rect 800 73648 160792 76088
rect 880 73368 160712 73648
rect 800 71608 160792 73368
rect 880 71328 160792 71608
rect 800 70928 160792 71328
rect 800 70648 160712 70928
rect 800 68888 160792 70648
rect 880 68608 160712 68888
rect 800 66848 160792 68608
rect 880 66568 160792 66848
rect 800 66168 160792 66568
rect 800 65888 160712 66168
rect 800 64128 160792 65888
rect 880 63848 160792 64128
rect 800 63448 160792 63848
rect 800 63168 160712 63448
rect 800 61408 160792 63168
rect 880 61128 160712 61408
rect 800 59368 160792 61128
rect 880 59088 160792 59368
rect 800 58688 160792 59088
rect 800 58408 160712 58688
rect 800 56648 160792 58408
rect 880 56368 160712 56648
rect 800 53928 160792 56368
rect 880 53648 160712 53928
rect 800 51888 160792 53648
rect 880 51608 160792 51888
rect 800 51208 160792 51608
rect 800 50928 160712 51208
rect 800 49168 160792 50928
rect 880 48888 160712 49168
rect 800 46448 160792 48888
rect 880 46168 160712 46448
rect 800 44408 160792 46168
rect 880 44128 160792 44408
rect 800 43728 160792 44128
rect 800 43448 160712 43728
rect 800 41688 160792 43448
rect 880 41408 160712 41688
rect 800 39648 160792 41408
rect 880 39368 160792 39648
rect 800 38968 160792 39368
rect 800 38688 160712 38968
rect 800 36928 160792 38688
rect 880 36648 160712 36928
rect 800 34208 160792 36648
rect 880 33928 160712 34208
rect 800 32168 160792 33928
rect 880 31888 160792 32168
rect 800 31488 160792 31888
rect 800 31208 160712 31488
rect 800 29448 160792 31208
rect 880 29168 160712 29448
rect 800 26728 160792 29168
rect 880 26448 160712 26728
rect 800 24688 160792 26448
rect 880 24408 160792 24688
rect 800 24008 160792 24408
rect 800 23728 160712 24008
rect 800 21968 160792 23728
rect 880 21688 160712 21968
rect 800 19928 160792 21688
rect 880 19648 160792 19928
rect 800 19248 160792 19648
rect 800 18968 160712 19248
rect 800 17208 160792 18968
rect 880 16928 160792 17208
rect 800 16528 160792 16928
rect 800 16248 160712 16528
rect 800 14488 160792 16248
rect 880 14208 160712 14488
rect 800 12448 160792 14208
rect 880 12168 160792 12448
rect 800 11768 160792 12168
rect 800 11488 160712 11768
rect 800 9728 160792 11488
rect 880 9448 160712 9728
rect 800 7008 160792 9448
rect 880 6728 160712 7008
rect 800 4968 160792 6728
rect 880 4688 160792 4968
rect 800 4288 160792 4688
rect 800 4008 160712 4288
rect 800 2248 160792 4008
rect 880 1968 160712 2248
rect 800 1667 160792 1968
<< metal4 >>
rect 4208 2128 4528 161072
rect 19568 2128 19888 161072
rect 34928 2128 35248 161072
rect 50288 2128 50608 161072
rect 65648 2128 65968 161072
rect 81008 2128 81328 161072
rect 96368 2128 96688 161072
rect 111728 2128 112048 161072
rect 127088 2128 127408 161072
rect 142448 2128 142768 161072
rect 157808 2128 158128 161072
<< obsm4 >>
rect 22323 2048 34848 160173
rect 35328 2048 50208 160173
rect 50688 2048 65568 160173
rect 66048 2048 80928 160173
rect 81408 2048 96288 160173
rect 96768 2048 111648 160173
rect 112128 2048 116413 160173
rect 22323 1667 116413 2048
<< labels >>
rlabel metal2 s 57334 162936 57390 163736 6 alu_output[0]
port 1 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 alu_output[10]
port 2 nsew signal output
rlabel metal2 s 27066 162936 27122 163736 6 alu_output[11]
port 3 nsew signal output
rlabel metal2 s 12898 162936 12954 163736 6 alu_output[12]
port 4 nsew signal output
rlabel metal2 s 36082 162936 36138 163736 6 alu_output[13]
port 5 nsew signal output
rlabel metal2 s 115938 162936 115994 163736 6 alu_output[14]
port 6 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 alu_output[15]
port 7 nsew signal output
rlabel metal3 s 0 59168 800 59288 6 alu_output[16]
port 8 nsew signal output
rlabel metal3 s 160792 48968 161592 49088 6 alu_output[17]
port 9 nsew signal output
rlabel metal2 s 123022 162936 123078 163736 6 alu_output[18]
port 10 nsew signal output
rlabel metal3 s 160792 26528 161592 26648 6 alu_output[19]
port 11 nsew signal output
rlabel metal2 s 126242 0 126298 800 6 alu_output[1]
port 12 nsew signal output
rlabel metal3 s 160792 95888 161592 96008 6 alu_output[20]
port 13 nsew signal output
rlabel metal2 s 127530 162936 127586 163736 6 alu_output[21]
port 14 nsew signal output
rlabel metal3 s 0 133288 800 133408 6 alu_output[22]
port 15 nsew signal output
rlabel metal3 s 160792 21768 161592 21888 6 alu_output[23]
port 16 nsew signal output
rlabel metal2 s 136546 162936 136602 163736 6 alu_output[24]
port 17 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 alu_output[25]
port 18 nsew signal output
rlabel metal2 s 15474 162936 15530 163736 6 alu_output[26]
port 19 nsew signal output
rlabel metal3 s 160792 140088 161592 140208 6 alu_output[27]
port 20 nsew signal output
rlabel metal3 s 160792 100648 161592 100768 6 alu_output[28]
port 21 nsew signal output
rlabel metal2 s 157798 162936 157854 163736 6 alu_output[29]
port 22 nsew signal output
rlabel metal2 s 78586 162936 78642 163736 6 alu_output[2]
port 23 nsew signal output
rlabel metal3 s 0 115608 800 115728 6 alu_output[30]
port 24 nsew signal output
rlabel metal3 s 160792 2048 161592 2168 6 alu_output[31]
port 25 nsew signal output
rlabel metal2 s 34150 162936 34206 163736 6 alu_output[3]
port 26 nsew signal output
rlabel metal2 s 80518 162936 80574 163736 6 alu_output[4]
port 27 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 alu_output[5]
port 28 nsew signal output
rlabel metal2 s 149426 0 149482 800 6 alu_output[6]
port 29 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 alu_output[7]
port 30 nsew signal output
rlabel metal2 s 97262 162936 97318 163736 6 alu_output[8]
port 31 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 alu_output[9]
port 32 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 clk
port 33 nsew signal input
rlabel metal2 s 90178 162936 90234 163736 6 funct3[0]
port 34 nsew signal input
rlabel metal3 s 160792 82968 161592 83088 6 funct3[1]
port 35 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 funct3[2]
port 36 nsew signal input
rlabel metal3 s 160792 85688 161592 85808 6 funct7[0]
port 37 nsew signal input
rlabel metal3 s 160792 65968 161592 66088 6 funct7[1]
port 38 nsew signal input
rlabel metal3 s 160792 147568 161592 147688 6 funct7[2]
port 39 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 funct7[3]
port 40 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 funct7[4]
port 41 nsew signal input
rlabel metal3 s 0 127848 800 127968 6 funct7[5]
port 42 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 funct7[6]
port 43 nsew signal input
rlabel metal2 s 129462 162936 129518 163736 6 immediate[0]
port 44 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 immediate[10]
port 45 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 immediate[11]
port 46 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 immediate[12]
port 47 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 immediate[13]
port 48 nsew signal input
rlabel metal3 s 0 113568 800 113688 6 immediate[14]
port 49 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 immediate[15]
port 50 nsew signal input
rlabel metal2 s 101770 162936 101826 163736 6 immediate[16]
port 51 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 immediate[17]
port 52 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 immediate[18]
port 53 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 immediate[19]
port 54 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 immediate[1]
port 55 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 immediate[20]
port 56 nsew signal input
rlabel metal3 s 0 86368 800 86488 6 immediate[21]
port 57 nsew signal input
rlabel metal2 s 76010 162936 76066 163736 6 immediate[22]
port 58 nsew signal input
rlabel metal3 s 160792 132608 161592 132728 6 immediate[23]
port 59 nsew signal input
rlabel metal2 s 68926 162936 68982 163736 6 immediate[24]
port 60 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 immediate[25]
port 61 nsew signal input
rlabel metal2 s 87602 162936 87658 163736 6 immediate[26]
port 62 nsew signal input
rlabel metal2 s 10322 162936 10378 163736 6 immediate[27]
port 63 nsew signal input
rlabel metal3 s 0 56448 800 56568 6 immediate[28]
port 64 nsew signal input
rlabel metal2 s 54758 162936 54814 163736 6 immediate[29]
port 65 nsew signal input
rlabel metal3 s 0 140088 800 140208 6 immediate[2]
port 66 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 immediate[30]
port 67 nsew signal input
rlabel metal3 s 160792 9528 161592 9648 6 immediate[31]
port 68 nsew signal input
rlabel metal2 s 66350 162936 66406 163736 6 immediate[3]
port 69 nsew signal input
rlabel metal3 s 0 83648 800 83768 6 immediate[4]
port 70 nsew signal input
rlabel metal2 s 1306 162936 1362 163736 6 immediate[5]
port 71 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 immediate[6]
port 72 nsew signal input
rlabel metal2 s 117870 162936 117926 163736 6 immediate[7]
port 73 nsew signal input
rlabel metal2 s 150714 162936 150770 163736 6 immediate[8]
port 74 nsew signal input
rlabel metal3 s 160792 137368 161592 137488 6 immediate[9]
port 75 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 immediate_sel
port 76 nsew signal input
rlabel metal3 s 160792 76168 161592 76288 6 instruction_type[0]
port 77 nsew signal input
rlabel metal3 s 160792 155048 161592 155168 6 instruction_type[1]
port 78 nsew signal input
rlabel metal3 s 160792 110168 161592 110288 6 instruction_type[2]
port 79 nsew signal input
rlabel metal2 s 17406 162936 17462 163736 6 instruction_type[3]
port 80 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 instruction_type[4]
port 81 nsew signal input
rlabel metal3 s 0 123088 800 123208 6 instruction_type[5]
port 82 nsew signal input
rlabel metal3 s 160792 125128 161592 125248 6 la_read_data[0]
port 83 nsew signal output
rlabel metal2 s 83094 162936 83150 163736 6 la_read_data[10]
port 84 nsew signal output
rlabel metal3 s 0 147568 800 147688 6 la_read_data[11]
port 85 nsew signal output
rlabel metal2 s 144918 0 144974 800 6 la_read_data[12]
port 86 nsew signal output
rlabel metal3 s 0 142808 800 142928 6 la_read_data[13]
port 87 nsew signal output
rlabel metal2 s 8390 162936 8446 163736 6 la_read_data[14]
port 88 nsew signal output
rlabel metal2 s 146850 0 146906 800 6 la_read_data[15]
port 89 nsew signal output
rlabel metal3 s 160792 43528 161592 43648 6 la_read_data[16]
port 90 nsew signal output
rlabel metal3 s 160792 88408 161592 88528 6 la_read_data[17]
port 91 nsew signal output
rlabel metal3 s 160792 90448 161592 90568 6 la_read_data[18]
port 92 nsew signal output
rlabel metal3 s 0 130568 800 130688 6 la_read_data[19]
port 93 nsew signal output
rlabel metal2 s 106278 162936 106334 163736 6 la_read_data[1]
port 94 nsew signal output
rlabel metal2 s 3238 162936 3294 163736 6 la_read_data[20]
port 95 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 la_read_data[21]
port 96 nsew signal output
rlabel metal2 s 142342 0 142398 800 6 la_read_data[22]
port 97 nsew signal output
rlabel metal2 s 132682 0 132738 800 6 la_read_data[23]
port 98 nsew signal output
rlabel metal3 s 0 80928 800 81048 6 la_read_data[24]
port 99 nsew signal output
rlabel metal3 s 0 110848 800 110968 6 la_read_data[25]
port 100 nsew signal output
rlabel metal3 s 0 135328 800 135448 6 la_read_data[26]
port 101 nsew signal output
rlabel metal2 s 158442 0 158498 800 6 la_read_data[27]
port 102 nsew signal output
rlabel metal2 s 45742 162936 45798 163736 6 la_read_data[28]
port 103 nsew signal output
rlabel metal2 s 153290 162936 153346 163736 6 la_read_data[29]
port 104 nsew signal output
rlabel metal2 s 43166 162936 43222 163736 6 la_read_data[2]
port 105 nsew signal output
rlabel metal3 s 160792 159808 161592 159928 6 la_read_data[30]
port 106 nsew signal output
rlabel metal3 s 0 155048 800 155168 6 la_read_data[31]
port 107 nsew signal output
rlabel metal2 s 112074 0 112130 800 6 la_read_data[3]
port 108 nsew signal output
rlabel metal3 s 0 95888 800 96008 6 la_read_data[4]
port 109 nsew signal output
rlabel metal2 s 38658 162936 38714 163736 6 la_read_data[5]
port 110 nsew signal output
rlabel metal2 s 71502 162936 71558 163736 6 la_read_data[6]
port 111 nsew signal output
rlabel metal3 s 160792 80928 161592 81048 6 la_read_data[7]
port 112 nsew signal output
rlabel metal3 s 0 160488 800 160608 6 la_read_data[8]
port 113 nsew signal output
rlabel metal3 s 160792 11568 161592 11688 6 la_read_data[9]
port 114 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 la_reg_select[0]
port 115 nsew signal input
rlabel metal3 s 160792 93168 161592 93288 6 la_reg_select[1]
port 116 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 la_reg_select[2]
port 117 nsew signal input
rlabel metal2 s 50250 162936 50306 163736 6 la_reg_select[3]
port 118 nsew signal input
rlabel metal3 s 0 103368 800 103488 6 la_reg_select[4]
port 119 nsew signal input
rlabel metal3 s 160792 61208 161592 61328 6 opcode[0]
port 120 nsew signal input
rlabel metal3 s 160792 46248 161592 46368 6 opcode[1]
port 121 nsew signal input
rlabel metal3 s 160792 129888 161592 130008 6 opcode[2]
port 122 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 opcode[3]
port 123 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 opcode[4]
port 124 nsew signal input
rlabel metal2 s 47674 162936 47730 163736 6 opcode[5]
port 125 nsew signal input
rlabel metal3 s 0 88408 800 88528 6 opcode[6]
port 126 nsew signal input
rlabel metal3 s 0 68688 800 68808 6 pc[0]
port 127 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 pc[10]
port 128 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 pc[11]
port 129 nsew signal input
rlabel metal2 s 141698 162936 141754 163736 6 pc[12]
port 130 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 pc[13]
port 131 nsew signal input
rlabel metal2 s 61842 162936 61898 163736 6 pc[14]
port 132 nsew signal input
rlabel metal2 s 31574 162936 31630 163736 6 pc[15]
port 133 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 pc[16]
port 134 nsew signal input
rlabel metal3 s 0 108128 800 108248 6 pc[17]
port 135 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 pc[18]
port 136 nsew signal input
rlabel metal3 s 160792 97928 161592 98048 6 pc[19]
port 137 nsew signal input
rlabel metal3 s 0 153008 800 153128 6 pc[1]
port 138 nsew signal input
rlabel metal2 s 5814 162936 5870 163736 6 pc[20]
port 139 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 pc[21]
port 140 nsew signal input
rlabel metal3 s 160792 16328 161592 16448 6 pc[22]
port 141 nsew signal input
rlabel metal3 s 160792 41488 161592 41608 6 pc[23]
port 142 nsew signal input
rlabel metal3 s 0 41488 800 41608 6 pc[24]
port 143 nsew signal input
rlabel metal2 s 155222 162936 155278 163736 6 pc[25]
port 144 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 pc[26]
port 145 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 pc[27]
port 146 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 pc[28]
port 147 nsew signal input
rlabel metal3 s 160792 23808 161592 23928 6 pc[29]
port 148 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 pc[2]
port 149 nsew signal input
rlabel metal3 s 160792 105408 161592 105528 6 pc[30]
port 150 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 pc[31]
port 151 nsew signal input
rlabel metal3 s 0 150288 800 150408 6 pc[3]
port 152 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 pc[4]
port 153 nsew signal input
rlabel metal2 s 104346 162936 104402 163736 6 pc[5]
port 154 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 pc[6]
port 155 nsew signal input
rlabel metal3 s 160792 29248 161592 29368 6 pc[7]
port 156 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 pc[8]
port 157 nsew signal input
rlabel metal3 s 160792 51008 161592 51128 6 pc[9]
port 158 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 rd[0]
port 159 nsew signal input
rlabel metal3 s 0 118328 800 118448 6 rd[1]
port 160 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 rd[2]
port 161 nsew signal input
rlabel metal3 s 160792 117648 161592 117768 6 rd[3]
port 162 nsew signal input
rlabel metal3 s 160792 68688 161592 68808 6 rd[4]
port 163 nsew signal input
rlabel metal2 s 124954 162936 125010 163736 6 read_data[0]
port 164 nsew signal input
rlabel metal2 s 134614 162936 134670 163736 6 read_data[10]
port 165 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 read_data[11]
port 166 nsew signal input
rlabel metal2 s 41234 162936 41290 163736 6 read_data[12]
port 167 nsew signal input
rlabel metal2 s 64418 162936 64474 163736 6 read_data[13]
port 168 nsew signal input
rlabel metal3 s 160792 150288 161592 150408 6 read_data[14]
port 169 nsew signal input
rlabel metal2 s 143630 162936 143686 163736 6 read_data[15]
port 170 nsew signal input
rlabel metal2 s 92110 162936 92166 163736 6 read_data[16]
port 171 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 read_data[17]
port 172 nsew signal input
rlabel metal3 s 0 106088 800 106208 6 read_data[18]
port 173 nsew signal input
rlabel metal3 s 160792 70728 161592 70848 6 read_data[19]
port 174 nsew signal input
rlabel metal3 s 160792 63248 161592 63368 6 read_data[1]
port 175 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 read_data[20]
port 176 nsew signal input
rlabel metal3 s 160792 56448 161592 56568 6 read_data[21]
port 177 nsew signal input
rlabel metal3 s 160792 14288 161592 14408 6 read_data[22]
port 178 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 read_data[23]
port 179 nsew signal input
rlabel metal3 s 160792 162528 161592 162648 6 read_data[24]
port 180 nsew signal input
rlabel metal3 s 160792 123088 161592 123208 6 read_data[25]
port 181 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 read_data[26]
port 182 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 read_data[27]
port 183 nsew signal input
rlabel metal3 s 160792 4088 161592 4208 6 read_data[28]
port 184 nsew signal input
rlabel metal2 s 85026 162936 85082 163736 6 read_data[29]
port 185 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 read_data[2]
port 186 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 read_data[30]
port 187 nsew signal input
rlabel metal2 s 113362 162936 113418 163736 6 read_data[31]
port 188 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 read_data[3]
port 189 nsew signal input
rlabel metal3 s 160792 112888 161592 113008 6 read_data[4]
port 190 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 read_data[5]
port 191 nsew signal input
rlabel metal3 s 160792 152328 161592 152448 6 read_data[6]
port 192 nsew signal input
rlabel metal3 s 160792 36728 161592 36848 6 read_data[7]
port 193 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 read_data[8]
port 194 nsew signal input
rlabel metal3 s 160792 157088 161592 157208 6 read_data[9]
port 195 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 reg_write
port 196 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 rs1[0]
port 197 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 rs1[1]
port 198 nsew signal input
rlabel metal2 s 139766 0 139822 800 6 rs1[2]
port 199 nsew signal input
rlabel metal3 s 160792 19048 161592 19168 6 rs1[3]
port 200 nsew signal input
rlabel metal2 s 99194 162936 99250 163736 6 rs1[4]
port 201 nsew signal input
rlabel metal3 s 160792 108128 161592 108248 6 rs1_data[0]
port 202 nsew signal output
rlabel metal2 s 19982 162936 20038 163736 6 rs1_data[10]
port 203 nsew signal output
rlabel metal2 s 28998 162936 29054 163736 6 rs1_data[11]
port 204 nsew signal output
rlabel metal2 s 24490 162936 24546 163736 6 rs1_data[12]
port 205 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 rs1_data[13]
port 206 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 rs1_data[14]
port 207 nsew signal output
rlabel metal3 s 160792 58488 161592 58608 6 rs1_data[15]
port 208 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 rs1_data[16]
port 209 nsew signal output
rlabel metal2 s 146206 162936 146262 163736 6 rs1_data[17]
port 210 nsew signal output
rlabel metal3 s 160792 144848 161592 144968 6 rs1_data[18]
port 211 nsew signal output
rlabel metal2 s 52826 162936 52882 163736 6 rs1_data[19]
port 212 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 rs1_data[1]
port 213 nsew signal output
rlabel metal3 s 160792 73448 161592 73568 6 rs1_data[20]
port 214 nsew signal output
rlabel metal3 s 160792 142808 161592 142928 6 rs1_data[21]
port 215 nsew signal output
rlabel metal3 s 0 145528 800 145648 6 rs1_data[22]
port 216 nsew signal output
rlabel metal3 s 160792 103368 161592 103488 6 rs1_data[23]
port 217 nsew signal output
rlabel metal3 s 160792 34008 161592 34128 6 rs1_data[24]
port 218 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 rs1_data[25]
port 219 nsew signal output
rlabel metal2 s 160374 162936 160430 163736 6 rs1_data[26]
port 220 nsew signal output
rlabel metal2 s 73434 162936 73490 163736 6 rs1_data[27]
port 221 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 rs1_data[28]
port 222 nsew signal output
rlabel metal3 s 0 91128 800 91248 6 rs1_data[29]
port 223 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 rs1_data[2]
port 224 nsew signal output
rlabel metal3 s 160792 31288 161592 31408 6 rs1_data[30]
port 225 nsew signal output
rlabel metal3 s 0 125808 800 125928 6 rs1_data[31]
port 226 nsew signal output
rlabel metal2 s 153934 0 153990 800 6 rs1_data[3]
port 227 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 rs1_data[4]
port 228 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 rs1_data[5]
port 229 nsew signal output
rlabel metal3 s 160792 53728 161592 53848 6 rs1_data[6]
port 230 nsew signal output
rlabel metal2 s 148782 162936 148838 163736 6 rs1_data[7]
port 231 nsew signal output
rlabel metal3 s 160792 127848 161592 127968 6 rs1_data[8]
port 232 nsew signal output
rlabel metal2 s 156510 0 156566 800 6 rs1_data[9]
port 233 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 rs2[0]
port 234 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 rs2[1]
port 235 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 rs2[2]
port 236 nsew signal input
rlabel metal3 s 160792 135328 161592 135448 6 rs2[3]
port 237 nsew signal input
rlabel metal2 s 139122 162936 139178 163736 6 rs2[4]
port 238 nsew signal input
rlabel metal3 s 160792 6808 161592 6928 6 rs2_data[0]
port 239 nsew signal output
rlabel metal2 s 132038 162936 132094 163736 6 rs2_data[10]
port 240 nsew signal output
rlabel metal3 s 0 71408 800 71528 6 rs2_data[11]
port 241 nsew signal output
rlabel metal3 s 0 76168 800 76288 6 rs2_data[12]
port 242 nsew signal output
rlabel metal2 s 102414 0 102470 800 6 rs2_data[13]
port 243 nsew signal output
rlabel metal2 s 18 0 74 800 6 rs2_data[14]
port 244 nsew signal output
rlabel metal2 s 121090 0 121146 800 6 rs2_data[15]
port 245 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 rs2_data[16]
port 246 nsew signal output
rlabel metal3 s 0 162528 800 162648 6 rs2_data[17]
port 247 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 rs2_data[18]
port 248 nsew signal output
rlabel metal3 s 0 73448 800 73568 6 rs2_data[19]
port 249 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 rs2_data[1]
port 250 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 rs2_data[20]
port 251 nsew signal output
rlabel metal2 s 94686 162936 94742 163736 6 rs2_data[21]
port 252 nsew signal output
rlabel metal2 s 59910 162936 59966 163736 6 rs2_data[22]
port 253 nsew signal output
rlabel metal2 s 83738 0 83794 800 6 rs2_data[23]
port 254 nsew signal output
rlabel metal2 s 120446 162936 120502 163736 6 rs2_data[24]
port 255 nsew signal output
rlabel metal3 s 160792 38768 161592 38888 6 rs2_data[25]
port 256 nsew signal output
rlabel metal3 s 0 120368 800 120488 6 rs2_data[26]
port 257 nsew signal output
rlabel metal3 s 160792 120368 161592 120488 6 rs2_data[27]
port 258 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 rs2_data[28]
port 259 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 rs2_data[29]
port 260 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 rs2_data[2]
port 261 nsew signal output
rlabel metal3 s 160792 115608 161592 115728 6 rs2_data[30]
port 262 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 rs2_data[31]
port 263 nsew signal output
rlabel metal2 s 110786 162936 110842 163736 6 rs2_data[3]
port 264 nsew signal output
rlabel metal2 s 108854 162936 108910 163736 6 rs2_data[4]
port 265 nsew signal output
rlabel metal3 s 0 157768 800 157888 6 rs2_data[5]
port 266 nsew signal output
rlabel metal2 s 21914 162936 21970 163736 6 rs2_data[6]
port 267 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 rs2_data[7]
port 268 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 rs2_data[8]
port 269 nsew signal output
rlabel metal3 s 0 138048 800 138168 6 rs2_data[9]
port 270 nsew signal output
rlabel metal3 s 160792 78208 161592 78328 6 rst_n
port 271 nsew signal input
rlabel metal4 s 4208 2128 4528 161072 6 vccd1
port 272 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 161072 6 vccd1
port 272 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 161072 6 vccd1
port 272 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 161072 6 vccd1
port 272 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 161072 6 vccd1
port 272 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 161072 6 vccd1
port 272 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 161072 6 vssd1
port 273 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 161072 6 vssd1
port 273 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 161072 6 vssd1
port 273 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 161072 6 vssd1
port 273 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 161072 6 vssd1
port 273 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 161592 163736
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 31813174
string GDS_FILE /home/drewarosa/RISC-V-Single-Cycle-CPU-Core/openlane/ALU/runs/22_09_16_16_48/results/signoff/ALU.magic.gds
string GDS_START 872968
<< end >>

