magic
tech sky130B
magscale 1 2
timestamp 1663701145
<< obsli1 >>
rect 1104 2159 148856 147441
<< obsm1 >>
rect 14 1844 148856 147472
<< metal2 >>
rect 662 149200 718 150000
rect 4526 149200 4582 150000
rect 8390 149200 8446 150000
rect 12898 149200 12954 150000
rect 16762 149200 16818 150000
rect 20626 149200 20682 150000
rect 25134 149200 25190 150000
rect 28998 149200 29054 150000
rect 33506 149200 33562 150000
rect 37370 149200 37426 150000
rect 41234 149200 41290 150000
rect 45742 149200 45798 150000
rect 49606 149200 49662 150000
rect 53470 149200 53526 150000
rect 57978 149200 58034 150000
rect 61842 149200 61898 150000
rect 65706 149200 65762 150000
rect 70214 149200 70270 150000
rect 74078 149200 74134 150000
rect 77942 149200 77998 150000
rect 82450 149200 82506 150000
rect 86314 149200 86370 150000
rect 90178 149200 90234 150000
rect 94686 149200 94742 150000
rect 98550 149200 98606 150000
rect 102414 149200 102470 150000
rect 106922 149200 106978 150000
rect 110786 149200 110842 150000
rect 115294 149200 115350 150000
rect 119158 149200 119214 150000
rect 123022 149200 123078 150000
rect 127530 149200 127586 150000
rect 131394 149200 131450 150000
rect 135258 149200 135314 150000
rect 139766 149200 139822 150000
rect 143630 149200 143686 150000
rect 147494 149200 147550 150000
rect 18 0 74 800
rect 3882 0 3938 800
rect 7746 0 7802 800
rect 12254 0 12310 800
rect 16118 0 16174 800
rect 19982 0 20038 800
rect 24490 0 24546 800
rect 28354 0 28410 800
rect 32218 0 32274 800
rect 36726 0 36782 800
rect 40590 0 40646 800
rect 44454 0 44510 800
rect 48962 0 49018 800
rect 52826 0 52882 800
rect 56690 0 56746 800
rect 61198 0 61254 800
rect 65062 0 65118 800
rect 68926 0 68982 800
rect 73434 0 73490 800
rect 77298 0 77354 800
rect 81162 0 81218 800
rect 85670 0 85726 800
rect 89534 0 89590 800
rect 94042 0 94098 800
rect 97906 0 97962 800
rect 101770 0 101826 800
rect 106278 0 106334 800
rect 110142 0 110198 800
rect 114006 0 114062 800
rect 118514 0 118570 800
rect 122378 0 122434 800
rect 126242 0 126298 800
rect 130750 0 130806 800
rect 134614 0 134670 800
rect 138478 0 138534 800
rect 142986 0 143042 800
rect 146850 0 146906 800
<< obsm2 >>
rect 20 149144 606 149200
rect 774 149144 4470 149200
rect 4638 149144 8334 149200
rect 8502 149144 12842 149200
rect 13010 149144 16706 149200
rect 16874 149144 20570 149200
rect 20738 149144 25078 149200
rect 25246 149144 28942 149200
rect 29110 149144 33450 149200
rect 33618 149144 37314 149200
rect 37482 149144 41178 149200
rect 41346 149144 45686 149200
rect 45854 149144 49550 149200
rect 49718 149144 53414 149200
rect 53582 149144 57922 149200
rect 58090 149144 61786 149200
rect 61954 149144 65650 149200
rect 65818 149144 70158 149200
rect 70326 149144 74022 149200
rect 74190 149144 77886 149200
rect 78054 149144 82394 149200
rect 82562 149144 86258 149200
rect 86426 149144 90122 149200
rect 90290 149144 94630 149200
rect 94798 149144 98494 149200
rect 98662 149144 102358 149200
rect 102526 149144 106866 149200
rect 107034 149144 110730 149200
rect 110898 149144 115238 149200
rect 115406 149144 119102 149200
rect 119270 149144 122966 149200
rect 123134 149144 127474 149200
rect 127642 149144 131338 149200
rect 131506 149144 135202 149200
rect 135370 149144 139710 149200
rect 139878 149144 143574 149200
rect 143742 149144 147438 149200
rect 147606 149144 148194 149200
rect 20 856 148194 149144
rect 130 734 3826 856
rect 3994 734 7690 856
rect 7858 734 12198 856
rect 12366 734 16062 856
rect 16230 734 19926 856
rect 20094 734 24434 856
rect 24602 734 28298 856
rect 28466 734 32162 856
rect 32330 734 36670 856
rect 36838 734 40534 856
rect 40702 734 44398 856
rect 44566 734 48906 856
rect 49074 734 52770 856
rect 52938 734 56634 856
rect 56802 734 61142 856
rect 61310 734 65006 856
rect 65174 734 68870 856
rect 69038 734 73378 856
rect 73546 734 77242 856
rect 77410 734 81106 856
rect 81274 734 85614 856
rect 85782 734 89478 856
rect 89646 734 93986 856
rect 94154 734 97850 856
rect 98018 734 101714 856
rect 101882 734 106222 856
rect 106390 734 110086 856
rect 110254 734 113950 856
rect 114118 734 118458 856
rect 118626 734 122322 856
rect 122490 734 126186 856
rect 126354 734 130694 856
rect 130862 734 134558 856
rect 134726 734 138422 856
rect 138590 734 142930 856
rect 143098 734 146794 856
rect 146962 734 148194 856
<< metal3 >>
rect 149200 147568 150000 147688
rect 0 146208 800 146328
rect 149200 143488 150000 143608
rect 0 142128 800 142248
rect 149200 139408 150000 139528
rect 0 138048 800 138168
rect 149200 134648 150000 134768
rect 0 133288 800 133408
rect 149200 130568 150000 130688
rect 0 129208 800 129328
rect 149200 126488 150000 126608
rect 0 125128 800 125248
rect 149200 121728 150000 121848
rect 0 120368 800 120488
rect 149200 117648 150000 117768
rect 0 116288 800 116408
rect 149200 113568 150000 113688
rect 0 112208 800 112328
rect 149200 108808 150000 108928
rect 0 107448 800 107568
rect 149200 104728 150000 104848
rect 0 103368 800 103488
rect 149200 99968 150000 100088
rect 0 99288 800 99408
rect 149200 95888 150000 96008
rect 0 94528 800 94648
rect 149200 91808 150000 91928
rect 0 90448 800 90568
rect 149200 87048 150000 87168
rect 0 85688 800 85808
rect 149200 82968 150000 83088
rect 0 81608 800 81728
rect 149200 78888 150000 79008
rect 0 77528 800 77648
rect 149200 74128 150000 74248
rect 0 72768 800 72888
rect 149200 70048 150000 70168
rect 0 68688 800 68808
rect 149200 65968 150000 66088
rect 0 64608 800 64728
rect 149200 61208 150000 61328
rect 0 59848 800 59968
rect 149200 57128 150000 57248
rect 0 55768 800 55888
rect 149200 53048 150000 53168
rect 0 51688 800 51808
rect 149200 48288 150000 48408
rect 0 46928 800 47048
rect 149200 44208 150000 44328
rect 0 42848 800 42968
rect 149200 40128 150000 40248
rect 0 38768 800 38888
rect 149200 35368 150000 35488
rect 0 34008 800 34128
rect 149200 31288 150000 31408
rect 0 29928 800 30048
rect 149200 27208 150000 27328
rect 0 25848 800 25968
rect 149200 22448 150000 22568
rect 0 21088 800 21208
rect 149200 18368 150000 18488
rect 0 17008 800 17128
rect 149200 13608 150000 13728
rect 0 12928 800 13048
rect 149200 9528 150000 9648
rect 0 8168 800 8288
rect 149200 5448 150000 5568
rect 0 4088 800 4208
rect 149200 688 150000 808
<< obsm3 >>
rect 749 146408 149200 147457
rect 880 146128 149200 146408
rect 749 143688 149200 146128
rect 749 143408 149120 143688
rect 749 142328 149200 143408
rect 880 142048 149200 142328
rect 749 139608 149200 142048
rect 749 139328 149120 139608
rect 749 138248 149200 139328
rect 880 137968 149200 138248
rect 749 134848 149200 137968
rect 749 134568 149120 134848
rect 749 133488 149200 134568
rect 880 133208 149200 133488
rect 749 130768 149200 133208
rect 749 130488 149120 130768
rect 749 129408 149200 130488
rect 880 129128 149200 129408
rect 749 126688 149200 129128
rect 749 126408 149120 126688
rect 749 125328 149200 126408
rect 880 125048 149200 125328
rect 749 121928 149200 125048
rect 749 121648 149120 121928
rect 749 120568 149200 121648
rect 880 120288 149200 120568
rect 749 117848 149200 120288
rect 749 117568 149120 117848
rect 749 116488 149200 117568
rect 880 116208 149200 116488
rect 749 113768 149200 116208
rect 749 113488 149120 113768
rect 749 112408 149200 113488
rect 880 112128 149200 112408
rect 749 109008 149200 112128
rect 749 108728 149120 109008
rect 749 107648 149200 108728
rect 880 107368 149200 107648
rect 749 104928 149200 107368
rect 749 104648 149120 104928
rect 749 103568 149200 104648
rect 880 103288 149200 103568
rect 749 100168 149200 103288
rect 749 99888 149120 100168
rect 749 99488 149200 99888
rect 880 99208 149200 99488
rect 749 96088 149200 99208
rect 749 95808 149120 96088
rect 749 94728 149200 95808
rect 880 94448 149200 94728
rect 749 92008 149200 94448
rect 749 91728 149120 92008
rect 749 90648 149200 91728
rect 880 90368 149200 90648
rect 749 87248 149200 90368
rect 749 86968 149120 87248
rect 749 85888 149200 86968
rect 880 85608 149200 85888
rect 749 83168 149200 85608
rect 749 82888 149120 83168
rect 749 81808 149200 82888
rect 880 81528 149200 81808
rect 749 79088 149200 81528
rect 749 78808 149120 79088
rect 749 77728 149200 78808
rect 880 77448 149200 77728
rect 749 74328 149200 77448
rect 749 74048 149120 74328
rect 749 72968 149200 74048
rect 880 72688 149200 72968
rect 749 70248 149200 72688
rect 749 69968 149120 70248
rect 749 68888 149200 69968
rect 880 68608 149200 68888
rect 749 66168 149200 68608
rect 749 65888 149120 66168
rect 749 64808 149200 65888
rect 880 64528 149200 64808
rect 749 61408 149200 64528
rect 749 61128 149120 61408
rect 749 60048 149200 61128
rect 880 59768 149200 60048
rect 749 57328 149200 59768
rect 749 57048 149120 57328
rect 749 55968 149200 57048
rect 880 55688 149200 55968
rect 749 53248 149200 55688
rect 749 52968 149120 53248
rect 749 51888 149200 52968
rect 880 51608 149200 51888
rect 749 48488 149200 51608
rect 749 48208 149120 48488
rect 749 47128 149200 48208
rect 880 46848 149200 47128
rect 749 44408 149200 46848
rect 749 44128 149120 44408
rect 749 43048 149200 44128
rect 880 42768 149200 43048
rect 749 40328 149200 42768
rect 749 40048 149120 40328
rect 749 38968 149200 40048
rect 880 38688 149200 38968
rect 749 35568 149200 38688
rect 749 35288 149120 35568
rect 749 34208 149200 35288
rect 880 33928 149200 34208
rect 749 31488 149200 33928
rect 749 31208 149120 31488
rect 749 30128 149200 31208
rect 880 29848 149200 30128
rect 749 27408 149200 29848
rect 749 27128 149120 27408
rect 749 26048 149200 27128
rect 880 25768 149200 26048
rect 749 22648 149200 25768
rect 749 22368 149120 22648
rect 749 21288 149200 22368
rect 880 21008 149200 21288
rect 749 18568 149200 21008
rect 749 18288 149120 18568
rect 749 17208 149200 18288
rect 880 16928 149200 17208
rect 749 13808 149200 16928
rect 749 13528 149120 13808
rect 749 13128 149200 13528
rect 880 12848 149200 13128
rect 749 9728 149200 12848
rect 749 9448 149120 9728
rect 749 8368 149200 9448
rect 880 8088 149200 8368
rect 749 5648 149200 8088
rect 749 5368 149120 5648
rect 749 4288 149200 5368
rect 880 4008 149200 4288
rect 749 1939 149200 4008
<< metal4 >>
rect 4208 2128 4528 147472
rect 19568 2128 19888 147472
rect 34928 2128 35248 147472
rect 50288 2128 50608 147472
rect 65648 2128 65968 147472
rect 81008 2128 81328 147472
rect 96368 2128 96688 147472
rect 111728 2128 112048 147472
rect 127088 2128 127408 147472
rect 142448 2128 142768 147472
<< obsm4 >>
rect 2451 2048 4128 146981
rect 4608 2048 19488 146981
rect 19968 2048 34848 146981
rect 35328 2048 50208 146981
rect 50688 2048 65568 146981
rect 66048 2048 71885 146981
rect 2451 1939 71885 2048
<< labels >>
rlabel metal2 s 44454 0 44510 800 6 clk
port 1 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 funct3[0]
port 2 nsew signal input
rlabel metal3 s 149200 44208 150000 44328 6 funct3[1]
port 3 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 funct3[2]
port 4 nsew signal input
rlabel metal2 s 135258 149200 135314 150000 6 la_dram_select[0]
port 5 nsew signal input
rlabel metal2 s 139766 149200 139822 150000 6 la_dram_select[1]
port 6 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 la_dram_select[2]
port 7 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 la_dram_select[3]
port 8 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 la_read_data[0]
port 9 nsew signal output
rlabel metal2 s 130750 0 130806 800 6 la_read_data[10]
port 10 nsew signal output
rlabel metal3 s 149200 126488 150000 126608 6 la_read_data[11]
port 11 nsew signal output
rlabel metal2 s 98550 149200 98606 150000 6 la_read_data[12]
port 12 nsew signal output
rlabel metal3 s 149200 108808 150000 108928 6 la_read_data[13]
port 13 nsew signal output
rlabel metal2 s 45742 149200 45798 150000 6 la_read_data[14]
port 14 nsew signal output
rlabel metal3 s 0 107448 800 107568 6 la_read_data[15]
port 15 nsew signal output
rlabel metal2 s 74078 149200 74134 150000 6 la_read_data[16]
port 16 nsew signal output
rlabel metal3 s 149200 134648 150000 134768 6 la_read_data[17]
port 17 nsew signal output
rlabel metal2 s 77298 0 77354 800 6 la_read_data[18]
port 18 nsew signal output
rlabel metal3 s 149200 104728 150000 104848 6 la_read_data[19]
port 19 nsew signal output
rlabel metal2 s 94686 149200 94742 150000 6 la_read_data[1]
port 20 nsew signal output
rlabel metal3 s 149200 117648 150000 117768 6 la_read_data[20]
port 21 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 la_read_data[21]
port 22 nsew signal output
rlabel metal2 s 8390 149200 8446 150000 6 la_read_data[22]
port 23 nsew signal output
rlabel metal2 s 77942 149200 77998 150000 6 la_read_data[23]
port 24 nsew signal output
rlabel metal3 s 149200 31288 150000 31408 6 la_read_data[24]
port 25 nsew signal output
rlabel metal3 s 0 68688 800 68808 6 la_read_data[25]
port 26 nsew signal output
rlabel metal2 s 25134 149200 25190 150000 6 la_read_data[26]
port 27 nsew signal output
rlabel metal2 s 20626 149200 20682 150000 6 la_read_data[27]
port 28 nsew signal output
rlabel metal2 s 123022 149200 123078 150000 6 la_read_data[28]
port 29 nsew signal output
rlabel metal2 s 70214 149200 70270 150000 6 la_read_data[29]
port 30 nsew signal output
rlabel metal3 s 149200 91808 150000 91928 6 la_read_data[2]
port 31 nsew signal output
rlabel metal2 s 662 149200 718 150000 6 la_read_data[30]
port 32 nsew signal output
rlabel metal3 s 149200 99968 150000 100088 6 la_read_data[31]
port 33 nsew signal output
rlabel metal3 s 0 116288 800 116408 6 la_read_data[3]
port 34 nsew signal output
rlabel metal3 s 0 133288 800 133408 6 la_read_data[4]
port 35 nsew signal output
rlabel metal3 s 149200 5448 150000 5568 6 la_read_data[5]
port 36 nsew signal output
rlabel metal3 s 0 99288 800 99408 6 la_read_data[6]
port 37 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 la_read_data[7]
port 38 nsew signal output
rlabel metal2 s 119158 149200 119214 150000 6 la_read_data[8]
port 39 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 la_read_data[9]
port 40 nsew signal output
rlabel metal2 s 126242 0 126298 800 6 mem_write
port 41 nsew signal input
rlabel metal3 s 149200 65968 150000 66088 6 memory_address[0]
port 42 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 memory_address[10]
port 43 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 memory_address[11]
port 44 nsew signal input
rlabel metal2 s 61842 149200 61898 150000 6 memory_address[12]
port 45 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 memory_address[13]
port 46 nsew signal input
rlabel metal3 s 149200 48288 150000 48408 6 memory_address[14]
port 47 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 memory_address[15]
port 48 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 memory_address[16]
port 49 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 memory_address[17]
port 50 nsew signal input
rlabel metal3 s 149200 121728 150000 121848 6 memory_address[18]
port 51 nsew signal input
rlabel metal3 s 149200 9528 150000 9648 6 memory_address[19]
port 52 nsew signal input
rlabel metal2 s 49606 149200 49662 150000 6 memory_address[1]
port 53 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 memory_address[20]
port 54 nsew signal input
rlabel metal2 s 33506 149200 33562 150000 6 memory_address[21]
port 55 nsew signal input
rlabel metal3 s 149200 143488 150000 143608 6 memory_address[22]
port 56 nsew signal input
rlabel metal2 s 86314 149200 86370 150000 6 memory_address[23]
port 57 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 memory_address[24]
port 58 nsew signal input
rlabel metal2 s 12898 149200 12954 150000 6 memory_address[25]
port 59 nsew signal input
rlabel metal3 s 149200 53048 150000 53168 6 memory_address[26]
port 60 nsew signal input
rlabel metal2 s 16762 149200 16818 150000 6 memory_address[27]
port 61 nsew signal input
rlabel metal3 s 149200 688 150000 808 6 memory_address[28]
port 62 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 memory_address[29]
port 63 nsew signal input
rlabel metal2 s 57978 149200 58034 150000 6 memory_address[2]
port 64 nsew signal input
rlabel metal2 s 41234 149200 41290 150000 6 memory_address[30]
port 65 nsew signal input
rlabel metal3 s 0 146208 800 146328 6 memory_address[31]
port 66 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 memory_address[3]
port 67 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 memory_address[4]
port 68 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 memory_address[5]
port 69 nsew signal input
rlabel metal2 s 127530 149200 127586 150000 6 memory_address[6]
port 70 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 memory_address[7]
port 71 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 memory_address[8]
port 72 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 memory_address[9]
port 73 nsew signal input
rlabel metal3 s 149200 18368 150000 18488 6 rd[0]
port 74 nsew signal input
rlabel metal2 s 102414 149200 102470 150000 6 rd[1]
port 75 nsew signal input
rlabel metal3 s 149200 147568 150000 147688 6 rd[2]
port 76 nsew signal input
rlabel metal2 s 65706 149200 65762 150000 6 rd[3]
port 77 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 rd[4]
port 78 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 read_data[0]
port 79 nsew signal output
rlabel metal2 s 146850 0 146906 800 6 read_data[10]
port 80 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 read_data[11]
port 81 nsew signal output
rlabel metal3 s 149200 78888 150000 79008 6 read_data[12]
port 82 nsew signal output
rlabel metal3 s 149200 57128 150000 57248 6 read_data[13]
port 83 nsew signal output
rlabel metal2 s 147494 149200 147550 150000 6 read_data[14]
port 84 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 read_data[15]
port 85 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 read_data[16]
port 86 nsew signal output
rlabel metal3 s 149200 61208 150000 61328 6 read_data[17]
port 87 nsew signal output
rlabel metal3 s 0 103368 800 103488 6 read_data[18]
port 88 nsew signal output
rlabel metal3 s 149200 35368 150000 35488 6 read_data[19]
port 89 nsew signal output
rlabel metal2 s 138478 0 138534 800 6 read_data[1]
port 90 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 read_data[20]
port 91 nsew signal output
rlabel metal3 s 149200 82968 150000 83088 6 read_data[21]
port 92 nsew signal output
rlabel metal2 s 143630 149200 143686 150000 6 read_data[22]
port 93 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 read_data[23]
port 94 nsew signal output
rlabel metal3 s 149200 27208 150000 27328 6 read_data[24]
port 95 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 read_data[25]
port 96 nsew signal output
rlabel metal2 s 142986 0 143042 800 6 read_data[26]
port 97 nsew signal output
rlabel metal2 s 53470 149200 53526 150000 6 read_data[27]
port 98 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 read_data[28]
port 99 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 read_data[29]
port 100 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 read_data[2]
port 101 nsew signal output
rlabel metal3 s 149200 13608 150000 13728 6 read_data[30]
port 102 nsew signal output
rlabel metal3 s 149200 113568 150000 113688 6 read_data[31]
port 103 nsew signal output
rlabel metal3 s 149200 74128 150000 74248 6 read_data[3]
port 104 nsew signal output
rlabel metal2 s 122378 0 122434 800 6 read_data[4]
port 105 nsew signal output
rlabel metal3 s 0 90448 800 90568 6 read_data[5]
port 106 nsew signal output
rlabel metal3 s 149200 40128 150000 40248 6 read_data[6]
port 107 nsew signal output
rlabel metal3 s 0 120368 800 120488 6 read_data[7]
port 108 nsew signal output
rlabel metal3 s 149200 87048 150000 87168 6 read_data[8]
port 109 nsew signal output
rlabel metal3 s 149200 130568 150000 130688 6 read_data[9]
port 110 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 rst_n
port 111 nsew signal input
rlabel metal4 s 4208 2128 4528 147472 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 147472 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 147472 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 147472 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 147472 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 147472 6 vssd1
port 113 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 147472 6 vssd1
port 113 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 147472 6 vssd1
port 113 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 147472 6 vssd1
port 113 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 147472 6 vssd1
port 113 nsew ground bidirectional
rlabel metal3 s 149200 139408 150000 139528 6 write_data[0]
port 114 nsew signal input
rlabel metal3 s 0 125128 800 125248 6 write_data[10]
port 115 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 write_data[11]
port 116 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 write_data[12]
port 117 nsew signal input
rlabel metal2 s 18 0 74 800 6 write_data[13]
port 118 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 write_data[14]
port 119 nsew signal input
rlabel metal3 s 0 142128 800 142248 6 write_data[15]
port 120 nsew signal input
rlabel metal2 s 37370 149200 37426 150000 6 write_data[16]
port 121 nsew signal input
rlabel metal2 s 90178 149200 90234 150000 6 write_data[17]
port 122 nsew signal input
rlabel metal3 s 0 112208 800 112328 6 write_data[18]
port 123 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 write_data[19]
port 124 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 write_data[1]
port 125 nsew signal input
rlabel metal2 s 115294 149200 115350 150000 6 write_data[20]
port 126 nsew signal input
rlabel metal2 s 82450 149200 82506 150000 6 write_data[21]
port 127 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 write_data[22]
port 128 nsew signal input
rlabel metal2 s 131394 149200 131450 150000 6 write_data[23]
port 129 nsew signal input
rlabel metal3 s 149200 22448 150000 22568 6 write_data[24]
port 130 nsew signal input
rlabel metal3 s 0 138048 800 138168 6 write_data[25]
port 131 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 write_data[26]
port 132 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 write_data[27]
port 133 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 write_data[28]
port 134 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 write_data[29]
port 135 nsew signal input
rlabel metal3 s 149200 95888 150000 96008 6 write_data[2]
port 136 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 write_data[30]
port 137 nsew signal input
rlabel metal2 s 110786 149200 110842 150000 6 write_data[31]
port 138 nsew signal input
rlabel metal2 s 106922 149200 106978 150000 6 write_data[3]
port 139 nsew signal input
rlabel metal2 s 4526 149200 4582 150000 6 write_data[4]
port 140 nsew signal input
rlabel metal2 s 28998 149200 29054 150000 6 write_data[5]
port 141 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 write_data[6]
port 142 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 write_data[7]
port 143 nsew signal input
rlabel metal3 s 0 129208 800 129328 6 write_data[8]
port 144 nsew signal input
rlabel metal3 s 149200 70048 150000 70168 6 write_data[9]
port 145 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 150000 150000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 18354662
string GDS_FILE /home/drewarosa/RISC-V-Single-Cycle-CPU-Core/openlane/DMemory/runs/22_09_20_15_07/results/signoff/DMemory.magic.gds
string GDS_START 500430
<< end >>

