magic
tech sky130B
magscale 1 2
timestamp 1663703974
<< obsli1 >>
rect 1104 2159 248860 247537
<< obsm1 >>
rect 14 8 248860 247852
<< metal2 >>
rect 18 249200 74 250000
rect 3882 249200 3938 250000
rect 7102 249200 7158 250000
rect 10966 249200 11022 250000
rect 14830 249200 14886 250000
rect 18050 249200 18106 250000
rect 21914 249200 21970 250000
rect 25134 249200 25190 250000
rect 28998 249200 29054 250000
rect 32862 249200 32918 250000
rect 36082 249200 36138 250000
rect 39946 249200 40002 250000
rect 43166 249200 43222 250000
rect 47030 249200 47086 250000
rect 50250 249200 50306 250000
rect 54114 249200 54170 250000
rect 57978 249200 58034 250000
rect 61198 249200 61254 250000
rect 65062 249200 65118 250000
rect 68282 249200 68338 250000
rect 72146 249200 72202 250000
rect 76010 249200 76066 250000
rect 79230 249200 79286 250000
rect 83094 249200 83150 250000
rect 86314 249200 86370 250000
rect 90178 249200 90234 250000
rect 93398 249200 93454 250000
rect 97262 249200 97318 250000
rect 101126 249200 101182 250000
rect 104346 249200 104402 250000
rect 108210 249200 108266 250000
rect 111430 249200 111486 250000
rect 115294 249200 115350 250000
rect 119158 249200 119214 250000
rect 122378 249200 122434 250000
rect 126242 249200 126298 250000
rect 129462 249200 129518 250000
rect 133326 249200 133382 250000
rect 137190 249200 137246 250000
rect 140410 249200 140466 250000
rect 144274 249200 144330 250000
rect 147494 249200 147550 250000
rect 151358 249200 151414 250000
rect 154578 249200 154634 250000
rect 158442 249200 158498 250000
rect 162306 249200 162362 250000
rect 165526 249200 165582 250000
rect 169390 249200 169446 250000
rect 172610 249200 172666 250000
rect 176474 249200 176530 250000
rect 180338 249200 180394 250000
rect 183558 249200 183614 250000
rect 187422 249200 187478 250000
rect 190642 249200 190698 250000
rect 194506 249200 194562 250000
rect 197726 249200 197782 250000
rect 201590 249200 201646 250000
rect 205454 249200 205510 250000
rect 208674 249200 208730 250000
rect 212538 249200 212594 250000
rect 215758 249200 215814 250000
rect 219622 249200 219678 250000
rect 223486 249200 223542 250000
rect 226706 249200 226762 250000
rect 230570 249200 230626 250000
rect 233790 249200 233846 250000
rect 237654 249200 237710 250000
rect 241518 249200 241574 250000
rect 244738 249200 244794 250000
rect 248602 249200 248658 250000
rect 18 0 74 800
rect 3238 0 3294 800
rect 7102 0 7158 800
rect 10322 0 10378 800
rect 14186 0 14242 800
rect 17406 0 17462 800
rect 21270 0 21326 800
rect 25134 0 25190 800
rect 28354 0 28410 800
rect 32218 0 32274 800
rect 35438 0 35494 800
rect 39302 0 39358 800
rect 43166 0 43222 800
rect 46386 0 46442 800
rect 50250 0 50306 800
rect 53470 0 53526 800
rect 57334 0 57390 800
rect 60554 0 60610 800
rect 64418 0 64474 800
rect 68282 0 68338 800
rect 71502 0 71558 800
rect 75366 0 75422 800
rect 78586 0 78642 800
rect 82450 0 82506 800
rect 86314 0 86370 800
rect 89534 0 89590 800
rect 93398 0 93454 800
rect 96618 0 96674 800
rect 100482 0 100538 800
rect 104346 0 104402 800
rect 107566 0 107622 800
rect 111430 0 111486 800
rect 114650 0 114706 800
rect 118514 0 118570 800
rect 121734 0 121790 800
rect 125598 0 125654 800
rect 129462 0 129518 800
rect 132682 0 132738 800
rect 136546 0 136602 800
rect 139766 0 139822 800
rect 143630 0 143686 800
rect 147494 0 147550 800
rect 150714 0 150770 800
rect 154578 0 154634 800
rect 157798 0 157854 800
rect 161662 0 161718 800
rect 164882 0 164938 800
rect 168746 0 168802 800
rect 172610 0 172666 800
rect 175830 0 175886 800
rect 179694 0 179750 800
rect 182914 0 182970 800
rect 186778 0 186834 800
rect 190642 0 190698 800
rect 193862 0 193918 800
rect 197726 0 197782 800
rect 200946 0 201002 800
rect 204810 0 204866 800
rect 208674 0 208730 800
rect 211894 0 211950 800
rect 215758 0 215814 800
rect 218978 0 219034 800
rect 222842 0 222898 800
rect 226062 0 226118 800
rect 229926 0 229982 800
rect 233790 0 233846 800
rect 237010 0 237066 800
rect 240874 0 240930 800
rect 244094 0 244150 800
rect 247958 0 248014 800
<< obsm2 >>
rect 130 249144 3826 249234
rect 3994 249144 7046 249234
rect 7214 249144 10910 249234
rect 11078 249144 14774 249234
rect 14942 249144 17994 249234
rect 18162 249144 21858 249234
rect 22026 249144 25078 249234
rect 25246 249144 28942 249234
rect 29110 249144 32806 249234
rect 32974 249144 36026 249234
rect 36194 249144 39890 249234
rect 40058 249144 43110 249234
rect 43278 249144 46974 249234
rect 47142 249144 50194 249234
rect 50362 249144 54058 249234
rect 54226 249144 57922 249234
rect 58090 249144 61142 249234
rect 61310 249144 65006 249234
rect 65174 249144 68226 249234
rect 68394 249144 72090 249234
rect 72258 249144 75954 249234
rect 76122 249144 79174 249234
rect 79342 249144 83038 249234
rect 83206 249144 86258 249234
rect 86426 249144 90122 249234
rect 90290 249144 93342 249234
rect 93510 249144 97206 249234
rect 97374 249144 101070 249234
rect 101238 249144 104290 249234
rect 104458 249144 108154 249234
rect 108322 249144 111374 249234
rect 111542 249144 115238 249234
rect 115406 249144 119102 249234
rect 119270 249144 122322 249234
rect 122490 249144 126186 249234
rect 126354 249144 129406 249234
rect 129574 249144 133270 249234
rect 133438 249144 137134 249234
rect 137302 249144 140354 249234
rect 140522 249144 144218 249234
rect 144386 249144 147438 249234
rect 147606 249144 151302 249234
rect 151470 249144 154522 249234
rect 154690 249144 158386 249234
rect 158554 249144 162250 249234
rect 162418 249144 165470 249234
rect 165638 249144 169334 249234
rect 169502 249144 172554 249234
rect 172722 249144 176418 249234
rect 176586 249144 180282 249234
rect 180450 249144 183502 249234
rect 183670 249144 187366 249234
rect 187534 249144 190586 249234
rect 190754 249144 194450 249234
rect 194618 249144 197670 249234
rect 197838 249144 201534 249234
rect 201702 249144 205398 249234
rect 205566 249144 208618 249234
rect 208786 249144 212482 249234
rect 212650 249144 215702 249234
rect 215870 249144 219566 249234
rect 219734 249144 223430 249234
rect 223598 249144 226650 249234
rect 226818 249144 230514 249234
rect 230682 249144 233734 249234
rect 233902 249144 237598 249234
rect 237766 249144 241462 249234
rect 241630 249144 244682 249234
rect 244850 249144 248546 249234
rect 20 856 248656 249144
rect 130 2 3182 856
rect 3350 2 7046 856
rect 7214 2 10266 856
rect 10434 2 14130 856
rect 14298 2 17350 856
rect 17518 2 21214 856
rect 21382 2 25078 856
rect 25246 2 28298 856
rect 28466 2 32162 856
rect 32330 2 35382 856
rect 35550 2 39246 856
rect 39414 2 43110 856
rect 43278 2 46330 856
rect 46498 2 50194 856
rect 50362 2 53414 856
rect 53582 2 57278 856
rect 57446 2 60498 856
rect 60666 2 64362 856
rect 64530 2 68226 856
rect 68394 2 71446 856
rect 71614 2 75310 856
rect 75478 2 78530 856
rect 78698 2 82394 856
rect 82562 2 86258 856
rect 86426 2 89478 856
rect 89646 2 93342 856
rect 93510 2 96562 856
rect 96730 2 100426 856
rect 100594 2 104290 856
rect 104458 2 107510 856
rect 107678 2 111374 856
rect 111542 2 114594 856
rect 114762 2 118458 856
rect 118626 2 121678 856
rect 121846 2 125542 856
rect 125710 2 129406 856
rect 129574 2 132626 856
rect 132794 2 136490 856
rect 136658 2 139710 856
rect 139878 2 143574 856
rect 143742 2 147438 856
rect 147606 2 150658 856
rect 150826 2 154522 856
rect 154690 2 157742 856
rect 157910 2 161606 856
rect 161774 2 164826 856
rect 164994 2 168690 856
rect 168858 2 172554 856
rect 172722 2 175774 856
rect 175942 2 179638 856
rect 179806 2 182858 856
rect 183026 2 186722 856
rect 186890 2 190586 856
rect 190754 2 193806 856
rect 193974 2 197670 856
rect 197838 2 200890 856
rect 201058 2 204754 856
rect 204922 2 208618 856
rect 208786 2 211838 856
rect 212006 2 215702 856
rect 215870 2 218922 856
rect 219090 2 222786 856
rect 222954 2 226006 856
rect 226174 2 229870 856
rect 230038 2 233734 856
rect 233902 2 236954 856
rect 237122 2 240818 856
rect 240986 2 244038 856
rect 244206 2 247902 856
rect 248070 2 248656 856
<< metal3 >>
rect 249200 248208 250000 248328
rect 0 246848 800 246968
rect 249200 244128 250000 244248
rect 0 242768 800 242888
rect 249200 240728 250000 240848
rect 0 238688 800 238808
rect 249200 236648 250000 236768
rect 0 235288 800 235408
rect 249200 232568 250000 232688
rect 0 231208 800 231328
rect 249200 229168 250000 229288
rect 0 227808 800 227928
rect 249200 225088 250000 225208
rect 0 223728 800 223848
rect 249200 221688 250000 221808
rect 0 220328 800 220448
rect 249200 217608 250000 217728
rect 0 216248 800 216368
rect 249200 213528 250000 213648
rect 0 212168 800 212288
rect 249200 210128 250000 210248
rect 0 208768 800 208888
rect 249200 206048 250000 206168
rect 0 204688 800 204808
rect 249200 202648 250000 202768
rect 0 201288 800 201408
rect 249200 198568 250000 198688
rect 0 197208 800 197328
rect 249200 194488 250000 194608
rect 0 193128 800 193248
rect 249200 191088 250000 191208
rect 0 189728 800 189848
rect 249200 187008 250000 187128
rect 0 185648 800 185768
rect 249200 183608 250000 183728
rect 0 182248 800 182368
rect 249200 179528 250000 179648
rect 0 178168 800 178288
rect 249200 176128 250000 176248
rect 0 174088 800 174208
rect 249200 172048 250000 172168
rect 0 170688 800 170808
rect 249200 167968 250000 168088
rect 0 166608 800 166728
rect 249200 164568 250000 164688
rect 0 163208 800 163328
rect 249200 160488 250000 160608
rect 0 159128 800 159248
rect 249200 157088 250000 157208
rect 0 155728 800 155848
rect 249200 153008 250000 153128
rect 0 151648 800 151768
rect 249200 148928 250000 149048
rect 0 147568 800 147688
rect 249200 145528 250000 145648
rect 0 144168 800 144288
rect 249200 141448 250000 141568
rect 0 140088 800 140208
rect 249200 138048 250000 138168
rect 0 136688 800 136808
rect 249200 133968 250000 134088
rect 0 132608 800 132728
rect 249200 130568 250000 130688
rect 0 128528 800 128648
rect 249200 126488 250000 126608
rect 0 125128 800 125248
rect 249200 122408 250000 122528
rect 0 121048 800 121168
rect 249200 119008 250000 119128
rect 0 117648 800 117768
rect 249200 114928 250000 115048
rect 0 113568 800 113688
rect 249200 111528 250000 111648
rect 0 110168 800 110288
rect 249200 107448 250000 107568
rect 0 106088 800 106208
rect 249200 103368 250000 103488
rect 0 102008 800 102128
rect 249200 99968 250000 100088
rect 0 98608 800 98728
rect 249200 95888 250000 96008
rect 0 94528 800 94648
rect 249200 92488 250000 92608
rect 0 91128 800 91248
rect 249200 88408 250000 88528
rect 0 87048 800 87168
rect 249200 84328 250000 84448
rect 0 82968 800 83088
rect 249200 80928 250000 81048
rect 0 79568 800 79688
rect 249200 76848 250000 76968
rect 0 75488 800 75608
rect 249200 73448 250000 73568
rect 0 72088 800 72208
rect 249200 69368 250000 69488
rect 0 68008 800 68128
rect 249200 65968 250000 66088
rect 0 63928 800 64048
rect 249200 61888 250000 62008
rect 0 60528 800 60648
rect 249200 57808 250000 57928
rect 0 56448 800 56568
rect 249200 54408 250000 54528
rect 0 53048 800 53168
rect 249200 50328 250000 50448
rect 0 48968 800 49088
rect 249200 46928 250000 47048
rect 0 45568 800 45688
rect 249200 42848 250000 42968
rect 0 41488 800 41608
rect 249200 38768 250000 38888
rect 0 37408 800 37528
rect 249200 35368 250000 35488
rect 0 34008 800 34128
rect 249200 31288 250000 31408
rect 0 29928 800 30048
rect 249200 27888 250000 28008
rect 0 26528 800 26648
rect 249200 23808 250000 23928
rect 0 22448 800 22568
rect 249200 20408 250000 20528
rect 0 18368 800 18488
rect 249200 16328 250000 16448
rect 0 14968 800 15088
rect 249200 12248 250000 12368
rect 0 10888 800 11008
rect 249200 8848 250000 8968
rect 0 7488 800 7608
rect 249200 4768 250000 4888
rect 0 3408 800 3528
rect 249200 1368 250000 1488
<< obsm3 >>
rect 800 248128 249120 248301
rect 800 247048 249200 248128
rect 880 246768 249200 247048
rect 800 244328 249200 246768
rect 800 244048 249120 244328
rect 800 242968 249200 244048
rect 880 242688 249200 242968
rect 800 240928 249200 242688
rect 800 240648 249120 240928
rect 800 238888 249200 240648
rect 880 238608 249200 238888
rect 800 236848 249200 238608
rect 800 236568 249120 236848
rect 800 235488 249200 236568
rect 880 235208 249200 235488
rect 800 232768 249200 235208
rect 800 232488 249120 232768
rect 800 231408 249200 232488
rect 880 231128 249200 231408
rect 800 229368 249200 231128
rect 800 229088 249120 229368
rect 800 228008 249200 229088
rect 880 227728 249200 228008
rect 800 225288 249200 227728
rect 800 225008 249120 225288
rect 800 223928 249200 225008
rect 880 223648 249200 223928
rect 800 221888 249200 223648
rect 800 221608 249120 221888
rect 800 220528 249200 221608
rect 880 220248 249200 220528
rect 800 217808 249200 220248
rect 800 217528 249120 217808
rect 800 216448 249200 217528
rect 880 216168 249200 216448
rect 800 213728 249200 216168
rect 800 213448 249120 213728
rect 800 212368 249200 213448
rect 880 212088 249200 212368
rect 800 210328 249200 212088
rect 800 210048 249120 210328
rect 800 208968 249200 210048
rect 880 208688 249200 208968
rect 800 206248 249200 208688
rect 800 205968 249120 206248
rect 800 204888 249200 205968
rect 880 204608 249200 204888
rect 800 202848 249200 204608
rect 800 202568 249120 202848
rect 800 201488 249200 202568
rect 880 201208 249200 201488
rect 800 198768 249200 201208
rect 800 198488 249120 198768
rect 800 197408 249200 198488
rect 880 197128 249200 197408
rect 800 194688 249200 197128
rect 800 194408 249120 194688
rect 800 193328 249200 194408
rect 880 193048 249200 193328
rect 800 191288 249200 193048
rect 800 191008 249120 191288
rect 800 189928 249200 191008
rect 880 189648 249200 189928
rect 800 187208 249200 189648
rect 800 186928 249120 187208
rect 800 185848 249200 186928
rect 880 185568 249200 185848
rect 800 183808 249200 185568
rect 800 183528 249120 183808
rect 800 182448 249200 183528
rect 880 182168 249200 182448
rect 800 179728 249200 182168
rect 800 179448 249120 179728
rect 800 178368 249200 179448
rect 880 178088 249200 178368
rect 800 176328 249200 178088
rect 800 176048 249120 176328
rect 800 174288 249200 176048
rect 880 174008 249200 174288
rect 800 172248 249200 174008
rect 800 171968 249120 172248
rect 800 170888 249200 171968
rect 880 170608 249200 170888
rect 800 168168 249200 170608
rect 800 167888 249120 168168
rect 800 166808 249200 167888
rect 880 166528 249200 166808
rect 800 164768 249200 166528
rect 800 164488 249120 164768
rect 800 163408 249200 164488
rect 880 163128 249200 163408
rect 800 160688 249200 163128
rect 800 160408 249120 160688
rect 800 159328 249200 160408
rect 880 159048 249200 159328
rect 800 157288 249200 159048
rect 800 157008 249120 157288
rect 800 155928 249200 157008
rect 880 155648 249200 155928
rect 800 153208 249200 155648
rect 800 152928 249120 153208
rect 800 151848 249200 152928
rect 880 151568 249200 151848
rect 800 149128 249200 151568
rect 800 148848 249120 149128
rect 800 147768 249200 148848
rect 880 147488 249200 147768
rect 800 145728 249200 147488
rect 800 145448 249120 145728
rect 800 144368 249200 145448
rect 880 144088 249200 144368
rect 800 141648 249200 144088
rect 800 141368 249120 141648
rect 800 140288 249200 141368
rect 880 140008 249200 140288
rect 800 138248 249200 140008
rect 800 137968 249120 138248
rect 800 136888 249200 137968
rect 880 136608 249200 136888
rect 800 134168 249200 136608
rect 800 133888 249120 134168
rect 800 132808 249200 133888
rect 880 132528 249200 132808
rect 800 130768 249200 132528
rect 800 130488 249120 130768
rect 800 128728 249200 130488
rect 880 128448 249200 128728
rect 800 126688 249200 128448
rect 800 126408 249120 126688
rect 800 125328 249200 126408
rect 880 125048 249200 125328
rect 800 122608 249200 125048
rect 800 122328 249120 122608
rect 800 121248 249200 122328
rect 880 120968 249200 121248
rect 800 119208 249200 120968
rect 800 118928 249120 119208
rect 800 117848 249200 118928
rect 880 117568 249200 117848
rect 800 115128 249200 117568
rect 800 114848 249120 115128
rect 800 113768 249200 114848
rect 880 113488 249200 113768
rect 800 111728 249200 113488
rect 800 111448 249120 111728
rect 800 110368 249200 111448
rect 880 110088 249200 110368
rect 800 107648 249200 110088
rect 800 107368 249120 107648
rect 800 106288 249200 107368
rect 880 106008 249200 106288
rect 800 103568 249200 106008
rect 800 103288 249120 103568
rect 800 102208 249200 103288
rect 880 101928 249200 102208
rect 800 100168 249200 101928
rect 800 99888 249120 100168
rect 800 98808 249200 99888
rect 880 98528 249200 98808
rect 800 96088 249200 98528
rect 800 95808 249120 96088
rect 800 94728 249200 95808
rect 880 94448 249200 94728
rect 800 92688 249200 94448
rect 800 92408 249120 92688
rect 800 91328 249200 92408
rect 880 91048 249200 91328
rect 800 88608 249200 91048
rect 800 88328 249120 88608
rect 800 87248 249200 88328
rect 880 86968 249200 87248
rect 800 84528 249200 86968
rect 800 84248 249120 84528
rect 800 83168 249200 84248
rect 880 82888 249200 83168
rect 800 81128 249200 82888
rect 800 80848 249120 81128
rect 800 79768 249200 80848
rect 880 79488 249200 79768
rect 800 77048 249200 79488
rect 800 76768 249120 77048
rect 800 75688 249200 76768
rect 880 75408 249200 75688
rect 800 73648 249200 75408
rect 800 73368 249120 73648
rect 800 72288 249200 73368
rect 880 72008 249200 72288
rect 800 69568 249200 72008
rect 800 69288 249120 69568
rect 800 68208 249200 69288
rect 880 67928 249200 68208
rect 800 66168 249200 67928
rect 800 65888 249120 66168
rect 800 64128 249200 65888
rect 880 63848 249200 64128
rect 800 62088 249200 63848
rect 800 61808 249120 62088
rect 800 60728 249200 61808
rect 880 60448 249200 60728
rect 800 58008 249200 60448
rect 800 57728 249120 58008
rect 800 56648 249200 57728
rect 880 56368 249200 56648
rect 800 54608 249200 56368
rect 800 54328 249120 54608
rect 800 53248 249200 54328
rect 880 52968 249200 53248
rect 800 50528 249200 52968
rect 800 50248 249120 50528
rect 800 49168 249200 50248
rect 880 48888 249200 49168
rect 800 47128 249200 48888
rect 800 46848 249120 47128
rect 800 45768 249200 46848
rect 880 45488 249200 45768
rect 800 43048 249200 45488
rect 800 42768 249120 43048
rect 800 41688 249200 42768
rect 880 41408 249200 41688
rect 800 38968 249200 41408
rect 800 38688 249120 38968
rect 800 37608 249200 38688
rect 880 37328 249200 37608
rect 800 35568 249200 37328
rect 800 35288 249120 35568
rect 800 34208 249200 35288
rect 880 33928 249200 34208
rect 800 31488 249200 33928
rect 800 31208 249120 31488
rect 800 30128 249200 31208
rect 880 29848 249200 30128
rect 800 28088 249200 29848
rect 800 27808 249120 28088
rect 800 26728 249200 27808
rect 880 26448 249200 26728
rect 800 24008 249200 26448
rect 800 23728 249120 24008
rect 800 22648 249200 23728
rect 880 22368 249200 22648
rect 800 20608 249200 22368
rect 800 20328 249120 20608
rect 800 18568 249200 20328
rect 880 18288 249200 18568
rect 800 16528 249200 18288
rect 800 16248 249120 16528
rect 800 15168 249200 16248
rect 880 14888 249200 15168
rect 800 12448 249200 14888
rect 800 12168 249120 12448
rect 800 11088 249200 12168
rect 880 10808 249200 11088
rect 800 9048 249200 10808
rect 800 8768 249120 9048
rect 800 7688 249200 8768
rect 880 7408 249200 7688
rect 800 4968 249200 7408
rect 800 4688 249120 4968
rect 800 3608 249200 4688
rect 880 3328 249200 3608
rect 800 1568 249200 3328
rect 800 1288 249120 1568
rect 800 171 249200 1288
<< metal4 >>
rect 4208 2128 4528 247568
rect 19568 2128 19888 247568
rect 34928 2128 35248 247568
rect 50288 2128 50608 247568
rect 65648 2128 65968 247568
rect 81008 2128 81328 247568
rect 96368 2128 96688 247568
rect 111728 2128 112048 247568
rect 127088 2128 127408 247568
rect 142448 2128 142768 247568
rect 157808 2128 158128 247568
rect 173168 2128 173488 247568
rect 188528 2128 188848 247568
rect 203888 2128 204208 247568
rect 219248 2128 219568 247568
rect 234608 2128 234928 247568
<< obsm4 >>
rect 8155 2048 19488 247213
rect 19968 2048 34848 247213
rect 35328 2048 50208 247213
rect 50688 2048 65568 247213
rect 66048 2048 80928 247213
rect 81408 2048 96288 247213
rect 96768 2048 111648 247213
rect 112128 2048 127008 247213
rect 127488 2048 132605 247213
rect 8155 171 132605 2048
<< labels >>
rlabel metal2 s 90178 249200 90234 250000 6 alu_output[0]
port 1 nsew signal output
rlabel metal2 s 104346 0 104402 800 6 alu_output[10]
port 2 nsew signal output
rlabel metal2 s 43166 249200 43222 250000 6 alu_output[11]
port 3 nsew signal output
rlabel metal2 s 21914 249200 21970 250000 6 alu_output[12]
port 4 nsew signal output
rlabel metal2 s 57978 249200 58034 250000 6 alu_output[13]
port 5 nsew signal output
rlabel metal2 s 180338 249200 180394 250000 6 alu_output[14]
port 6 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 alu_output[15]
port 7 nsew signal output
rlabel metal3 s 0 91128 800 91248 6 alu_output[16]
port 8 nsew signal output
rlabel metal3 s 249200 73448 250000 73568 6 alu_output[17]
port 9 nsew signal output
rlabel metal2 s 190642 249200 190698 250000 6 alu_output[18]
port 10 nsew signal output
rlabel metal3 s 249200 38768 250000 38888 6 alu_output[19]
port 11 nsew signal output
rlabel metal2 s 193862 0 193918 800 6 alu_output[1]
port 12 nsew signal output
rlabel metal3 s 249200 145528 250000 145648 6 alu_output[20]
port 13 nsew signal output
rlabel metal2 s 197726 249200 197782 250000 6 alu_output[21]
port 14 nsew signal output
rlabel metal3 s 0 204688 800 204808 6 alu_output[22]
port 15 nsew signal output
rlabel metal3 s 249200 31288 250000 31408 6 alu_output[23]
port 16 nsew signal output
rlabel metal2 s 212538 249200 212594 250000 6 alu_output[24]
port 17 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 alu_output[25]
port 18 nsew signal output
rlabel metal2 s 25134 249200 25190 250000 6 alu_output[26]
port 19 nsew signal output
rlabel metal3 s 249200 213528 250000 213648 6 alu_output[27]
port 20 nsew signal output
rlabel metal3 s 249200 153008 250000 153128 6 alu_output[28]
port 21 nsew signal output
rlabel metal2 s 244738 249200 244794 250000 6 alu_output[29]
port 22 nsew signal output
rlabel metal2 s 122378 249200 122434 250000 6 alu_output[2]
port 23 nsew signal output
rlabel metal3 s 0 178168 800 178288 6 alu_output[30]
port 24 nsew signal output
rlabel metal3 s 249200 1368 250000 1488 6 alu_output[31]
port 25 nsew signal output
rlabel metal2 s 54114 249200 54170 250000 6 alu_output[3]
port 26 nsew signal output
rlabel metal2 s 126242 249200 126298 250000 6 alu_output[4]
port 27 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 alu_output[5]
port 28 nsew signal output
rlabel metal2 s 229926 0 229982 800 6 alu_output[6]
port 29 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 alu_output[7]
port 30 nsew signal output
rlabel metal2 s 151358 249200 151414 250000 6 alu_output[8]
port 31 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 alu_output[9]
port 32 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 clk
port 33 nsew signal input
rlabel metal2 s 140410 249200 140466 250000 6 funct3[0]
port 34 nsew signal input
rlabel metal3 s 249200 126488 250000 126608 6 funct3[1]
port 35 nsew signal input
rlabel metal2 s 190642 0 190698 800 6 funct3[2]
port 36 nsew signal input
rlabel metal3 s 249200 130568 250000 130688 6 funct7[0]
port 37 nsew signal input
rlabel metal3 s 249200 99968 250000 100088 6 funct7[1]
port 38 nsew signal input
rlabel metal3 s 249200 225088 250000 225208 6 funct7[2]
port 39 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 funct7[3]
port 40 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 funct7[4]
port 41 nsew signal input
rlabel metal3 s 0 197208 800 197328 6 funct7[5]
port 42 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 funct7[6]
port 43 nsew signal input
rlabel metal2 s 201590 249200 201646 250000 6 immediate[0]
port 44 nsew signal input
rlabel metal2 s 211894 0 211950 800 6 immediate[10]
port 45 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 immediate[11]
port 46 nsew signal input
rlabel metal2 s 200946 0 201002 800 6 immediate[12]
port 47 nsew signal input
rlabel metal2 s 150714 0 150770 800 6 immediate[13]
port 48 nsew signal input
rlabel metal3 s 0 174088 800 174208 6 immediate[14]
port 49 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 immediate[15]
port 50 nsew signal input
rlabel metal2 s 158442 249200 158498 250000 6 immediate[16]
port 51 nsew signal input
rlabel metal2 s 247958 0 248014 800 6 immediate[17]
port 52 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 immediate[18]
port 53 nsew signal input
rlabel metal2 s 179694 0 179750 800 6 immediate[19]
port 54 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 immediate[1]
port 55 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 immediate[20]
port 56 nsew signal input
rlabel metal3 s 0 132608 800 132728 6 immediate[21]
port 57 nsew signal input
rlabel metal2 s 119158 249200 119214 250000 6 immediate[22]
port 58 nsew signal input
rlabel metal3 s 249200 202648 250000 202768 6 immediate[23]
port 59 nsew signal input
rlabel metal2 s 108210 249200 108266 250000 6 immediate[24]
port 60 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 immediate[25]
port 61 nsew signal input
rlabel metal2 s 137190 249200 137246 250000 6 immediate[26]
port 62 nsew signal input
rlabel metal2 s 18050 249200 18106 250000 6 immediate[27]
port 63 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 immediate[28]
port 64 nsew signal input
rlabel metal2 s 86314 249200 86370 250000 6 immediate[29]
port 65 nsew signal input
rlabel metal3 s 0 216248 800 216368 6 immediate[2]
port 66 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 immediate[30]
port 67 nsew signal input
rlabel metal3 s 249200 12248 250000 12368 6 immediate[31]
port 68 nsew signal input
rlabel metal2 s 104346 249200 104402 250000 6 immediate[3]
port 69 nsew signal input
rlabel metal3 s 0 128528 800 128648 6 immediate[4]
port 70 nsew signal input
rlabel metal2 s 3882 249200 3938 250000 6 immediate[5]
port 71 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 immediate[6]
port 72 nsew signal input
rlabel metal2 s 183558 249200 183614 250000 6 immediate[7]
port 73 nsew signal input
rlabel metal2 s 233790 249200 233846 250000 6 immediate[8]
port 74 nsew signal input
rlabel metal3 s 249200 210128 250000 210248 6 immediate[9]
port 75 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 immediate_sel
port 76 nsew signal input
rlabel metal3 s 249200 114928 250000 115048 6 instruction_type[0]
port 77 nsew signal input
rlabel metal3 s 249200 236648 250000 236768 6 instruction_type[1]
port 78 nsew signal input
rlabel metal3 s 249200 167968 250000 168088 6 instruction_type[2]
port 79 nsew signal input
rlabel metal2 s 28998 249200 29054 250000 6 instruction_type[3]
port 80 nsew signal input
rlabel metal2 s 139766 0 139822 800 6 instruction_type[4]
port 81 nsew signal input
rlabel metal3 s 0 189728 800 189848 6 instruction_type[5]
port 82 nsew signal input
rlabel metal3 s 249200 191088 250000 191208 6 la_read_data[0]
port 83 nsew signal output
rlabel metal2 s 129462 249200 129518 250000 6 la_read_data[10]
port 84 nsew signal output
rlabel metal3 s 0 227808 800 227928 6 la_read_data[11]
port 85 nsew signal output
rlabel metal2 s 222842 0 222898 800 6 la_read_data[12]
port 86 nsew signal output
rlabel metal3 s 0 220328 800 220448 6 la_read_data[13]
port 87 nsew signal output
rlabel metal2 s 14830 249200 14886 250000 6 la_read_data[14]
port 88 nsew signal output
rlabel metal2 s 226062 0 226118 800 6 la_read_data[15]
port 89 nsew signal output
rlabel metal3 s 249200 65968 250000 66088 6 la_read_data[16]
port 90 nsew signal output
rlabel metal3 s 249200 133968 250000 134088 6 la_read_data[17]
port 91 nsew signal output
rlabel metal3 s 249200 138048 250000 138168 6 la_read_data[18]
port 92 nsew signal output
rlabel metal3 s 0 201288 800 201408 6 la_read_data[19]
port 93 nsew signal output
rlabel metal2 s 165526 249200 165582 250000 6 la_read_data[1]
port 94 nsew signal output
rlabel metal2 s 7102 249200 7158 250000 6 la_read_data[20]
port 95 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 la_read_data[21]
port 96 nsew signal output
rlabel metal2 s 218978 0 219034 800 6 la_read_data[22]
port 97 nsew signal output
rlabel metal2 s 204810 0 204866 800 6 la_read_data[23]
port 98 nsew signal output
rlabel metal3 s 0 125128 800 125248 6 la_read_data[24]
port 99 nsew signal output
rlabel metal3 s 0 170688 800 170808 6 la_read_data[25]
port 100 nsew signal output
rlabel metal3 s 0 208768 800 208888 6 la_read_data[26]
port 101 nsew signal output
rlabel metal2 s 244094 0 244150 800 6 la_read_data[27]
port 102 nsew signal output
rlabel metal2 s 72146 249200 72202 250000 6 la_read_data[28]
port 103 nsew signal output
rlabel metal2 s 237654 249200 237710 250000 6 la_read_data[29]
port 104 nsew signal output
rlabel metal2 s 68282 249200 68338 250000 6 la_read_data[2]
port 105 nsew signal output
rlabel metal3 s 249200 244128 250000 244248 6 la_read_data[30]
port 106 nsew signal output
rlabel metal3 s 0 238688 800 238808 6 la_read_data[31]
port 107 nsew signal output
rlabel metal2 s 172610 0 172666 800 6 la_read_data[3]
port 108 nsew signal output
rlabel metal3 s 0 147568 800 147688 6 la_read_data[4]
port 109 nsew signal output
rlabel metal2 s 61198 249200 61254 250000 6 la_read_data[5]
port 110 nsew signal output
rlabel metal2 s 111430 249200 111486 250000 6 la_read_data[6]
port 111 nsew signal output
rlabel metal3 s 249200 122408 250000 122528 6 la_read_data[7]
port 112 nsew signal output
rlabel metal3 s 0 246848 800 246968 6 la_read_data[8]
port 113 nsew signal output
rlabel metal3 s 249200 16328 250000 16448 6 la_read_data[9]
port 114 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 la_reg_select[0]
port 115 nsew signal input
rlabel metal3 s 249200 141448 250000 141568 6 la_reg_select[1]
port 116 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 la_reg_select[2]
port 117 nsew signal input
rlabel metal2 s 79230 249200 79286 250000 6 la_reg_select[3]
port 118 nsew signal input
rlabel metal3 s 0 159128 800 159248 6 la_reg_select[4]
port 119 nsew signal input
rlabel metal3 s 249200 92488 250000 92608 6 opcode[0]
port 120 nsew signal input
rlabel metal3 s 249200 69368 250000 69488 6 opcode[1]
port 121 nsew signal input
rlabel metal3 s 249200 198568 250000 198688 6 opcode[2]
port 122 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 opcode[3]
port 123 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 opcode[4]
port 124 nsew signal input
rlabel metal2 s 76010 249200 76066 250000 6 opcode[5]
port 125 nsew signal input
rlabel metal3 s 0 136688 800 136808 6 opcode[6]
port 126 nsew signal input
rlabel metal3 s 0 106088 800 106208 6 pc[0]
port 127 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 pc[10]
port 128 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 pc[11]
port 129 nsew signal input
rlabel metal2 s 219622 249200 219678 250000 6 pc[12]
port 130 nsew signal input
rlabel metal3 s 0 56448 800 56568 6 pc[13]
port 131 nsew signal input
rlabel metal2 s 97262 249200 97318 250000 6 pc[14]
port 132 nsew signal input
rlabel metal2 s 50250 249200 50306 250000 6 pc[15]
port 133 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 pc[16]
port 134 nsew signal input
rlabel metal3 s 0 166608 800 166728 6 pc[17]
port 135 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 pc[18]
port 136 nsew signal input
rlabel metal3 s 249200 148928 250000 149048 6 pc[19]
port 137 nsew signal input
rlabel metal3 s 0 235288 800 235408 6 pc[1]
port 138 nsew signal input
rlabel metal2 s 10966 249200 11022 250000 6 pc[20]
port 139 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 pc[21]
port 140 nsew signal input
rlabel metal3 s 249200 23808 250000 23928 6 pc[22]
port 141 nsew signal input
rlabel metal3 s 249200 61888 250000 62008 6 pc[23]
port 142 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 pc[24]
port 143 nsew signal input
rlabel metal2 s 241518 249200 241574 250000 6 pc[25]
port 144 nsew signal input
rlabel metal2 s 182914 0 182970 800 6 pc[26]
port 145 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 pc[27]
port 146 nsew signal input
rlabel metal3 s 0 151648 800 151768 6 pc[28]
port 147 nsew signal input
rlabel metal3 s 249200 35368 250000 35488 6 pc[29]
port 148 nsew signal input
rlabel metal3 s 0 41488 800 41608 6 pc[2]
port 149 nsew signal input
rlabel metal3 s 249200 160488 250000 160608 6 pc[30]
port 150 nsew signal input
rlabel metal2 s 208674 0 208730 800 6 pc[31]
port 151 nsew signal input
rlabel metal3 s 0 231208 800 231328 6 pc[3]
port 152 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 pc[4]
port 153 nsew signal input
rlabel metal2 s 162306 249200 162362 250000 6 pc[5]
port 154 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 pc[6]
port 155 nsew signal input
rlabel metal3 s 249200 42848 250000 42968 6 pc[7]
port 156 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 pc[8]
port 157 nsew signal input
rlabel metal3 s 249200 76848 250000 76968 6 pc[9]
port 158 nsew signal input
rlabel metal3 s 0 82968 800 83088 6 rd[0]
port 159 nsew signal input
rlabel metal3 s 0 182248 800 182368 6 rd[1]
port 160 nsew signal input
rlabel metal3 s 0 121048 800 121168 6 rd[2]
port 161 nsew signal input
rlabel metal3 s 249200 179528 250000 179648 6 rd[3]
port 162 nsew signal input
rlabel metal3 s 249200 103368 250000 103488 6 rd[4]
port 163 nsew signal input
rlabel metal2 s 194506 249200 194562 250000 6 read_data[0]
port 164 nsew signal input
rlabel metal2 s 208674 249200 208730 250000 6 read_data[10]
port 165 nsew signal input
rlabel metal2 s 233790 0 233846 800 6 read_data[11]
port 166 nsew signal input
rlabel metal2 s 65062 249200 65118 250000 6 read_data[12]
port 167 nsew signal input
rlabel metal2 s 101126 249200 101182 250000 6 read_data[13]
port 168 nsew signal input
rlabel metal3 s 249200 229168 250000 229288 6 read_data[14]
port 169 nsew signal input
rlabel metal2 s 223486 249200 223542 250000 6 read_data[15]
port 170 nsew signal input
rlabel metal2 s 144274 249200 144330 250000 6 read_data[16]
port 171 nsew signal input
rlabel metal3 s 0 144168 800 144288 6 read_data[17]
port 172 nsew signal input
rlabel metal3 s 0 163208 800 163328 6 read_data[18]
port 173 nsew signal input
rlabel metal3 s 249200 107448 250000 107568 6 read_data[19]
port 174 nsew signal input
rlabel metal3 s 249200 95888 250000 96008 6 read_data[1]
port 175 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 read_data[20]
port 176 nsew signal input
rlabel metal3 s 249200 84328 250000 84448 6 read_data[21]
port 177 nsew signal input
rlabel metal3 s 249200 20408 250000 20528 6 read_data[22]
port 178 nsew signal input
rlabel metal2 s 197726 0 197782 800 6 read_data[23]
port 179 nsew signal input
rlabel metal3 s 249200 248208 250000 248328 6 read_data[24]
port 180 nsew signal input
rlabel metal3 s 249200 187008 250000 187128 6 read_data[25]
port 181 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 read_data[26]
port 182 nsew signal input
rlabel metal2 s 168746 0 168802 800 6 read_data[27]
port 183 nsew signal input
rlabel metal3 s 249200 4768 250000 4888 6 read_data[28]
port 184 nsew signal input
rlabel metal2 s 133326 249200 133382 250000 6 read_data[29]
port 185 nsew signal input
rlabel metal2 s 114650 0 114706 800 6 read_data[2]
port 186 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 read_data[30]
port 187 nsew signal input
rlabel metal2 s 176474 249200 176530 250000 6 read_data[31]
port 188 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 read_data[3]
port 189 nsew signal input
rlabel metal3 s 249200 172048 250000 172168 6 read_data[4]
port 190 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 read_data[5]
port 191 nsew signal input
rlabel metal3 s 249200 232568 250000 232688 6 read_data[6]
port 192 nsew signal input
rlabel metal3 s 249200 54408 250000 54528 6 read_data[7]
port 193 nsew signal input
rlabel metal2 s 164882 0 164938 800 6 read_data[8]
port 194 nsew signal input
rlabel metal3 s 249200 240728 250000 240848 6 read_data[9]
port 195 nsew signal input
rlabel metal2 s 161662 0 161718 800 6 reg_write
port 196 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 rs1[0]
port 197 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 rs1[1]
port 198 nsew signal input
rlabel metal2 s 215758 0 215814 800 6 rs1[2]
port 199 nsew signal input
rlabel metal3 s 249200 27888 250000 28008 6 rs1[3]
port 200 nsew signal input
rlabel metal2 s 154578 249200 154634 250000 6 rs1[4]
port 201 nsew signal input
rlabel metal3 s 249200 164568 250000 164688 6 rs1_data[0]
port 202 nsew signal output
rlabel metal2 s 32862 249200 32918 250000 6 rs1_data[10]
port 203 nsew signal output
rlabel metal2 s 47030 249200 47086 250000 6 rs1_data[11]
port 204 nsew signal output
rlabel metal2 s 39946 249200 40002 250000 6 rs1_data[12]
port 205 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 rs1_data[13]
port 206 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 rs1_data[14]
port 207 nsew signal output
rlabel metal3 s 249200 88408 250000 88528 6 rs1_data[15]
port 208 nsew signal output
rlabel metal2 s 125598 0 125654 800 6 rs1_data[16]
port 209 nsew signal output
rlabel metal2 s 226706 249200 226762 250000 6 rs1_data[17]
port 210 nsew signal output
rlabel metal3 s 249200 221688 250000 221808 6 rs1_data[18]
port 211 nsew signal output
rlabel metal2 s 83094 249200 83150 250000 6 rs1_data[19]
port 212 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 rs1_data[1]
port 213 nsew signal output
rlabel metal3 s 249200 111528 250000 111648 6 rs1_data[20]
port 214 nsew signal output
rlabel metal3 s 249200 217608 250000 217728 6 rs1_data[21]
port 215 nsew signal output
rlabel metal3 s 0 223728 800 223848 6 rs1_data[22]
port 216 nsew signal output
rlabel metal3 s 249200 157088 250000 157208 6 rs1_data[23]
port 217 nsew signal output
rlabel metal3 s 249200 50328 250000 50448 6 rs1_data[24]
port 218 nsew signal output
rlabel metal2 s 154578 0 154634 800 6 rs1_data[25]
port 219 nsew signal output
rlabel metal2 s 248602 249200 248658 250000 6 rs1_data[26]
port 220 nsew signal output
rlabel metal2 s 115294 249200 115350 250000 6 rs1_data[27]
port 221 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 rs1_data[28]
port 222 nsew signal output
rlabel metal3 s 0 140088 800 140208 6 rs1_data[29]
port 223 nsew signal output
rlabel metal3 s 0 102008 800 102128 6 rs1_data[2]
port 224 nsew signal output
rlabel metal3 s 249200 46928 250000 47048 6 rs1_data[30]
port 225 nsew signal output
rlabel metal3 s 0 193128 800 193248 6 rs1_data[31]
port 226 nsew signal output
rlabel metal2 s 237010 0 237066 800 6 rs1_data[3]
port 227 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 rs1_data[4]
port 228 nsew signal output
rlabel metal2 s 111430 0 111486 800 6 rs1_data[5]
port 229 nsew signal output
rlabel metal3 s 249200 80928 250000 81048 6 rs1_data[6]
port 230 nsew signal output
rlabel metal2 s 230570 249200 230626 250000 6 rs1_data[7]
port 231 nsew signal output
rlabel metal3 s 249200 194488 250000 194608 6 rs1_data[8]
port 232 nsew signal output
rlabel metal2 s 240874 0 240930 800 6 rs1_data[9]
port 233 nsew signal output
rlabel metal3 s 0 79568 800 79688 6 rs2[0]
port 234 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 rs2[1]
port 235 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 rs2[2]
port 236 nsew signal input
rlabel metal3 s 249200 206048 250000 206168 6 rs2[3]
port 237 nsew signal input
rlabel metal2 s 215758 249200 215814 250000 6 rs2[4]
port 238 nsew signal input
rlabel metal3 s 249200 8848 250000 8968 6 rs2_data[0]
port 239 nsew signal output
rlabel metal2 s 205454 249200 205510 250000 6 rs2_data[10]
port 240 nsew signal output
rlabel metal3 s 0 110168 800 110288 6 rs2_data[11]
port 241 nsew signal output
rlabel metal3 s 0 117648 800 117768 6 rs2_data[12]
port 242 nsew signal output
rlabel metal2 s 157798 0 157854 800 6 rs2_data[13]
port 243 nsew signal output
rlabel metal2 s 18 0 74 800 6 rs2_data[14]
port 244 nsew signal output
rlabel metal2 s 186778 0 186834 800 6 rs2_data[15]
port 245 nsew signal output
rlabel metal3 s 0 155728 800 155848 6 rs2_data[16]
port 246 nsew signal output
rlabel metal2 s 18 249200 74 250000 6 rs2_data[17]
port 247 nsew signal output
rlabel metal3 s 0 72088 800 72208 6 rs2_data[18]
port 248 nsew signal output
rlabel metal3 s 0 113568 800 113688 6 rs2_data[19]
port 249 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 rs2_data[1]
port 250 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 rs2_data[20]
port 251 nsew signal output
rlabel metal2 s 147494 249200 147550 250000 6 rs2_data[21]
port 252 nsew signal output
rlabel metal2 s 93398 249200 93454 250000 6 rs2_data[22]
port 253 nsew signal output
rlabel metal2 s 129462 0 129518 800 6 rs2_data[23]
port 254 nsew signal output
rlabel metal2 s 187422 249200 187478 250000 6 rs2_data[24]
port 255 nsew signal output
rlabel metal3 s 249200 57808 250000 57928 6 rs2_data[25]
port 256 nsew signal output
rlabel metal3 s 0 185648 800 185768 6 rs2_data[26]
port 257 nsew signal output
rlabel metal3 s 249200 183608 250000 183728 6 rs2_data[27]
port 258 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 rs2_data[28]
port 259 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 rs2_data[29]
port 260 nsew signal output
rlabel metal2 s 143630 0 143686 800 6 rs2_data[2]
port 261 nsew signal output
rlabel metal3 s 249200 176128 250000 176248 6 rs2_data[30]
port 262 nsew signal output
rlabel metal2 s 147494 0 147550 800 6 rs2_data[31]
port 263 nsew signal output
rlabel metal2 s 172610 249200 172666 250000 6 rs2_data[3]
port 264 nsew signal output
rlabel metal2 s 169390 249200 169446 250000 6 rs2_data[4]
port 265 nsew signal output
rlabel metal3 s 0 242768 800 242888 6 rs2_data[5]
port 266 nsew signal output
rlabel metal2 s 36082 249200 36138 250000 6 rs2_data[6]
port 267 nsew signal output
rlabel metal2 s 175830 0 175886 800 6 rs2_data[7]
port 268 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 rs2_data[8]
port 269 nsew signal output
rlabel metal3 s 0 212168 800 212288 6 rs2_data[9]
port 270 nsew signal output
rlabel metal3 s 249200 119008 250000 119128 6 rst_n
port 271 nsew signal input
rlabel metal4 s 4208 2128 4528 247568 6 vccd1
port 272 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 247568 6 vccd1
port 272 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 247568 6 vccd1
port 272 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 247568 6 vccd1
port 272 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 247568 6 vccd1
port 272 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 247568 6 vccd1
port 272 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 247568 6 vccd1
port 272 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 247568 6 vccd1
port 272 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 247568 6 vssd1
port 273 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 247568 6 vssd1
port 273 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 247568 6 vssd1
port 273 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 247568 6 vssd1
port 273 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 247568 6 vssd1
port 273 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 247568 6 vssd1
port 273 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 247568 6 vssd1
port 273 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 247568 6 vssd1
port 273 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 250000 250000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 44801716
string GDS_FILE /home/drewarosa/RISC-V-Single-Cycle-CPU-Core/openlane/ALU/runs/22_09_20_15_38/results/signoff/ALU.magic.gds
string GDS_START 894054
<< end >>

