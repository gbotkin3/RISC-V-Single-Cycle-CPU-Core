magic
tech sky130B
magscale 1 2
timestamp 1663699927
<< obsli1 >>
rect 1104 2159 48852 47345
<< obsm1 >>
rect 14 1776 49666 47796
<< metal2 >>
rect 18 49200 74 50000
rect 1950 49200 2006 50000
rect 3882 49200 3938 50000
rect 5814 49200 5870 50000
rect 7746 49200 7802 50000
rect 9678 49200 9734 50000
rect 11610 49200 11666 50000
rect 13542 49200 13598 50000
rect 15474 49200 15530 50000
rect 17406 49200 17462 50000
rect 19338 49200 19394 50000
rect 21270 49200 21326 50000
rect 23202 49200 23258 50000
rect 25134 49200 25190 50000
rect 27066 49200 27122 50000
rect 28998 49200 29054 50000
rect 30930 49200 30986 50000
rect 32862 49200 32918 50000
rect 34794 49200 34850 50000
rect 36726 49200 36782 50000
rect 38658 49200 38714 50000
rect 40590 49200 40646 50000
rect 42522 49200 42578 50000
rect 44454 49200 44510 50000
rect 46386 49200 46442 50000
rect 48318 49200 48374 50000
rect 49606 49200 49662 50000
rect 18 0 74 800
rect 1306 0 1362 800
rect 3238 0 3294 800
rect 5170 0 5226 800
rect 7102 0 7158 800
rect 9034 0 9090 800
rect 10966 0 11022 800
rect 12898 0 12954 800
rect 14830 0 14886 800
rect 16762 0 16818 800
rect 18694 0 18750 800
rect 20626 0 20682 800
rect 22558 0 22614 800
rect 24490 0 24546 800
rect 26422 0 26478 800
rect 28354 0 28410 800
rect 30286 0 30342 800
rect 32218 0 32274 800
rect 34150 0 34206 800
rect 36082 0 36138 800
rect 38014 0 38070 800
rect 39946 0 40002 800
rect 41878 0 41934 800
rect 43810 0 43866 800
rect 45742 0 45798 800
rect 47674 0 47730 800
rect 49606 0 49662 800
<< obsm2 >>
rect 130 49144 1894 49314
rect 2062 49144 3826 49314
rect 3994 49144 5758 49314
rect 5926 49144 7690 49314
rect 7858 49144 9622 49314
rect 9790 49144 11554 49314
rect 11722 49144 13486 49314
rect 13654 49144 15418 49314
rect 15586 49144 17350 49314
rect 17518 49144 19282 49314
rect 19450 49144 21214 49314
rect 21382 49144 23146 49314
rect 23314 49144 25078 49314
rect 25246 49144 27010 49314
rect 27178 49144 28942 49314
rect 29110 49144 30874 49314
rect 31042 49144 32806 49314
rect 32974 49144 34738 49314
rect 34906 49144 36670 49314
rect 36838 49144 38602 49314
rect 38770 49144 40534 49314
rect 40702 49144 42466 49314
rect 42634 49144 44398 49314
rect 44566 49144 46330 49314
rect 46498 49144 48262 49314
rect 48430 49144 49550 49314
rect 20 856 49660 49144
rect 130 800 1250 856
rect 1418 800 3182 856
rect 3350 800 5114 856
rect 5282 800 7046 856
rect 7214 800 8978 856
rect 9146 800 10910 856
rect 11078 800 12842 856
rect 13010 800 14774 856
rect 14942 800 16706 856
rect 16874 800 18638 856
rect 18806 800 20570 856
rect 20738 800 22502 856
rect 22670 800 24434 856
rect 24602 800 26366 856
rect 26534 800 28298 856
rect 28466 800 30230 856
rect 30398 800 32162 856
rect 32330 800 34094 856
rect 34262 800 36026 856
rect 36194 800 37958 856
rect 38126 800 39890 856
rect 40058 800 41822 856
rect 41990 800 43754 856
rect 43922 800 45686 856
rect 45854 800 47618 856
rect 47786 800 49550 856
<< metal3 >>
rect 0 48288 800 48408
rect 49200 48288 50000 48408
rect 0 46248 800 46368
rect 49200 46248 50000 46368
rect 0 44208 800 44328
rect 49200 44208 50000 44328
rect 0 42168 800 42288
rect 49200 42168 50000 42288
rect 0 40128 800 40248
rect 49200 40128 50000 40248
rect 0 38088 800 38208
rect 49200 38088 50000 38208
rect 0 36048 800 36168
rect 49200 36048 50000 36168
rect 0 34008 800 34128
rect 49200 34008 50000 34128
rect 0 31968 800 32088
rect 49200 31968 50000 32088
rect 0 29928 800 30048
rect 49200 29928 50000 30048
rect 0 27888 800 28008
rect 49200 27888 50000 28008
rect 0 25848 800 25968
rect 49200 25848 50000 25968
rect 0 23808 800 23928
rect 49200 23808 50000 23928
rect 0 21768 800 21888
rect 49200 21768 50000 21888
rect 0 19728 800 19848
rect 49200 19728 50000 19848
rect 0 17688 800 17808
rect 49200 17688 50000 17808
rect 0 15648 800 15768
rect 49200 15648 50000 15768
rect 0 13608 800 13728
rect 49200 13608 50000 13728
rect 0 11568 800 11688
rect 49200 11568 50000 11688
rect 0 9528 800 9648
rect 49200 9528 50000 9648
rect 0 7488 800 7608
rect 49200 7488 50000 7608
rect 0 5448 800 5568
rect 49200 5448 50000 5568
rect 0 3408 800 3528
rect 49200 3408 50000 3528
rect 0 1368 800 1488
rect 49200 1368 50000 1488
<< obsm3 >>
rect 880 48208 49120 48381
rect 800 46448 49200 48208
rect 880 46168 49120 46448
rect 800 44408 49200 46168
rect 880 44128 49120 44408
rect 800 42368 49200 44128
rect 880 42088 49120 42368
rect 800 40328 49200 42088
rect 880 40048 49120 40328
rect 800 38288 49200 40048
rect 880 38008 49120 38288
rect 800 36248 49200 38008
rect 880 35968 49120 36248
rect 800 34208 49200 35968
rect 880 33928 49120 34208
rect 800 32168 49200 33928
rect 880 31888 49120 32168
rect 800 30128 49200 31888
rect 880 29848 49120 30128
rect 800 28088 49200 29848
rect 880 27808 49120 28088
rect 800 26048 49200 27808
rect 880 25768 49120 26048
rect 800 24008 49200 25768
rect 880 23728 49120 24008
rect 800 21968 49200 23728
rect 880 21688 49120 21968
rect 800 19928 49200 21688
rect 880 19648 49120 19928
rect 800 17888 49200 19648
rect 880 17608 49120 17888
rect 800 15848 49200 17608
rect 880 15568 49120 15848
rect 800 13808 49200 15568
rect 880 13528 49120 13808
rect 800 11768 49200 13528
rect 880 11488 49120 11768
rect 800 9728 49200 11488
rect 880 9448 49120 9728
rect 800 7688 49200 9448
rect 880 7408 49120 7688
rect 800 5648 49200 7408
rect 880 5368 49120 5648
rect 800 3608 49200 5368
rect 880 3328 49120 3608
rect 800 1568 49200 3328
rect 880 1395 49120 1568
<< metal4 >>
rect 4208 2128 4528 47376
rect 19568 2128 19888 47376
rect 34928 2128 35248 47376
<< obsm4 >>
rect 14963 2483 19488 47021
rect 19968 2483 34848 47021
rect 35328 2483 35453 47021
<< labels >>
rlabel metal3 s 49200 7488 50000 7608 6 alu_branch
port 1 nsew signal input
rlabel metal3 s 49200 42168 50000 42288 6 branch
port 2 nsew signal input
rlabel metal2 s 28998 49200 29054 50000 6 clk
port 3 nsew signal input
rlabel metal3 s 49200 48288 50000 48408 6 immediate[0]
port 4 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 immediate[10]
port 5 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 immediate[11]
port 6 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 immediate[12]
port 7 nsew signal input
rlabel metal2 s 48318 49200 48374 50000 6 immediate[13]
port 8 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 immediate[14]
port 9 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 immediate[15]
port 10 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 immediate[16]
port 11 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 immediate[17]
port 12 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 immediate[18]
port 13 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 immediate[19]
port 14 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 immediate[1]
port 15 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 immediate[20]
port 16 nsew signal input
rlabel metal3 s 49200 36048 50000 36168 6 immediate[21]
port 17 nsew signal input
rlabel metal2 s 23202 49200 23258 50000 6 immediate[22]
port 18 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 immediate[23]
port 19 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 immediate[24]
port 20 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 immediate[25]
port 21 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 immediate[26]
port 22 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 immediate[27]
port 23 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 immediate[28]
port 24 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 immediate[29]
port 25 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 immediate[2]
port 26 nsew signal input
rlabel metal3 s 49200 25848 50000 25968 6 immediate[30]
port 27 nsew signal input
rlabel metal2 s 30930 49200 30986 50000 6 immediate[31]
port 28 nsew signal input
rlabel metal2 s 17406 49200 17462 50000 6 immediate[3]
port 29 nsew signal input
rlabel metal3 s 49200 46248 50000 46368 6 immediate[4]
port 30 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 immediate[5]
port 31 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 immediate[6]
port 32 nsew signal input
rlabel metal3 s 49200 44208 50000 44328 6 immediate[7]
port 33 nsew signal input
rlabel metal2 s 19338 49200 19394 50000 6 immediate[8]
port 34 nsew signal input
rlabel metal3 s 49200 11568 50000 11688 6 immediate[9]
port 35 nsew signal input
rlabel metal3 s 49200 15648 50000 15768 6 jump_jal
port 36 nsew signal input
rlabel metal2 s 21270 49200 21326 50000 6 jump_jalr
port 37 nsew signal input
rlabel metal2 s 13542 49200 13598 50000 6 pc_out[0]
port 38 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 pc_out[10]
port 39 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 pc_out[11]
port 40 nsew signal output
rlabel metal3 s 49200 38088 50000 38208 6 pc_out[12]
port 41 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 pc_out[13]
port 42 nsew signal output
rlabel metal3 s 49200 19728 50000 19848 6 pc_out[14]
port 43 nsew signal output
rlabel metal2 s 36726 49200 36782 50000 6 pc_out[15]
port 44 nsew signal output
rlabel metal2 s 15474 49200 15530 50000 6 pc_out[16]
port 45 nsew signal output
rlabel metal3 s 49200 1368 50000 1488 6 pc_out[17]
port 46 nsew signal output
rlabel metal3 s 49200 40128 50000 40248 6 pc_out[18]
port 47 nsew signal output
rlabel metal2 s 46386 49200 46442 50000 6 pc_out[19]
port 48 nsew signal output
rlabel metal2 s 27066 49200 27122 50000 6 pc_out[1]
port 49 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 pc_out[20]
port 50 nsew signal output
rlabel metal3 s 49200 9528 50000 9648 6 pc_out[21]
port 51 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 pc_out[22]
port 52 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 pc_out[23]
port 53 nsew signal output
rlabel metal2 s 32862 49200 32918 50000 6 pc_out[24]
port 54 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 pc_out[25]
port 55 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 pc_out[26]
port 56 nsew signal output
rlabel metal2 s 42522 49200 42578 50000 6 pc_out[27]
port 57 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 pc_out[28]
port 58 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 pc_out[29]
port 59 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 pc_out[2]
port 60 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 pc_out[30]
port 61 nsew signal output
rlabel metal3 s 49200 21768 50000 21888 6 pc_out[31]
port 62 nsew signal output
rlabel metal3 s 49200 13608 50000 13728 6 pc_out[3]
port 63 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 pc_out[4]
port 64 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 pc_out[5]
port 65 nsew signal output
rlabel metal3 s 49200 3408 50000 3528 6 pc_out[6]
port 66 nsew signal output
rlabel metal2 s 5814 49200 5870 50000 6 pc_out[7]
port 67 nsew signal output
rlabel metal3 s 49200 17688 50000 17808 6 pc_out[8]
port 68 nsew signal output
rlabel metal3 s 49200 31968 50000 32088 6 pc_out[9]
port 69 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 rs1_data[0]
port 70 nsew signal input
rlabel metal3 s 49200 34008 50000 34128 6 rs1_data[10]
port 71 nsew signal input
rlabel metal2 s 7746 49200 7802 50000 6 rs1_data[11]
port 72 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 rs1_data[12]
port 73 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 rs1_data[13]
port 74 nsew signal input
rlabel metal2 s 18 0 74 800 6 rs1_data[14]
port 75 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 rs1_data[15]
port 76 nsew signal input
rlabel metal2 s 9678 49200 9734 50000 6 rs1_data[16]
port 77 nsew signal input
rlabel metal2 s 25134 49200 25190 50000 6 rs1_data[17]
port 78 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 rs1_data[18]
port 79 nsew signal input
rlabel metal2 s 18 49200 74 50000 6 rs1_data[19]
port 80 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 rs1_data[1]
port 81 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 rs1_data[20]
port 82 nsew signal input
rlabel metal2 s 44454 49200 44510 50000 6 rs1_data[21]
port 83 nsew signal input
rlabel metal2 s 34794 49200 34850 50000 6 rs1_data[22]
port 84 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 rs1_data[23]
port 85 nsew signal input
rlabel metal2 s 49606 49200 49662 50000 6 rs1_data[24]
port 86 nsew signal input
rlabel metal3 s 49200 5448 50000 5568 6 rs1_data[25]
port 87 nsew signal input
rlabel metal2 s 1950 49200 2006 50000 6 rs1_data[26]
port 88 nsew signal input
rlabel metal3 s 49200 27888 50000 28008 6 rs1_data[27]
port 89 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 rs1_data[28]
port 90 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 rs1_data[29]
port 91 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 rs1_data[2]
port 92 nsew signal input
rlabel metal3 s 49200 29928 50000 30048 6 rs1_data[30]
port 93 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 rs1_data[31]
port 94 nsew signal input
rlabel metal2 s 40590 49200 40646 50000 6 rs1_data[3]
port 95 nsew signal input
rlabel metal2 s 38658 49200 38714 50000 6 rs1_data[4]
port 96 nsew signal input
rlabel metal2 s 3882 49200 3938 50000 6 rs1_data[5]
port 97 nsew signal input
rlabel metal2 s 11610 49200 11666 50000 6 rs1_data[6]
port 98 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 rs1_data[7]
port 99 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 rs1_data[8]
port 100 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 rs1_data[9]
port 101 nsew signal input
rlabel metal3 s 49200 23808 50000 23928 6 rst_n
port 102 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 103 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 103 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 104 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 50000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3562972
string GDS_FILE /home/drewarosa/RISC-V-Single-Cycle-CPU-Core/openlane/pc/runs/22_09_20_14_49/results/signoff/pc.magic.gds
string GDS_START 531454
<< end >>

