magic
tech sky130B
magscale 1 2
timestamp 1661896804
<< obsli1 >>
rect 1104 2159 221352 221969
<< obsm1 >>
rect 1104 2128 221352 222000
<< metal2 >>
rect 1950 223859 2006 224659
rect 3882 223859 3938 224659
rect 6458 223859 6514 224659
rect 8390 223859 8446 224659
rect 10966 223859 11022 224659
rect 12898 223859 12954 224659
rect 15474 223859 15530 224659
rect 17406 223859 17462 224659
rect 19982 223859 20038 224659
rect 21914 223859 21970 224659
rect 24490 223859 24546 224659
rect 26422 223859 26478 224659
rect 28998 223859 29054 224659
rect 30930 223859 30986 224659
rect 33506 223859 33562 224659
rect 35438 223859 35494 224659
rect 38014 223859 38070 224659
rect 39946 223859 40002 224659
rect 42522 223859 42578 224659
rect 44454 223859 44510 224659
rect 47030 223859 47086 224659
rect 48962 223859 49018 224659
rect 51538 223859 51594 224659
rect 53470 223859 53526 224659
rect 56046 223859 56102 224659
rect 58622 223859 58678 224659
rect 60554 223859 60610 224659
rect 63130 223859 63186 224659
rect 65062 223859 65118 224659
rect 67638 223859 67694 224659
rect 69570 223859 69626 224659
rect 72146 223859 72202 224659
rect 74078 223859 74134 224659
rect 76654 223859 76710 224659
rect 78586 223859 78642 224659
rect 81162 223859 81218 224659
rect 83094 223859 83150 224659
rect 85670 223859 85726 224659
rect 87602 223859 87658 224659
rect 90178 223859 90234 224659
rect 92110 223859 92166 224659
rect 94686 223859 94742 224659
rect 96618 223859 96674 224659
rect 99194 223859 99250 224659
rect 101126 223859 101182 224659
rect 103702 223859 103758 224659
rect 105634 223859 105690 224659
rect 108210 223859 108266 224659
rect 110142 223859 110198 224659
rect 112718 223859 112774 224659
rect 114650 223859 114706 224659
rect 117226 223859 117282 224659
rect 119158 223859 119214 224659
rect 121734 223859 121790 224659
rect 124310 223859 124366 224659
rect 126242 223859 126298 224659
rect 128818 223859 128874 224659
rect 130750 223859 130806 224659
rect 133326 223859 133382 224659
rect 135258 223859 135314 224659
rect 137834 223859 137890 224659
rect 139766 223859 139822 224659
rect 142342 223859 142398 224659
rect 144274 223859 144330 224659
rect 146850 223859 146906 224659
rect 148782 223859 148838 224659
rect 151358 223859 151414 224659
rect 153290 223859 153346 224659
rect 155866 223859 155922 224659
rect 157798 223859 157854 224659
rect 160374 223859 160430 224659
rect 162306 223859 162362 224659
rect 164882 223859 164938 224659
rect 166814 223859 166870 224659
rect 169390 223859 169446 224659
rect 171322 223859 171378 224659
rect 173898 223859 173954 224659
rect 175830 223859 175886 224659
rect 178406 223859 178462 224659
rect 180338 223859 180394 224659
rect 182914 223859 182970 224659
rect 184846 223859 184902 224659
rect 187422 223859 187478 224659
rect 189998 223859 190054 224659
rect 191930 223859 191986 224659
rect 194506 223859 194562 224659
rect 196438 223859 196494 224659
rect 199014 223859 199070 224659
rect 200946 223859 201002 224659
rect 203522 223859 203578 224659
rect 205454 223859 205510 224659
rect 208030 223859 208086 224659
rect 209962 223859 210018 224659
rect 212538 223859 212594 224659
rect 214470 223859 214526 224659
rect 217046 223859 217102 224659
rect 218978 223859 219034 224659
rect 221554 223859 221610 224659
rect 18 0 74 800
rect 1950 0 2006 800
rect 4526 0 4582 800
rect 6458 0 6514 800
rect 9034 0 9090 800
rect 10966 0 11022 800
rect 13542 0 13598 800
rect 15474 0 15530 800
rect 18050 0 18106 800
rect 19982 0 20038 800
rect 22558 0 22614 800
rect 24490 0 24546 800
rect 27066 0 27122 800
rect 28998 0 29054 800
rect 31574 0 31630 800
rect 33506 0 33562 800
rect 36082 0 36138 800
rect 38014 0 38070 800
rect 40590 0 40646 800
rect 42522 0 42578 800
rect 45098 0 45154 800
rect 47030 0 47086 800
rect 49606 0 49662 800
rect 51538 0 51594 800
rect 54114 0 54170 800
rect 56046 0 56102 800
rect 58622 0 58678 800
rect 60554 0 60610 800
rect 63130 0 63186 800
rect 65062 0 65118 800
rect 67638 0 67694 800
rect 70214 0 70270 800
rect 72146 0 72202 800
rect 74722 0 74778 800
rect 76654 0 76710 800
rect 79230 0 79286 800
rect 81162 0 81218 800
rect 83738 0 83794 800
rect 85670 0 85726 800
rect 88246 0 88302 800
rect 90178 0 90234 800
rect 92754 0 92810 800
rect 94686 0 94742 800
rect 97262 0 97318 800
rect 99194 0 99250 800
rect 101770 0 101826 800
rect 103702 0 103758 800
rect 106278 0 106334 800
rect 108210 0 108266 800
rect 110786 0 110842 800
rect 112718 0 112774 800
rect 115294 0 115350 800
rect 117226 0 117282 800
rect 119802 0 119858 800
rect 121734 0 121790 800
rect 124310 0 124366 800
rect 126242 0 126298 800
rect 128818 0 128874 800
rect 130750 0 130806 800
rect 133326 0 133382 800
rect 135902 0 135958 800
rect 137834 0 137890 800
rect 140410 0 140466 800
rect 142342 0 142398 800
rect 144918 0 144974 800
rect 146850 0 146906 800
rect 149426 0 149482 800
rect 151358 0 151414 800
rect 153934 0 153990 800
rect 155866 0 155922 800
rect 158442 0 158498 800
rect 160374 0 160430 800
rect 162950 0 163006 800
rect 164882 0 164938 800
rect 167458 0 167514 800
rect 169390 0 169446 800
rect 171966 0 172022 800
rect 173898 0 173954 800
rect 176474 0 176530 800
rect 178406 0 178462 800
rect 180982 0 181038 800
rect 182914 0 182970 800
rect 185490 0 185546 800
rect 187422 0 187478 800
rect 189998 0 190054 800
rect 191930 0 191986 800
rect 194506 0 194562 800
rect 196438 0 196494 800
rect 199014 0 199070 800
rect 201590 0 201646 800
rect 203522 0 203578 800
rect 206098 0 206154 800
rect 208030 0 208086 800
rect 210606 0 210662 800
rect 212538 0 212594 800
rect 215114 0 215170 800
rect 217046 0 217102 800
rect 219622 0 219678 800
rect 221554 0 221610 800
<< obsm2 >>
rect 1398 223803 1894 223859
rect 2062 223803 3826 223859
rect 3994 223803 6402 223859
rect 6570 223803 8334 223859
rect 8502 223803 10910 223859
rect 11078 223803 12842 223859
rect 13010 223803 15418 223859
rect 15586 223803 17350 223859
rect 17518 223803 19926 223859
rect 20094 223803 21858 223859
rect 22026 223803 24434 223859
rect 24602 223803 26366 223859
rect 26534 223803 28942 223859
rect 29110 223803 30874 223859
rect 31042 223803 33450 223859
rect 33618 223803 35382 223859
rect 35550 223803 37958 223859
rect 38126 223803 39890 223859
rect 40058 223803 42466 223859
rect 42634 223803 44398 223859
rect 44566 223803 46974 223859
rect 47142 223803 48906 223859
rect 49074 223803 51482 223859
rect 51650 223803 53414 223859
rect 53582 223803 55990 223859
rect 56158 223803 58566 223859
rect 58734 223803 60498 223859
rect 60666 223803 63074 223859
rect 63242 223803 65006 223859
rect 65174 223803 67582 223859
rect 67750 223803 69514 223859
rect 69682 223803 72090 223859
rect 72258 223803 74022 223859
rect 74190 223803 76598 223859
rect 76766 223803 78530 223859
rect 78698 223803 81106 223859
rect 81274 223803 83038 223859
rect 83206 223803 85614 223859
rect 85782 223803 87546 223859
rect 87714 223803 90122 223859
rect 90290 223803 92054 223859
rect 92222 223803 94630 223859
rect 94798 223803 96562 223859
rect 96730 223803 99138 223859
rect 99306 223803 101070 223859
rect 101238 223803 103646 223859
rect 103814 223803 105578 223859
rect 105746 223803 108154 223859
rect 108322 223803 110086 223859
rect 110254 223803 112662 223859
rect 112830 223803 114594 223859
rect 114762 223803 117170 223859
rect 117338 223803 119102 223859
rect 119270 223803 121678 223859
rect 121846 223803 124254 223859
rect 124422 223803 126186 223859
rect 126354 223803 128762 223859
rect 128930 223803 130694 223859
rect 130862 223803 133270 223859
rect 133438 223803 135202 223859
rect 135370 223803 137778 223859
rect 137946 223803 139710 223859
rect 139878 223803 142286 223859
rect 142454 223803 144218 223859
rect 144386 223803 146794 223859
rect 146962 223803 148726 223859
rect 148894 223803 151302 223859
rect 151470 223803 153234 223859
rect 153402 223803 155810 223859
rect 155978 223803 157742 223859
rect 157910 223803 160318 223859
rect 160486 223803 162250 223859
rect 162418 223803 164826 223859
rect 164994 223803 166758 223859
rect 166926 223803 169334 223859
rect 169502 223803 171266 223859
rect 171434 223803 173842 223859
rect 174010 223803 175774 223859
rect 175942 223803 178350 223859
rect 178518 223803 180282 223859
rect 180450 223803 182858 223859
rect 183026 223803 184790 223859
rect 184958 223803 187366 223859
rect 187534 223803 189942 223859
rect 190110 223803 191874 223859
rect 192042 223803 194450 223859
rect 194618 223803 196382 223859
rect 196550 223803 198958 223859
rect 199126 223803 200890 223859
rect 201058 223803 203466 223859
rect 203634 223803 205398 223859
rect 205566 223803 207974 223859
rect 208142 223803 209906 223859
rect 210074 223803 212482 223859
rect 212650 223803 214414 223859
rect 214582 223803 216990 223859
rect 217158 223803 218922 223859
rect 219090 223803 220782 223859
rect 1398 856 220782 223803
rect 1398 734 1894 856
rect 2062 734 4470 856
rect 4638 734 6402 856
rect 6570 734 8978 856
rect 9146 734 10910 856
rect 11078 734 13486 856
rect 13654 734 15418 856
rect 15586 734 17994 856
rect 18162 734 19926 856
rect 20094 734 22502 856
rect 22670 734 24434 856
rect 24602 734 27010 856
rect 27178 734 28942 856
rect 29110 734 31518 856
rect 31686 734 33450 856
rect 33618 734 36026 856
rect 36194 734 37958 856
rect 38126 734 40534 856
rect 40702 734 42466 856
rect 42634 734 45042 856
rect 45210 734 46974 856
rect 47142 734 49550 856
rect 49718 734 51482 856
rect 51650 734 54058 856
rect 54226 734 55990 856
rect 56158 734 58566 856
rect 58734 734 60498 856
rect 60666 734 63074 856
rect 63242 734 65006 856
rect 65174 734 67582 856
rect 67750 734 70158 856
rect 70326 734 72090 856
rect 72258 734 74666 856
rect 74834 734 76598 856
rect 76766 734 79174 856
rect 79342 734 81106 856
rect 81274 734 83682 856
rect 83850 734 85614 856
rect 85782 734 88190 856
rect 88358 734 90122 856
rect 90290 734 92698 856
rect 92866 734 94630 856
rect 94798 734 97206 856
rect 97374 734 99138 856
rect 99306 734 101714 856
rect 101882 734 103646 856
rect 103814 734 106222 856
rect 106390 734 108154 856
rect 108322 734 110730 856
rect 110898 734 112662 856
rect 112830 734 115238 856
rect 115406 734 117170 856
rect 117338 734 119746 856
rect 119914 734 121678 856
rect 121846 734 124254 856
rect 124422 734 126186 856
rect 126354 734 128762 856
rect 128930 734 130694 856
rect 130862 734 133270 856
rect 133438 734 135846 856
rect 136014 734 137778 856
rect 137946 734 140354 856
rect 140522 734 142286 856
rect 142454 734 144862 856
rect 145030 734 146794 856
rect 146962 734 149370 856
rect 149538 734 151302 856
rect 151470 734 153878 856
rect 154046 734 155810 856
rect 155978 734 158386 856
rect 158554 734 160318 856
rect 160486 734 162894 856
rect 163062 734 164826 856
rect 164994 734 167402 856
rect 167570 734 169334 856
rect 169502 734 171910 856
rect 172078 734 173842 856
rect 174010 734 176418 856
rect 176586 734 178350 856
rect 178518 734 180926 856
rect 181094 734 182858 856
rect 183026 734 185434 856
rect 185602 734 187366 856
rect 187534 734 189942 856
rect 190110 734 191874 856
rect 192042 734 194450 856
rect 194618 734 196382 856
rect 196550 734 198958 856
rect 199126 734 201534 856
rect 201702 734 203466 856
rect 203634 734 206042 856
rect 206210 734 207974 856
rect 208142 734 210550 856
rect 210718 734 212482 856
rect 212650 734 215058 856
rect 215226 734 216990 856
rect 217158 734 219566 856
rect 219734 734 220782 856
<< metal3 >>
rect 0 224408 800 224528
rect 221715 223728 222515 223848
rect 0 222368 800 222488
rect 221715 221008 222515 221128
rect 0 219648 800 219768
rect 221715 218968 222515 219088
rect 0 217608 800 217728
rect 221715 216248 222515 216368
rect 0 214888 800 215008
rect 221715 214208 222515 214328
rect 0 212848 800 212968
rect 221715 211488 222515 211608
rect 0 210128 800 210248
rect 221715 209448 222515 209568
rect 0 207408 800 207528
rect 221715 206728 222515 206848
rect 0 205368 800 205488
rect 221715 204688 222515 204808
rect 0 202648 800 202768
rect 221715 201968 222515 202088
rect 0 200608 800 200728
rect 221715 199928 222515 200048
rect 0 197888 800 198008
rect 221715 197208 222515 197328
rect 0 195848 800 195968
rect 221715 195168 222515 195288
rect 0 193128 800 193248
rect 221715 192448 222515 192568
rect 0 191088 800 191208
rect 221715 190408 222515 190528
rect 0 188368 800 188488
rect 221715 187688 222515 187808
rect 0 186328 800 186448
rect 221715 184968 222515 185088
rect 0 183608 800 183728
rect 221715 182928 222515 183048
rect 0 181568 800 181688
rect 221715 180208 222515 180328
rect 0 178848 800 178968
rect 221715 178168 222515 178288
rect 0 176808 800 176928
rect 221715 175448 222515 175568
rect 0 174088 800 174208
rect 221715 173408 222515 173528
rect 0 172048 800 172168
rect 221715 170688 222515 170808
rect 0 169328 800 169448
rect 221715 168648 222515 168768
rect 0 167288 800 167408
rect 221715 165928 222515 166048
rect 0 164568 800 164688
rect 221715 163888 222515 164008
rect 0 162528 800 162648
rect 221715 161168 222515 161288
rect 0 159808 800 159928
rect 221715 159128 222515 159248
rect 0 157768 800 157888
rect 221715 156408 222515 156528
rect 0 155048 800 155168
rect 221715 154368 222515 154488
rect 0 153008 800 153128
rect 221715 151648 222515 151768
rect 0 150288 800 150408
rect 221715 149608 222515 149728
rect 0 148248 800 148368
rect 221715 146888 222515 147008
rect 0 145528 800 145648
rect 221715 144848 222515 144968
rect 0 143488 800 143608
rect 221715 142128 222515 142248
rect 0 140768 800 140888
rect 221715 140088 222515 140208
rect 0 138048 800 138168
rect 221715 137368 222515 137488
rect 0 136008 800 136128
rect 221715 135328 222515 135448
rect 0 133288 800 133408
rect 221715 132608 222515 132728
rect 0 131248 800 131368
rect 221715 130568 222515 130688
rect 0 128528 800 128648
rect 221715 127848 222515 127968
rect 0 126488 800 126608
rect 221715 125808 222515 125928
rect 0 123768 800 123888
rect 221715 123088 222515 123208
rect 0 121728 800 121848
rect 221715 121048 222515 121168
rect 0 119008 800 119128
rect 221715 118328 222515 118448
rect 0 116968 800 117088
rect 221715 115608 222515 115728
rect 0 114248 800 114368
rect 221715 113568 222515 113688
rect 0 112208 800 112328
rect 221715 110848 222515 110968
rect 0 109488 800 109608
rect 221715 108808 222515 108928
rect 0 107448 800 107568
rect 221715 106088 222515 106208
rect 0 104728 800 104848
rect 221715 104048 222515 104168
rect 0 102688 800 102808
rect 221715 101328 222515 101448
rect 0 99968 800 100088
rect 221715 99288 222515 99408
rect 0 97928 800 98048
rect 221715 96568 222515 96688
rect 0 95208 800 95328
rect 221715 94528 222515 94648
rect 0 93168 800 93288
rect 221715 91808 222515 91928
rect 0 90448 800 90568
rect 221715 89768 222515 89888
rect 0 88408 800 88528
rect 221715 87048 222515 87168
rect 0 85688 800 85808
rect 221715 85008 222515 85128
rect 0 83648 800 83768
rect 221715 82288 222515 82408
rect 0 80928 800 81048
rect 221715 80248 222515 80368
rect 0 78888 800 79008
rect 221715 77528 222515 77648
rect 0 76168 800 76288
rect 221715 75488 222515 75608
rect 0 74128 800 74248
rect 221715 72768 222515 72888
rect 0 71408 800 71528
rect 221715 70728 222515 70848
rect 0 68688 800 68808
rect 221715 68008 222515 68128
rect 0 66648 800 66768
rect 221715 65968 222515 66088
rect 0 63928 800 64048
rect 221715 63248 222515 63368
rect 0 61888 800 62008
rect 221715 61208 222515 61328
rect 0 59168 800 59288
rect 221715 58488 222515 58608
rect 0 57128 800 57248
rect 221715 56448 222515 56568
rect 0 54408 800 54528
rect 221715 53728 222515 53848
rect 0 52368 800 52488
rect 221715 51688 222515 51808
rect 0 49648 800 49768
rect 221715 48968 222515 49088
rect 0 47608 800 47728
rect 221715 46248 222515 46368
rect 0 44888 800 45008
rect 221715 44208 222515 44328
rect 0 42848 800 42968
rect 221715 41488 222515 41608
rect 0 40128 800 40248
rect 221715 39448 222515 39568
rect 0 38088 800 38208
rect 221715 36728 222515 36848
rect 0 35368 800 35488
rect 221715 34688 222515 34808
rect 0 33328 800 33448
rect 221715 31968 222515 32088
rect 0 30608 800 30728
rect 221715 29928 222515 30048
rect 0 28568 800 28688
rect 221715 27208 222515 27328
rect 0 25848 800 25968
rect 221715 25168 222515 25288
rect 0 23808 800 23928
rect 221715 22448 222515 22568
rect 0 21088 800 21208
rect 221715 20408 222515 20528
rect 0 19048 800 19168
rect 221715 17688 222515 17808
rect 0 16328 800 16448
rect 221715 15648 222515 15768
rect 0 14288 800 14408
rect 221715 12928 222515 13048
rect 0 11568 800 11688
rect 221715 10888 222515 11008
rect 0 9528 800 9648
rect 221715 8168 222515 8288
rect 0 6808 800 6928
rect 221715 6128 222515 6248
rect 0 4768 800 4888
rect 221715 3408 222515 3528
rect 0 2048 800 2168
rect 221715 1368 222515 1488
<< obsm3 >>
rect 800 223648 221635 223821
rect 800 222568 221715 223648
rect 880 222288 221715 222568
rect 800 221208 221715 222288
rect 800 220928 221635 221208
rect 800 219848 221715 220928
rect 880 219568 221715 219848
rect 800 219168 221715 219568
rect 800 218888 221635 219168
rect 800 217808 221715 218888
rect 880 217528 221715 217808
rect 800 216448 221715 217528
rect 800 216168 221635 216448
rect 800 215088 221715 216168
rect 880 214808 221715 215088
rect 800 214408 221715 214808
rect 800 214128 221635 214408
rect 800 213048 221715 214128
rect 880 212768 221715 213048
rect 800 211688 221715 212768
rect 800 211408 221635 211688
rect 800 210328 221715 211408
rect 880 210048 221715 210328
rect 800 209648 221715 210048
rect 800 209368 221635 209648
rect 800 207608 221715 209368
rect 880 207328 221715 207608
rect 800 206928 221715 207328
rect 800 206648 221635 206928
rect 800 205568 221715 206648
rect 880 205288 221715 205568
rect 800 204888 221715 205288
rect 800 204608 221635 204888
rect 800 202848 221715 204608
rect 880 202568 221715 202848
rect 800 202168 221715 202568
rect 800 201888 221635 202168
rect 800 200808 221715 201888
rect 880 200528 221715 200808
rect 800 200128 221715 200528
rect 800 199848 221635 200128
rect 800 198088 221715 199848
rect 880 197808 221715 198088
rect 800 197408 221715 197808
rect 800 197128 221635 197408
rect 800 196048 221715 197128
rect 880 195768 221715 196048
rect 800 195368 221715 195768
rect 800 195088 221635 195368
rect 800 193328 221715 195088
rect 880 193048 221715 193328
rect 800 192648 221715 193048
rect 800 192368 221635 192648
rect 800 191288 221715 192368
rect 880 191008 221715 191288
rect 800 190608 221715 191008
rect 800 190328 221635 190608
rect 800 188568 221715 190328
rect 880 188288 221715 188568
rect 800 187888 221715 188288
rect 800 187608 221635 187888
rect 800 186528 221715 187608
rect 880 186248 221715 186528
rect 800 185168 221715 186248
rect 800 184888 221635 185168
rect 800 183808 221715 184888
rect 880 183528 221715 183808
rect 800 183128 221715 183528
rect 800 182848 221635 183128
rect 800 181768 221715 182848
rect 880 181488 221715 181768
rect 800 180408 221715 181488
rect 800 180128 221635 180408
rect 800 179048 221715 180128
rect 880 178768 221715 179048
rect 800 178368 221715 178768
rect 800 178088 221635 178368
rect 800 177008 221715 178088
rect 880 176728 221715 177008
rect 800 175648 221715 176728
rect 800 175368 221635 175648
rect 800 174288 221715 175368
rect 880 174008 221715 174288
rect 800 173608 221715 174008
rect 800 173328 221635 173608
rect 800 172248 221715 173328
rect 880 171968 221715 172248
rect 800 170888 221715 171968
rect 800 170608 221635 170888
rect 800 169528 221715 170608
rect 880 169248 221715 169528
rect 800 168848 221715 169248
rect 800 168568 221635 168848
rect 800 167488 221715 168568
rect 880 167208 221715 167488
rect 800 166128 221715 167208
rect 800 165848 221635 166128
rect 800 164768 221715 165848
rect 880 164488 221715 164768
rect 800 164088 221715 164488
rect 800 163808 221635 164088
rect 800 162728 221715 163808
rect 880 162448 221715 162728
rect 800 161368 221715 162448
rect 800 161088 221635 161368
rect 800 160008 221715 161088
rect 880 159728 221715 160008
rect 800 159328 221715 159728
rect 800 159048 221635 159328
rect 800 157968 221715 159048
rect 880 157688 221715 157968
rect 800 156608 221715 157688
rect 800 156328 221635 156608
rect 800 155248 221715 156328
rect 880 154968 221715 155248
rect 800 154568 221715 154968
rect 800 154288 221635 154568
rect 800 153208 221715 154288
rect 880 152928 221715 153208
rect 800 151848 221715 152928
rect 800 151568 221635 151848
rect 800 150488 221715 151568
rect 880 150208 221715 150488
rect 800 149808 221715 150208
rect 800 149528 221635 149808
rect 800 148448 221715 149528
rect 880 148168 221715 148448
rect 800 147088 221715 148168
rect 800 146808 221635 147088
rect 800 145728 221715 146808
rect 880 145448 221715 145728
rect 800 145048 221715 145448
rect 800 144768 221635 145048
rect 800 143688 221715 144768
rect 880 143408 221715 143688
rect 800 142328 221715 143408
rect 800 142048 221635 142328
rect 800 140968 221715 142048
rect 880 140688 221715 140968
rect 800 140288 221715 140688
rect 800 140008 221635 140288
rect 800 138248 221715 140008
rect 880 137968 221715 138248
rect 800 137568 221715 137968
rect 800 137288 221635 137568
rect 800 136208 221715 137288
rect 880 135928 221715 136208
rect 800 135528 221715 135928
rect 800 135248 221635 135528
rect 800 133488 221715 135248
rect 880 133208 221715 133488
rect 800 132808 221715 133208
rect 800 132528 221635 132808
rect 800 131448 221715 132528
rect 880 131168 221715 131448
rect 800 130768 221715 131168
rect 800 130488 221635 130768
rect 800 128728 221715 130488
rect 880 128448 221715 128728
rect 800 128048 221715 128448
rect 800 127768 221635 128048
rect 800 126688 221715 127768
rect 880 126408 221715 126688
rect 800 126008 221715 126408
rect 800 125728 221635 126008
rect 800 123968 221715 125728
rect 880 123688 221715 123968
rect 800 123288 221715 123688
rect 800 123008 221635 123288
rect 800 121928 221715 123008
rect 880 121648 221715 121928
rect 800 121248 221715 121648
rect 800 120968 221635 121248
rect 800 119208 221715 120968
rect 880 118928 221715 119208
rect 800 118528 221715 118928
rect 800 118248 221635 118528
rect 800 117168 221715 118248
rect 880 116888 221715 117168
rect 800 115808 221715 116888
rect 800 115528 221635 115808
rect 800 114448 221715 115528
rect 880 114168 221715 114448
rect 800 113768 221715 114168
rect 800 113488 221635 113768
rect 800 112408 221715 113488
rect 880 112128 221715 112408
rect 800 111048 221715 112128
rect 800 110768 221635 111048
rect 800 109688 221715 110768
rect 880 109408 221715 109688
rect 800 109008 221715 109408
rect 800 108728 221635 109008
rect 800 107648 221715 108728
rect 880 107368 221715 107648
rect 800 106288 221715 107368
rect 800 106008 221635 106288
rect 800 104928 221715 106008
rect 880 104648 221715 104928
rect 800 104248 221715 104648
rect 800 103968 221635 104248
rect 800 102888 221715 103968
rect 880 102608 221715 102888
rect 800 101528 221715 102608
rect 800 101248 221635 101528
rect 800 100168 221715 101248
rect 880 99888 221715 100168
rect 800 99488 221715 99888
rect 800 99208 221635 99488
rect 800 98128 221715 99208
rect 880 97848 221715 98128
rect 800 96768 221715 97848
rect 800 96488 221635 96768
rect 800 95408 221715 96488
rect 880 95128 221715 95408
rect 800 94728 221715 95128
rect 800 94448 221635 94728
rect 800 93368 221715 94448
rect 880 93088 221715 93368
rect 800 92008 221715 93088
rect 800 91728 221635 92008
rect 800 90648 221715 91728
rect 880 90368 221715 90648
rect 800 89968 221715 90368
rect 800 89688 221635 89968
rect 800 88608 221715 89688
rect 880 88328 221715 88608
rect 800 87248 221715 88328
rect 800 86968 221635 87248
rect 800 85888 221715 86968
rect 880 85608 221715 85888
rect 800 85208 221715 85608
rect 800 84928 221635 85208
rect 800 83848 221715 84928
rect 880 83568 221715 83848
rect 800 82488 221715 83568
rect 800 82208 221635 82488
rect 800 81128 221715 82208
rect 880 80848 221715 81128
rect 800 80448 221715 80848
rect 800 80168 221635 80448
rect 800 79088 221715 80168
rect 880 78808 221715 79088
rect 800 77728 221715 78808
rect 800 77448 221635 77728
rect 800 76368 221715 77448
rect 880 76088 221715 76368
rect 800 75688 221715 76088
rect 800 75408 221635 75688
rect 800 74328 221715 75408
rect 880 74048 221715 74328
rect 800 72968 221715 74048
rect 800 72688 221635 72968
rect 800 71608 221715 72688
rect 880 71328 221715 71608
rect 800 70928 221715 71328
rect 800 70648 221635 70928
rect 800 68888 221715 70648
rect 880 68608 221715 68888
rect 800 68208 221715 68608
rect 800 67928 221635 68208
rect 800 66848 221715 67928
rect 880 66568 221715 66848
rect 800 66168 221715 66568
rect 800 65888 221635 66168
rect 800 64128 221715 65888
rect 880 63848 221715 64128
rect 800 63448 221715 63848
rect 800 63168 221635 63448
rect 800 62088 221715 63168
rect 880 61808 221715 62088
rect 800 61408 221715 61808
rect 800 61128 221635 61408
rect 800 59368 221715 61128
rect 880 59088 221715 59368
rect 800 58688 221715 59088
rect 800 58408 221635 58688
rect 800 57328 221715 58408
rect 880 57048 221715 57328
rect 800 56648 221715 57048
rect 800 56368 221635 56648
rect 800 54608 221715 56368
rect 880 54328 221715 54608
rect 800 53928 221715 54328
rect 800 53648 221635 53928
rect 800 52568 221715 53648
rect 880 52288 221715 52568
rect 800 51888 221715 52288
rect 800 51608 221635 51888
rect 800 49848 221715 51608
rect 880 49568 221715 49848
rect 800 49168 221715 49568
rect 800 48888 221635 49168
rect 800 47808 221715 48888
rect 880 47528 221715 47808
rect 800 46448 221715 47528
rect 800 46168 221635 46448
rect 800 45088 221715 46168
rect 880 44808 221715 45088
rect 800 44408 221715 44808
rect 800 44128 221635 44408
rect 800 43048 221715 44128
rect 880 42768 221715 43048
rect 800 41688 221715 42768
rect 800 41408 221635 41688
rect 800 40328 221715 41408
rect 880 40048 221715 40328
rect 800 39648 221715 40048
rect 800 39368 221635 39648
rect 800 38288 221715 39368
rect 880 38008 221715 38288
rect 800 36928 221715 38008
rect 800 36648 221635 36928
rect 800 35568 221715 36648
rect 880 35288 221715 35568
rect 800 34888 221715 35288
rect 800 34608 221635 34888
rect 800 33528 221715 34608
rect 880 33248 221715 33528
rect 800 32168 221715 33248
rect 800 31888 221635 32168
rect 800 30808 221715 31888
rect 880 30528 221715 30808
rect 800 30128 221715 30528
rect 800 29848 221635 30128
rect 800 28768 221715 29848
rect 880 28488 221715 28768
rect 800 27408 221715 28488
rect 800 27128 221635 27408
rect 800 26048 221715 27128
rect 880 25768 221715 26048
rect 800 25368 221715 25768
rect 800 25088 221635 25368
rect 800 24008 221715 25088
rect 880 23728 221715 24008
rect 800 22648 221715 23728
rect 800 22368 221635 22648
rect 800 21288 221715 22368
rect 880 21008 221715 21288
rect 800 20608 221715 21008
rect 800 20328 221635 20608
rect 800 19248 221715 20328
rect 880 18968 221715 19248
rect 800 17888 221715 18968
rect 800 17608 221635 17888
rect 800 16528 221715 17608
rect 880 16248 221715 16528
rect 800 15848 221715 16248
rect 800 15568 221635 15848
rect 800 14488 221715 15568
rect 880 14208 221715 14488
rect 800 13128 221715 14208
rect 800 12848 221635 13128
rect 800 11768 221715 12848
rect 880 11488 221715 11768
rect 800 11088 221715 11488
rect 800 10808 221635 11088
rect 800 9728 221715 10808
rect 880 9448 221715 9728
rect 800 8368 221715 9448
rect 800 8088 221635 8368
rect 800 7008 221715 8088
rect 880 6728 221715 7008
rect 800 6328 221715 6728
rect 800 6048 221635 6328
rect 800 4968 221715 6048
rect 880 4688 221715 4968
rect 800 3608 221715 4688
rect 800 3328 221635 3608
rect 800 2248 221715 3328
rect 880 2075 221715 2248
<< metal4 >>
rect 4208 2128 4528 222000
rect 19568 2128 19888 222000
rect 34928 2128 35248 222000
rect 50288 2128 50608 222000
rect 65648 2128 65968 222000
rect 81008 2128 81328 222000
rect 96368 2128 96688 222000
rect 111728 2128 112048 222000
rect 127088 2128 127408 222000
rect 142448 2128 142768 222000
rect 157808 2128 158128 222000
rect 173168 2128 173488 222000
rect 188528 2128 188848 222000
rect 203888 2128 204208 222000
rect 219248 2128 219568 222000
<< obsm4 >>
rect 27659 2347 34848 221509
rect 35328 2347 50208 221509
rect 50688 2347 65568 221509
rect 66048 2347 80928 221509
rect 81408 2347 96288 221509
rect 96768 2347 111648 221509
rect 112128 2347 127008 221509
rect 127488 2347 142368 221509
rect 142848 2347 157728 221509
rect 158208 2347 160205 221509
<< labels >>
rlabel metal3 s 0 95208 800 95328 6 clk
port 1 nsew signal input
rlabel metal2 s 208030 223859 208086 224659 6 la_data_in[0]
port 2 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 la_data_in[100]
port 3 nsew signal input
rlabel metal2 s 182914 223859 182970 224659 6 la_data_in[101]
port 4 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 la_data_in[102]
port 5 nsew signal input
rlabel metal3 s 0 138048 800 138168 6 la_data_in[103]
port 6 nsew signal input
rlabel metal3 s 0 126488 800 126608 6 la_data_in[104]
port 7 nsew signal input
rlabel metal3 s 221715 36728 222515 36848 6 la_data_in[105]
port 8 nsew signal input
rlabel metal3 s 0 200608 800 200728 6 la_data_in[106]
port 9 nsew signal input
rlabel metal2 s 92110 223859 92166 224659 6 la_data_in[107]
port 10 nsew signal input
rlabel metal2 s 78586 223859 78642 224659 6 la_data_in[108]
port 11 nsew signal input
rlabel metal2 s 153290 223859 153346 224659 6 la_data_in[109]
port 12 nsew signal input
rlabel metal3 s 221715 46248 222515 46368 6 la_data_in[10]
port 13 nsew signal input
rlabel metal2 s 199014 223859 199070 224659 6 la_data_in[110]
port 14 nsew signal input
rlabel metal3 s 0 148248 800 148368 6 la_data_in[111]
port 15 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 la_data_in[112]
port 16 nsew signal input
rlabel metal3 s 221715 68008 222515 68128 6 la_data_in[113]
port 17 nsew signal input
rlabel metal2 s 214470 223859 214526 224659 6 la_data_in[114]
port 18 nsew signal input
rlabel metal3 s 0 183608 800 183728 6 la_data_in[115]
port 19 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 la_data_in[116]
port 20 nsew signal input
rlabel metal3 s 221715 211488 222515 211608 6 la_data_in[117]
port 21 nsew signal input
rlabel metal3 s 221715 132608 222515 132728 6 la_data_in[118]
port 22 nsew signal input
rlabel metal2 s 196438 0 196494 800 6 la_data_in[119]
port 23 nsew signal input
rlabel metal2 s 173898 223859 173954 224659 6 la_data_in[11]
port 24 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 la_data_in[120]
port 25 nsew signal input
rlabel metal3 s 0 224408 800 224528 6 la_data_in[121]
port 26 nsew signal input
rlabel metal2 s 87602 223859 87658 224659 6 la_data_in[122]
port 27 nsew signal input
rlabel metal3 s 221715 190408 222515 190528 6 la_data_in[123]
port 28 nsew signal input
rlabel metal3 s 221715 77528 222515 77648 6 la_data_in[124]
port 29 nsew signal input
rlabel metal3 s 0 219648 800 219768 6 la_data_in[125]
port 30 nsew signal input
rlabel metal2 s 166814 223859 166870 224659 6 la_data_in[126]
port 31 nsew signal input
rlabel metal3 s 221715 161168 222515 161288 6 la_data_in[127]
port 32 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 la_data_in[12]
port 33 nsew signal input
rlabel metal3 s 221715 115608 222515 115728 6 la_data_in[13]
port 34 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 la_data_in[14]
port 35 nsew signal input
rlabel metal2 s 212538 0 212594 800 6 la_data_in[15]
port 36 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 la_data_in[16]
port 37 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 la_data_in[17]
port 38 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 la_data_in[18]
port 39 nsew signal input
rlabel metal3 s 221715 48968 222515 49088 6 la_data_in[19]
port 40 nsew signal input
rlabel metal3 s 221715 209448 222515 209568 6 la_data_in[1]
port 41 nsew signal input
rlabel metal2 s 191930 0 191986 800 6 la_data_in[20]
port 42 nsew signal input
rlabel metal3 s 221715 149608 222515 149728 6 la_data_in[21]
port 43 nsew signal input
rlabel metal3 s 221715 223728 222515 223848 6 la_data_in[22]
port 44 nsew signal input
rlabel metal2 s 142342 0 142398 800 6 la_data_in[23]
port 45 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 la_data_in[24]
port 46 nsew signal input
rlabel metal2 s 58622 223859 58678 224659 6 la_data_in[25]
port 47 nsew signal input
rlabel metal2 s 53470 223859 53526 224659 6 la_data_in[26]
port 48 nsew signal input
rlabel metal2 s 114650 223859 114706 224659 6 la_data_in[27]
port 49 nsew signal input
rlabel metal3 s 0 172048 800 172168 6 la_data_in[28]
port 50 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 la_data_in[29]
port 51 nsew signal input
rlabel metal3 s 221715 178168 222515 178288 6 la_data_in[2]
port 52 nsew signal input
rlabel metal3 s 221715 106088 222515 106208 6 la_data_in[30]
port 53 nsew signal input
rlabel metal2 s 12898 223859 12954 224659 6 la_data_in[31]
port 54 nsew signal input
rlabel metal2 s 203522 0 203578 800 6 la_data_in[32]
port 55 nsew signal input
rlabel metal3 s 221715 25168 222515 25288 6 la_data_in[33]
port 56 nsew signal input
rlabel metal3 s 221715 137368 222515 137488 6 la_data_in[34]
port 57 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 la_data_in[35]
port 58 nsew signal input
rlabel metal3 s 221715 221008 222515 221128 6 la_data_in[36]
port 59 nsew signal input
rlabel metal3 s 221715 96568 222515 96688 6 la_data_in[37]
port 60 nsew signal input
rlabel metal3 s 221715 199928 222515 200048 6 la_data_in[38]
port 61 nsew signal input
rlabel metal3 s 0 167288 800 167408 6 la_data_in[39]
port 62 nsew signal input
rlabel metal2 s 144274 223859 144330 224659 6 la_data_in[3]
port 63 nsew signal input
rlabel metal3 s 0 178848 800 178968 6 la_data_in[40]
port 64 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 la_data_in[41]
port 65 nsew signal input
rlabel metal2 s 187422 0 187478 800 6 la_data_in[42]
port 66 nsew signal input
rlabel metal2 s 110142 223859 110198 224659 6 la_data_in[43]
port 67 nsew signal input
rlabel metal2 s 153934 0 153990 800 6 la_data_in[44]
port 68 nsew signal input
rlabel metal2 s 178406 223859 178462 224659 6 la_data_in[45]
port 69 nsew signal input
rlabel metal2 s 210606 0 210662 800 6 la_data_in[46]
port 70 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 la_data_in[47]
port 71 nsew signal input
rlabel metal2 s 130750 223859 130806 224659 6 la_data_in[48]
port 72 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 la_data_in[49]
port 73 nsew signal input
rlabel metal3 s 221715 180208 222515 180328 6 la_data_in[4]
port 74 nsew signal input
rlabel metal2 s 96618 223859 96674 224659 6 la_data_in[50]
port 75 nsew signal input
rlabel metal3 s 221715 113568 222515 113688 6 la_data_in[51]
port 76 nsew signal input
rlabel metal2 s 169390 0 169446 800 6 la_data_in[52]
port 77 nsew signal input
rlabel metal3 s 221715 168648 222515 168768 6 la_data_in[53]
port 78 nsew signal input
rlabel metal3 s 221715 165928 222515 166048 6 la_data_in[54]
port 79 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 la_data_in[55]
port 80 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 la_data_in[56]
port 81 nsew signal input
rlabel metal3 s 0 150288 800 150408 6 la_data_in[57]
port 82 nsew signal input
rlabel metal3 s 221715 39448 222515 39568 6 la_data_in[58]
port 83 nsew signal input
rlabel metal2 s 47030 223859 47086 224659 6 la_data_in[59]
port 84 nsew signal input
rlabel metal2 s 173898 0 173954 800 6 la_data_in[5]
port 85 nsew signal input
rlabel metal2 s 221554 0 221610 800 6 la_data_in[60]
port 86 nsew signal input
rlabel metal2 s 8390 223859 8446 224659 6 la_data_in[61]
port 87 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 la_data_in[62]
port 88 nsew signal input
rlabel metal3 s 221715 214208 222515 214328 6 la_data_in[63]
port 89 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_data_in[64]
port 90 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_data_in[65]
port 91 nsew signal input
rlabel metal2 s 39946 223859 40002 224659 6 la_data_in[66]
port 92 nsew signal input
rlabel metal3 s 221715 195168 222515 195288 6 la_data_in[67]
port 93 nsew signal input
rlabel metal2 s 60554 223859 60610 224659 6 la_data_in[68]
port 94 nsew signal input
rlabel metal2 s 17406 223859 17462 224659 6 la_data_in[69]
port 95 nsew signal input
rlabel metal3 s 0 174088 800 174208 6 la_data_in[6]
port 96 nsew signal input
rlabel metal2 s 35438 223859 35494 224659 6 la_data_in[70]
port 97 nsew signal input
rlabel metal3 s 221715 51688 222515 51808 6 la_data_in[71]
port 98 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_data_in[72]
port 99 nsew signal input
rlabel metal2 s 103702 223859 103758 224659 6 la_data_in[73]
port 100 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 la_data_in[74]
port 101 nsew signal input
rlabel metal2 s 112718 223859 112774 224659 6 la_data_in[75]
port 102 nsew signal input
rlabel metal3 s 221715 17688 222515 17808 6 la_data_in[76]
port 103 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_data_in[77]
port 104 nsew signal input
rlabel metal2 s 133326 223859 133382 224659 6 la_data_in[78]
port 105 nsew signal input
rlabel metal3 s 221715 151648 222515 151768 6 la_data_in[79]
port 106 nsew signal input
rlabel metal3 s 221715 10888 222515 11008 6 la_data_in[7]
port 107 nsew signal input
rlabel metal2 s 221554 223859 221610 224659 6 la_data_in[80]
port 108 nsew signal input
rlabel metal3 s 0 131248 800 131368 6 la_data_in[81]
port 109 nsew signal input
rlabel metal2 s 135258 223859 135314 224659 6 la_data_in[82]
port 110 nsew signal input
rlabel metal2 s 194506 223859 194562 224659 6 la_data_in[83]
port 111 nsew signal input
rlabel metal3 s 221715 184968 222515 185088 6 la_data_in[84]
port 112 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 la_data_in[85]
port 113 nsew signal input
rlabel metal3 s 221715 182928 222515 183048 6 la_data_in[86]
port 114 nsew signal input
rlabel metal3 s 0 99968 800 100088 6 la_data_in[87]
port 115 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 la_data_in[88]
port 116 nsew signal input
rlabel metal2 s 26422 223859 26478 224659 6 la_data_in[89]
port 117 nsew signal input
rlabel metal3 s 0 159808 800 159928 6 la_data_in[8]
port 118 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 la_data_in[90]
port 119 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 la_data_in[91]
port 120 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 la_data_in[92]
port 121 nsew signal input
rlabel metal2 s 189998 0 190054 800 6 la_data_in[93]
port 122 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_data_in[94]
port 123 nsew signal input
rlabel metal2 s 3882 223859 3938 224659 6 la_data_in[95]
port 124 nsew signal input
rlabel metal3 s 0 162528 800 162648 6 la_data_in[96]
port 125 nsew signal input
rlabel metal2 s 69570 223859 69626 224659 6 la_data_in[97]
port 126 nsew signal input
rlabel metal3 s 0 68688 800 68808 6 la_data_in[98]
port 127 nsew signal input
rlabel metal2 s 105634 223859 105690 224659 6 la_data_in[99]
port 128 nsew signal input
rlabel metal3 s 221715 82288 222515 82408 6 la_data_in[9]
port 129 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_data_out[0]
port 130 nsew signal output
rlabel metal3 s 221715 31968 222515 32088 6 la_data_out[100]
port 131 nsew signal output
rlabel metal2 s 6458 223859 6514 224659 6 la_data_out[101]
port 132 nsew signal output
rlabel metal3 s 221715 22448 222515 22568 6 la_data_out[102]
port 133 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 la_data_out[103]
port 134 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 la_data_out[104]
port 135 nsew signal output
rlabel metal2 s 199014 0 199070 800 6 la_data_out[105]
port 136 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 la_data_out[106]
port 137 nsew signal output
rlabel metal2 s 187422 223859 187478 224659 6 la_data_out[107]
port 138 nsew signal output
rlabel metal3 s 0 140768 800 140888 6 la_data_out[108]
port 139 nsew signal output
rlabel metal2 s 21914 223859 21970 224659 6 la_data_out[109]
port 140 nsew signal output
rlabel metal2 s 99194 0 99250 800 6 la_data_out[10]
port 141 nsew signal output
rlabel metal3 s 0 217608 800 217728 6 la_data_out[110]
port 142 nsew signal output
rlabel metal2 s 126242 223859 126298 224659 6 la_data_out[111]
port 143 nsew signal output
rlabel metal2 s 137834 223859 137890 224659 6 la_data_out[112]
port 144 nsew signal output
rlabel metal3 s 221715 44208 222515 44328 6 la_data_out[113]
port 145 nsew signal output
rlabel metal3 s 221715 201968 222515 202088 6 la_data_out[114]
port 146 nsew signal output
rlabel metal2 s 178406 0 178462 800 6 la_data_out[115]
port 147 nsew signal output
rlabel metal3 s 221715 75488 222515 75608 6 la_data_out[116]
port 148 nsew signal output
rlabel metal3 s 221715 80248 222515 80368 6 la_data_out[117]
port 149 nsew signal output
rlabel metal2 s 140410 0 140466 800 6 la_data_out[118]
port 150 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 la_data_out[119]
port 151 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 la_data_out[11]
port 152 nsew signal output
rlabel metal3 s 221715 56448 222515 56568 6 la_data_out[120]
port 153 nsew signal output
rlabel metal3 s 221715 175448 222515 175568 6 la_data_out[121]
port 154 nsew signal output
rlabel metal3 s 0 164568 800 164688 6 la_data_out[122]
port 155 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 la_data_out[123]
port 156 nsew signal output
rlabel metal3 s 221715 144848 222515 144968 6 la_data_out[124]
port 157 nsew signal output
rlabel metal3 s 0 143488 800 143608 6 la_data_out[125]
port 158 nsew signal output
rlabel metal3 s 221715 70728 222515 70848 6 la_data_out[126]
port 159 nsew signal output
rlabel metal2 s 15474 223859 15530 224659 6 la_data_out[127]
port 160 nsew signal output
rlabel metal3 s 221715 121048 222515 121168 6 la_data_out[12]
port 161 nsew signal output
rlabel metal2 s 139766 223859 139822 224659 6 la_data_out[13]
port 162 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 la_data_out[14]
port 163 nsew signal output
rlabel metal3 s 221715 34688 222515 34808 6 la_data_out[15]
port 164 nsew signal output
rlabel metal2 s 121734 223859 121790 224659 6 la_data_out[16]
port 165 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 la_data_out[17]
port 166 nsew signal output
rlabel metal2 s 51538 223859 51594 224659 6 la_data_out[18]
port 167 nsew signal output
rlabel metal3 s 221715 142128 222515 142248 6 la_data_out[19]
port 168 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 la_data_out[1]
port 169 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 la_data_out[20]
port 170 nsew signal output
rlabel metal3 s 221715 72768 222515 72888 6 la_data_out[21]
port 171 nsew signal output
rlabel metal2 s 74078 223859 74134 224659 6 la_data_out[22]
port 172 nsew signal output
rlabel metal2 s 38014 223859 38070 224659 6 la_data_out[23]
port 173 nsew signal output
rlabel metal3 s 221715 15648 222515 15768 6 la_data_out[24]
port 174 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 la_data_out[25]
port 175 nsew signal output
rlabel metal2 s 196438 223859 196494 224659 6 la_data_out[26]
port 176 nsew signal output
rlabel metal3 s 221715 146888 222515 147008 6 la_data_out[27]
port 177 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 la_data_out[28]
port 178 nsew signal output
rlabel metal3 s 0 222368 800 222488 6 la_data_out[29]
port 179 nsew signal output
rlabel metal3 s 0 93168 800 93288 6 la_data_out[2]
port 180 nsew signal output
rlabel metal2 s 126242 0 126298 800 6 la_data_out[30]
port 181 nsew signal output
rlabel metal2 s 56046 223859 56102 224659 6 la_data_out[31]
port 182 nsew signal output
rlabel metal2 s 189998 223859 190054 224659 6 la_data_out[32]
port 183 nsew signal output
rlabel metal3 s 221715 156408 222515 156528 6 la_data_out[33]
port 184 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 la_data_out[34]
port 185 nsew signal output
rlabel metal3 s 0 193128 800 193248 6 la_data_out[35]
port 186 nsew signal output
rlabel metal2 s 19982 223859 20038 224659 6 la_data_out[36]
port 187 nsew signal output
rlabel metal2 s 142342 223859 142398 224659 6 la_data_out[37]
port 188 nsew signal output
rlabel metal3 s 0 176808 800 176928 6 la_data_out[38]
port 189 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 la_data_out[39]
port 190 nsew signal output
rlabel metal2 s 182914 0 182970 800 6 la_data_out[3]
port 191 nsew signal output
rlabel metal3 s 221715 89768 222515 89888 6 la_data_out[40]
port 192 nsew signal output
rlabel metal3 s 221715 3408 222515 3528 6 la_data_out[41]
port 193 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 la_data_out[42]
port 194 nsew signal output
rlabel metal2 s 101126 223859 101182 224659 6 la_data_out[43]
port 195 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 la_data_out[44]
port 196 nsew signal output
rlabel metal2 s 1950 223859 2006 224659 6 la_data_out[45]
port 197 nsew signal output
rlabel metal2 s 103702 0 103758 800 6 la_data_out[46]
port 198 nsew signal output
rlabel metal3 s 221715 29928 222515 30048 6 la_data_out[47]
port 199 nsew signal output
rlabel metal2 s 200946 223859 201002 224659 6 la_data_out[48]
port 200 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 la_data_out[49]
port 201 nsew signal output
rlabel metal2 s 128818 223859 128874 224659 6 la_data_out[4]
port 202 nsew signal output
rlabel metal3 s 0 80928 800 81048 6 la_data_out[50]
port 203 nsew signal output
rlabel metal2 s 209962 223859 210018 224659 6 la_data_out[51]
port 204 nsew signal output
rlabel metal2 s 42522 223859 42578 224659 6 la_data_out[52]
port 205 nsew signal output
rlabel metal3 s 0 61888 800 62008 6 la_data_out[53]
port 206 nsew signal output
rlabel metal2 s 219622 0 219678 800 6 la_data_out[54]
port 207 nsew signal output
rlabel metal3 s 0 210128 800 210248 6 la_data_out[55]
port 208 nsew signal output
rlabel metal3 s 0 195848 800 195968 6 la_data_out[56]
port 209 nsew signal output
rlabel metal2 s 128818 0 128874 800 6 la_data_out[57]
port 210 nsew signal output
rlabel metal3 s 221715 85008 222515 85128 6 la_data_out[58]
port 211 nsew signal output
rlabel metal3 s 221715 63248 222515 63368 6 la_data_out[59]
port 212 nsew signal output
rlabel metal2 s 81162 223859 81218 224659 6 la_data_out[5]
port 213 nsew signal output
rlabel metal3 s 221715 104048 222515 104168 6 la_data_out[60]
port 214 nsew signal output
rlabel metal2 s 155866 0 155922 800 6 la_data_out[61]
port 215 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 la_data_out[62]
port 216 nsew signal output
rlabel metal2 s 151358 0 151414 800 6 la_data_out[63]
port 217 nsew signal output
rlabel metal2 s 180982 0 181038 800 6 la_data_out[64]
port 218 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 la_data_out[65]
port 219 nsew signal output
rlabel metal3 s 0 155048 800 155168 6 la_data_out[66]
port 220 nsew signal output
rlabel metal2 s 164882 0 164938 800 6 la_data_out[67]
port 221 nsew signal output
rlabel metal3 s 0 107448 800 107568 6 la_data_out[68]
port 222 nsew signal output
rlabel metal3 s 0 169328 800 169448 6 la_data_out[69]
port 223 nsew signal output
rlabel metal3 s 221715 218968 222515 219088 6 la_data_out[6]
port 224 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 la_data_out[70]
port 225 nsew signal output
rlabel metal3 s 0 123768 800 123888 6 la_data_out[71]
port 226 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 la_data_out[72]
port 227 nsew signal output
rlabel metal3 s 221715 118328 222515 118448 6 la_data_out[73]
port 228 nsew signal output
rlabel metal2 s 185490 0 185546 800 6 la_data_out[74]
port 229 nsew signal output
rlabel metal2 s 175830 223859 175886 224659 6 la_data_out[75]
port 230 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 la_data_out[76]
port 231 nsew signal output
rlabel metal2 s 48962 223859 49018 224659 6 la_data_out[77]
port 232 nsew signal output
rlabel metal3 s 221715 192448 222515 192568 6 la_data_out[78]
port 233 nsew signal output
rlabel metal3 s 0 83648 800 83768 6 la_data_out[79]
port 234 nsew signal output
rlabel metal3 s 221715 173408 222515 173528 6 la_data_out[7]
port 235 nsew signal output
rlabel metal2 s 124310 223859 124366 224659 6 la_data_out[80]
port 236 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 la_data_out[81]
port 237 nsew signal output
rlabel metal3 s 0 102688 800 102808 6 la_data_out[82]
port 238 nsew signal output
rlabel metal3 s 0 136008 800 136128 6 la_data_out[83]
port 239 nsew signal output
rlabel metal2 s 99194 223859 99250 224659 6 la_data_out[84]
port 240 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 la_data_out[85]
port 241 nsew signal output
rlabel metal2 s 65062 223859 65118 224659 6 la_data_out[86]
port 242 nsew signal output
rlabel metal2 s 108210 0 108266 800 6 la_data_out[87]
port 243 nsew signal output
rlabel metal2 s 217046 0 217102 800 6 la_data_out[88]
port 244 nsew signal output
rlabel metal3 s 221715 216248 222515 216368 6 la_data_out[89]
port 245 nsew signal output
rlabel metal3 s 221715 12928 222515 13048 6 la_data_out[8]
port 246 nsew signal output
rlabel metal2 s 108210 223859 108266 224659 6 la_data_out[90]
port 247 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 la_data_out[91]
port 248 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 la_data_out[92]
port 249 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 la_data_out[93]
port 250 nsew signal output
rlabel metal2 s 203522 223859 203578 224659 6 la_data_out[94]
port 251 nsew signal output
rlabel metal3 s 0 186328 800 186448 6 la_data_out[95]
port 252 nsew signal output
rlabel metal2 s 79230 0 79286 800 6 la_data_out[96]
port 253 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 la_data_out[97]
port 254 nsew signal output
rlabel metal3 s 221715 94528 222515 94648 6 la_data_out[98]
port 255 nsew signal output
rlabel metal3 s 0 207408 800 207528 6 la_data_out[99]
port 256 nsew signal output
rlabel metal2 s 162950 0 163006 800 6 la_data_out[9]
port 257 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 la_oenb[0]
port 258 nsew signal input
rlabel metal2 s 208030 0 208086 800 6 la_oenb[100]
port 259 nsew signal input
rlabel metal3 s 221715 127848 222515 127968 6 la_oenb[101]
port 260 nsew signal input
rlabel metal2 s 169390 223859 169446 224659 6 la_oenb[102]
port 261 nsew signal input
rlabel metal3 s 221715 101328 222515 101448 6 la_oenb[103]
port 262 nsew signal input
rlabel metal3 s 0 181568 800 181688 6 la_oenb[104]
port 263 nsew signal input
rlabel metal3 s 0 133288 800 133408 6 la_oenb[105]
port 264 nsew signal input
rlabel metal3 s 221715 8168 222515 8288 6 la_oenb[106]
port 265 nsew signal input
rlabel metal2 s 151358 223859 151414 224659 6 la_oenb[107]
port 266 nsew signal input
rlabel metal2 s 194506 0 194562 800 6 la_oenb[108]
port 267 nsew signal input
rlabel metal2 s 30930 223859 30986 224659 6 la_oenb[109]
port 268 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 la_oenb[10]
port 269 nsew signal input
rlabel metal3 s 221715 99288 222515 99408 6 la_oenb[110]
port 270 nsew signal input
rlabel metal2 s 10966 223859 11022 224659 6 la_oenb[111]
port 271 nsew signal input
rlabel metal3 s 221715 135328 222515 135448 6 la_oenb[112]
port 272 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 la_oenb[113]
port 273 nsew signal input
rlabel metal2 s 201590 0 201646 800 6 la_oenb[114]
port 274 nsew signal input
rlabel metal2 s 85670 223859 85726 224659 6 la_oenb[115]
port 275 nsew signal input
rlabel metal2 s 205454 223859 205510 224659 6 la_oenb[116]
port 276 nsew signal input
rlabel metal3 s 221715 159128 222515 159248 6 la_oenb[117]
port 277 nsew signal input
rlabel metal2 s 76654 223859 76710 224659 6 la_oenb[118]
port 278 nsew signal input
rlabel metal2 s 94686 223859 94742 224659 6 la_oenb[119]
port 279 nsew signal input
rlabel metal3 s 221715 27208 222515 27328 6 la_oenb[11]
port 280 nsew signal input
rlabel metal3 s 0 121728 800 121848 6 la_oenb[120]
port 281 nsew signal input
rlabel metal3 s 0 109488 800 109608 6 la_oenb[121]
port 282 nsew signal input
rlabel metal2 s 162306 223859 162362 224659 6 la_oenb[122]
port 283 nsew signal input
rlabel metal2 s 117226 223859 117282 224659 6 la_oenb[123]
port 284 nsew signal input
rlabel metal2 s 33506 223859 33562 224659 6 la_oenb[124]
port 285 nsew signal input
rlabel metal3 s 0 90448 800 90568 6 la_oenb[125]
port 286 nsew signal input
rlabel metal3 s 0 214888 800 215008 6 la_oenb[126]
port 287 nsew signal input
rlabel metal3 s 221715 154368 222515 154488 6 la_oenb[127]
port 288 nsew signal input
rlabel metal3 s 221715 140088 222515 140208 6 la_oenb[12]
port 289 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 la_oenb[13]
port 290 nsew signal input
rlabel metal3 s 221715 125808 222515 125928 6 la_oenb[14]
port 291 nsew signal input
rlabel metal3 s 0 112208 800 112328 6 la_oenb[15]
port 292 nsew signal input
rlabel metal2 s 206098 0 206154 800 6 la_oenb[16]
port 293 nsew signal input
rlabel metal2 s 155866 223859 155922 224659 6 la_oenb[17]
port 294 nsew signal input
rlabel metal2 s 217046 223859 217102 224659 6 la_oenb[18]
port 295 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 la_oenb[19]
port 296 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 la_oenb[1]
port 297 nsew signal input
rlabel metal3 s 221715 41488 222515 41608 6 la_oenb[20]
port 298 nsew signal input
rlabel metal2 s 44454 223859 44510 224659 6 la_oenb[21]
port 299 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 la_oenb[22]
port 300 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 la_oenb[23]
port 301 nsew signal input
rlabel metal2 s 90178 223859 90234 224659 6 la_oenb[24]
port 302 nsew signal input
rlabel metal3 s 0 88408 800 88528 6 la_oenb[25]
port 303 nsew signal input
rlabel metal3 s 221715 206728 222515 206848 6 la_oenb[26]
port 304 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 la_oenb[27]
port 305 nsew signal input
rlabel metal2 s 184846 223859 184902 224659 6 la_oenb[28]
port 306 nsew signal input
rlabel metal3 s 221715 87048 222515 87168 6 la_oenb[29]
port 307 nsew signal input
rlabel metal2 s 167458 0 167514 800 6 la_oenb[2]
port 308 nsew signal input
rlabel metal3 s 0 97928 800 98048 6 la_oenb[30]
port 309 nsew signal input
rlabel metal2 s 160374 0 160430 800 6 la_oenb[31]
port 310 nsew signal input
rlabel metal3 s 0 119008 800 119128 6 la_oenb[32]
port 311 nsew signal input
rlabel metal3 s 0 157768 800 157888 6 la_oenb[33]
port 312 nsew signal input
rlabel metal2 s 215114 0 215170 800 6 la_oenb[34]
port 313 nsew signal input
rlabel metal3 s 221715 53728 222515 53848 6 la_oenb[35]
port 314 nsew signal input
rlabel metal2 s 83094 223859 83150 224659 6 la_oenb[36]
port 315 nsew signal input
rlabel metal3 s 221715 187688 222515 187808 6 la_oenb[37]
port 316 nsew signal input
rlabel metal3 s 0 188368 800 188488 6 la_oenb[38]
port 317 nsew signal input
rlabel metal3 s 0 205368 800 205488 6 la_oenb[39]
port 318 nsew signal input
rlabel metal3 s 0 197888 800 198008 6 la_oenb[3]
port 319 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 la_oenb[40]
port 320 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 la_oenb[41]
port 321 nsew signal input
rlabel metal3 s 221715 110848 222515 110968 6 la_oenb[42]
port 322 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 la_oenb[43]
port 323 nsew signal input
rlabel metal2 s 160374 223859 160430 224659 6 la_oenb[44]
port 324 nsew signal input
rlabel metal2 s 212538 223859 212594 224659 6 la_oenb[45]
port 325 nsew signal input
rlabel metal2 s 24490 223859 24546 224659 6 la_oenb[46]
port 326 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 la_oenb[47]
port 327 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 la_oenb[48]
port 328 nsew signal input
rlabel metal2 s 218978 223859 219034 224659 6 la_oenb[49]
port 329 nsew signal input
rlabel metal3 s 0 145528 800 145648 6 la_oenb[4]
port 330 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 la_oenb[50]
port 331 nsew signal input
rlabel metal3 s 221715 65968 222515 66088 6 la_oenb[51]
port 332 nsew signal input
rlabel metal2 s 149426 0 149482 800 6 la_oenb[52]
port 333 nsew signal input
rlabel metal2 s 191930 223859 191986 224659 6 la_oenb[53]
port 334 nsew signal input
rlabel metal2 s 63130 223859 63186 224659 6 la_oenb[54]
port 335 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_oenb[55]
port 336 nsew signal input
rlabel metal3 s 221715 130568 222515 130688 6 la_oenb[56]
port 337 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 la_oenb[57]
port 338 nsew signal input
rlabel metal3 s 221715 61208 222515 61328 6 la_oenb[58]
port 339 nsew signal input
rlabel metal3 s 0 128528 800 128648 6 la_oenb[59]
port 340 nsew signal input
rlabel metal3 s 221715 1368 222515 1488 6 la_oenb[5]
port 341 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 la_oenb[60]
port 342 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 la_oenb[61]
port 343 nsew signal input
rlabel metal3 s 221715 91808 222515 91928 6 la_oenb[62]
port 344 nsew signal input
rlabel metal2 s 180338 223859 180394 224659 6 la_oenb[63]
port 345 nsew signal input
rlabel metal3 s 221715 197208 222515 197328 6 la_oenb[64]
port 346 nsew signal input
rlabel metal3 s 221715 6128 222515 6248 6 la_oenb[65]
port 347 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 la_oenb[66]
port 348 nsew signal input
rlabel metal3 s 221715 123088 222515 123208 6 la_oenb[67]
port 349 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 la_oenb[68]
port 350 nsew signal input
rlabel metal3 s 221715 204688 222515 204808 6 la_oenb[69]
port 351 nsew signal input
rlabel metal2 s 171322 223859 171378 224659 6 la_oenb[6]
port 352 nsew signal input
rlabel metal3 s 221715 20408 222515 20528 6 la_oenb[70]
port 353 nsew signal input
rlabel metal2 s 164882 223859 164938 224659 6 la_oenb[71]
port 354 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 la_oenb[72]
port 355 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 la_oenb[73]
port 356 nsew signal input
rlabel metal2 s 144918 0 144974 800 6 la_oenb[74]
port 357 nsew signal input
rlabel metal2 s 18 0 74 800 6 la_oenb[75]
port 358 nsew signal input
rlabel metal2 s 171966 0 172022 800 6 la_oenb[76]
port 359 nsew signal input
rlabel metal3 s 0 114248 800 114368 6 la_oenb[77]
port 360 nsew signal input
rlabel metal3 s 0 202648 800 202768 6 la_oenb[78]
port 361 nsew signal input
rlabel metal2 s 67638 223859 67694 224659 6 la_oenb[79]
port 362 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 la_oenb[7]
port 363 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 la_oenb[80]
port 364 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 la_oenb[81]
port 365 nsew signal input
rlabel metal2 s 119158 223859 119214 224659 6 la_oenb[82]
port 366 nsew signal input
rlabel metal2 s 72146 223859 72202 224659 6 la_oenb[83]
port 367 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 la_oenb[84]
port 368 nsew signal input
rlabel metal2 s 157798 223859 157854 224659 6 la_oenb[85]
port 369 nsew signal input
rlabel metal3 s 221715 58488 222515 58608 6 la_oenb[86]
port 370 nsew signal input
rlabel metal3 s 0 153008 800 153128 6 la_oenb[87]
port 371 nsew signal input
rlabel metal3 s 221715 170688 222515 170808 6 la_oenb[88]
port 372 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_oenb[89]
port 373 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_oenb[8]
port 374 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 la_oenb[90]
port 375 nsew signal input
rlabel metal3 s 221715 163888 222515 164008 6 la_oenb[91]
port 376 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 la_oenb[92]
port 377 nsew signal input
rlabel metal2 s 148782 223859 148838 224659 6 la_oenb[93]
port 378 nsew signal input
rlabel metal2 s 146850 223859 146906 224659 6 la_oenb[94]
port 379 nsew signal input
rlabel metal3 s 0 212848 800 212968 6 la_oenb[95]
port 380 nsew signal input
rlabel metal2 s 28998 223859 29054 224659 6 la_oenb[96]
port 381 nsew signal input
rlabel metal2 s 158442 0 158498 800 6 la_oenb[97]
port 382 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 la_oenb[98]
port 383 nsew signal input
rlabel metal3 s 0 191088 800 191208 6 la_oenb[99]
port 384 nsew signal input
rlabel metal3 s 221715 108808 222515 108928 6 la_oenb[9]
port 385 nsew signal input
rlabel metal4 s 4208 2128 4528 222000 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 222000 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 222000 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 222000 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 222000 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 222000 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 222000 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 222000 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 222000 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 222000 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 222000 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 222000 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 222000 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 222000 6 vssd1
port 387 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 222000 6 vssd1
port 387 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 222515 224659
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 60808848
string GDS_FILE /home/drewarosa/RISC-V-Single-Cycle-CPU-Core/openlane/risc_v/runs/22_08_30_17_25/results/signoff/RISC_V.magic.gds
string GDS_START 1085442
<< end >>

